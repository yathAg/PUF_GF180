magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect 5753 27606 7054 27622
rect 13132 27606 14433 27622
rect 1479 27468 7054 27606
rect 8858 27468 14433 27606
rect 23617 27562 24919 27681
rect 1479 26958 8341 27468
rect 8858 26958 15720 27468
rect 1479 26945 7054 26958
rect 8858 26945 14433 26958
rect 1479 25077 5469 26945
rect 8858 25156 12848 26945
rect 16524 25287 23175 27042
rect 23617 26980 26150 27562
rect 23617 26945 24919 26980
rect 6472 25135 7008 25136
rect 5958 25077 7008 25135
rect 1394 25058 7008 25077
rect 7649 25077 12848 25156
rect 13851 25135 14387 25136
rect 13337 25077 14387 25135
rect 7649 25058 14387 25077
rect 15028 25058 16138 25156
rect 1394 24683 16138 25058
rect 1637 22243 16138 24683
rect 16524 24513 28667 25287
rect 16438 24039 28667 24513
rect 1637 22242 8745 22243
rect 9016 22242 16124 22243
rect 1637 21381 6541 22242
rect 5264 21338 6541 21381
rect 7219 21338 8232 22242
rect 9016 21381 13920 22242
rect 12643 21338 13920 21381
rect 14598 21338 15611 22242
rect 16524 21769 28667 24039
rect 23173 21740 28667 21769
rect 5911 21336 6541 21338
rect 7602 21336 8232 21338
rect 13290 21336 13920 21338
rect 14981 21336 15611 21338
rect 7114 19567 7116 19568
rect 14493 19567 14495 19568
rect 23837 19567 24981 19568
rect 25528 19567 26671 19568
rect 27218 19567 28362 19568
rect 5489 18378 8806 19567
rect 12868 18378 16185 19567
rect 23353 18378 28362 19567
rect 1815 16637 20347 17092
rect 1815 16636 20281 16637
rect 1815 11908 20141 16636
rect 7270 8117 13921 8427
rect 1839 7013 13921 8117
rect 20706 8070 21480 8586
rect 1839 6558 14007 7013
rect 20739 6709 20904 6756
rect 1839 5143 13921 6558
rect 24661 5866 24705 10029
rect 25867 5253 25991 10029
rect 27119 5388 27222 10029
rect 1839 5113 7333 5143
rect 2019 1751 7028 2941
rect 8581 1311 9883 1422
rect 8581 1303 13811 1311
rect 7599 721 13811 1303
rect 8581 693 13811 721
rect 8581 686 9883 693
<< mvnmos >>
rect 1734 27745 1854 28653
rect 1958 27745 2078 28653
rect 2182 27745 2302 28653
rect 2406 27745 2526 28653
rect 2630 27745 2750 28653
rect 2854 27745 2974 28653
rect 3078 27745 3198 28653
rect 3302 27745 3422 28653
rect 3526 27745 3646 28653
rect 3750 27745 3870 28653
rect 3974 27745 4094 28653
rect 4198 27745 4318 28653
rect 4422 27745 4542 28653
rect 4646 27745 4766 28653
rect 4870 27745 4990 28653
rect 5094 27745 5214 28653
rect 6008 27821 6128 28095
rect 6232 27821 6352 28095
rect 7602 27817 7722 28009
rect 9113 27745 9233 28653
rect 9337 27745 9457 28653
rect 9561 27745 9681 28653
rect 9785 27745 9905 28653
rect 10009 27745 10129 28653
rect 10233 27745 10353 28653
rect 10457 27745 10577 28653
rect 10681 27745 10801 28653
rect 10905 27745 11025 28653
rect 11129 27745 11249 28653
rect 11353 27745 11473 28653
rect 11577 27745 11697 28653
rect 11801 27745 11921 28653
rect 12025 27745 12145 28653
rect 12249 27745 12369 28653
rect 12473 27745 12593 28653
rect 13387 27821 13507 28095
rect 13611 27821 13731 28095
rect 14981 27817 15101 28009
rect 6166 25336 6286 26744
rect 6680 25415 6800 26459
rect 7857 25336 7977 26744
rect 8371 25415 8491 26459
rect 16779 27181 16899 28089
rect 17003 27181 17123 28089
rect 17227 27181 17347 28089
rect 17451 27181 17571 28089
rect 17675 27181 17795 28089
rect 17899 27181 18019 28089
rect 18413 27181 18533 28089
rect 18637 27181 18757 28089
rect 18861 27181 18981 28089
rect 19085 27181 19205 28089
rect 19309 27181 19429 28089
rect 19533 27181 19653 28089
rect 20046 27181 20166 28089
rect 20270 27181 20390 28089
rect 20494 27181 20614 28089
rect 20718 27181 20838 28089
rect 20942 27181 21062 28089
rect 21166 27181 21286 28089
rect 21680 27181 21800 28089
rect 21904 27181 22024 28089
rect 22128 27181 22248 28089
rect 22352 27181 22472 28089
rect 22576 27181 22696 28089
rect 22800 27181 22920 28089
rect 23872 27821 23992 28203
rect 24096 27821 24216 28203
rect 25467 27817 25587 28089
rect 13545 25336 13665 26744
rect 14059 25415 14179 26459
rect 15236 25336 15356 26744
rect 15750 25415 15870 26459
rect 24031 25427 24151 26743
rect 24545 25427 24665 26743
rect 25721 25427 25841 26743
rect 26235 25427 26355 26743
rect 27412 25427 27532 26743
rect 27926 25427 28046 26743
rect 1892 18101 2012 20551
rect 2116 18101 2236 20551
rect 2920 18101 3040 20551
rect 3144 18101 3264 20551
rect 3684 18101 3804 20551
rect 3908 18101 4028 20551
rect 4712 18101 4832 20551
rect 4936 18101 5056 20551
rect 9271 18101 9391 20551
rect 9495 18101 9615 20551
rect 10299 18101 10419 20551
rect 10523 18101 10643 20551
rect 11063 18101 11183 20551
rect 11287 18101 11407 20551
rect 12091 18101 12211 20551
rect 12315 18101 12435 20551
rect 16779 18043 16899 20538
rect 17003 18043 17123 20538
rect 17227 18043 17347 20538
rect 17451 18043 17571 20538
rect 17675 18043 17795 20538
rect 17899 18043 18019 20538
rect 18413 18043 18533 20538
rect 18637 18043 18757 20538
rect 18861 18043 18981 20538
rect 19085 18043 19205 20538
rect 19309 18043 19429 20538
rect 19533 18043 19653 20538
rect 20046 18043 20166 20538
rect 20270 18043 20390 20538
rect 20494 18043 20614 20538
rect 20718 18043 20838 20538
rect 20942 18043 21062 20538
rect 21166 18043 21286 20538
rect 21680 18043 21800 20538
rect 21904 18043 22024 20538
rect 22128 18043 22248 20538
rect 22352 18043 22472 20538
rect 22576 18043 22696 20538
rect 22800 18043 22920 20538
rect 2070 9954 2190 11770
rect 2518 9954 2638 11770
rect 2742 9954 2862 11770
rect 2966 9954 3086 11770
rect 3190 9954 3310 11770
rect 3638 9954 3758 11770
rect 3862 9954 3982 11770
rect 4086 9954 4206 11770
rect 4310 9954 4430 11770
rect 4758 9954 4878 11770
rect 4982 9954 5102 11770
rect 5206 9954 5326 11770
rect 5430 9954 5550 11770
rect 5878 9954 5998 11770
rect 6102 9954 6222 11770
rect 6326 9954 6446 11770
rect 6550 9954 6670 11770
rect 6998 9954 7118 11770
rect 7222 9954 7342 11770
rect 7446 9954 7566 11770
rect 7670 9954 7790 11770
rect 8118 9954 8238 11770
rect 8342 9954 8462 11770
rect 8566 9954 8686 11770
rect 8790 9954 8910 11770
rect 9238 9954 9358 11770
rect 9462 9954 9582 11770
rect 9686 9954 9806 11770
rect 9910 9954 10030 11770
rect 10358 9954 10478 11770
rect 10582 9954 10702 11770
rect 10806 9954 10926 11770
rect 11030 9954 11150 11770
rect 11478 9954 11598 11770
rect 11702 9954 11822 11770
rect 11926 9954 12046 11770
rect 12150 9954 12270 11770
rect 12598 9954 12718 11770
rect 12822 9954 12942 11770
rect 13046 9954 13166 11770
rect 13270 9954 13390 11770
rect 13718 9954 13838 11770
rect 13942 9954 14062 11770
rect 14166 9954 14286 11770
rect 14390 9954 14510 11770
rect 14838 9954 14958 11770
rect 15062 9954 15182 11770
rect 15286 9954 15406 11770
rect 15510 9954 15630 11770
rect 15958 9954 16078 11770
rect 16182 9954 16302 11770
rect 16406 9954 16526 11770
rect 16630 9954 16750 11770
rect 17078 9954 17198 11770
rect 17302 9954 17422 11770
rect 17526 9954 17646 11770
rect 17750 9954 17870 11770
rect 18198 9954 18318 11770
rect 18422 9954 18542 11770
rect 18646 9954 18766 11770
rect 18870 9954 18990 11770
rect 19318 9954 19438 11770
rect 19542 9954 19662 11770
rect 19766 9954 19886 11770
rect 2696 8257 2816 9165
rect 3210 8257 3330 9165
rect 4387 8257 4507 9165
rect 4901 8257 5021 9165
rect 6078 8257 6198 9165
rect 6592 8257 6712 9165
rect 7525 8567 7645 9021
rect 7749 8567 7869 9021
rect 7973 8567 8093 9021
rect 8197 8567 8317 9021
rect 8421 8567 8541 9021
rect 8645 8567 8765 9021
rect 9158 8567 9278 9021
rect 9382 8567 9502 9021
rect 9606 8567 9726 9021
rect 9830 8567 9950 9021
rect 10054 8567 10174 9021
rect 10278 8567 10398 9021
rect 10792 8567 10912 9021
rect 11016 8567 11136 9021
rect 11240 8567 11360 9021
rect 11464 8567 11584 9021
rect 11688 8567 11808 9021
rect 11912 8567 12032 9021
rect 12426 8567 12546 9021
rect 12650 8567 12770 9021
rect 12874 8567 12994 9021
rect 13098 8567 13218 9021
rect 13322 8567 13442 9021
rect 13546 8567 13666 9021
rect 7526 2550 7646 3912
rect 7748 2550 7868 3912
rect 7972 2550 8092 3912
rect 8198 2550 8318 3912
rect 8422 2550 8542 3912
rect 8644 2550 8764 3912
rect 9159 2550 9279 3912
rect 9381 2550 9501 3912
rect 9605 2550 9725 3912
rect 9831 2550 9951 3912
rect 10055 2550 10175 3912
rect 10277 2550 10397 3912
rect 10793 2550 10913 3912
rect 11015 2550 11135 3912
rect 11239 2550 11359 3912
rect 11465 2550 11585 3912
rect 11689 2550 11809 3912
rect 11911 2550 12031 3912
rect 12427 2550 12547 3912
rect 12649 2550 12769 3912
rect 12873 2550 12993 3912
rect 13099 2550 13219 3912
rect 13323 2550 13443 3912
rect 13545 2550 13665 3912
rect 7913 1557 8033 1829
rect 9283 1562 9403 1944
rect 9507 1562 9627 1944
<< mvpmos >>
rect 1734 25197 1854 27465
rect 1958 25197 2078 27465
rect 2182 25197 2302 27465
rect 2406 25197 2526 27465
rect 2630 25197 2750 27465
rect 2854 25197 2974 27465
rect 3078 25197 3198 27465
rect 3302 25197 3422 27465
rect 3526 25197 3646 27465
rect 3750 25197 3870 27465
rect 3974 25197 4094 27465
rect 4198 25197 4318 27465
rect 4422 25197 4542 27465
rect 4646 25197 4766 27465
rect 4870 25197 4990 27465
rect 5094 25197 5214 27465
rect 6008 27086 6128 27427
rect 6231 27086 6351 27427
rect 6456 27086 6576 27427
rect 6679 27086 6799 27427
rect 7484 27100 7604 27328
rect 7708 27100 7828 27328
rect 9113 25197 9233 27465
rect 9337 25197 9457 27465
rect 9561 25197 9681 27465
rect 9785 25197 9905 27465
rect 10009 25197 10129 27465
rect 10233 25197 10353 27465
rect 10457 25197 10577 27465
rect 10681 25197 10801 27465
rect 10905 25197 11025 27465
rect 11129 25197 11249 27465
rect 11353 25197 11473 27465
rect 11577 25197 11697 27465
rect 11801 25197 11921 27465
rect 12025 25197 12145 27465
rect 12249 25197 12369 27465
rect 12473 25197 12593 27465
rect 13387 27086 13507 27427
rect 13610 27086 13730 27427
rect 13835 27086 13955 27427
rect 14058 27086 14178 27427
rect 14863 27100 14983 27328
rect 15087 27100 15207 27328
rect 23872 27086 23992 27541
rect 24096 27086 24216 27541
rect 24320 27086 24440 27541
rect 24544 27086 24664 27541
rect 25348 27100 25468 27442
rect 25572 27100 25692 27442
rect 1892 21523 2012 24563
rect 2116 21523 2236 24563
rect 2920 21523 3040 24563
rect 3144 21523 3264 24563
rect 3684 21523 3804 24563
rect 3908 21523 4028 24563
rect 4712 21523 4832 24563
rect 4936 21523 5056 24563
rect 6166 21477 6286 25015
rect 6680 22384 6800 25016
rect 7857 21477 7977 25015
rect 8371 22384 8491 25016
rect 9271 21523 9391 24563
rect 9495 21523 9615 24563
rect 10299 21523 10419 24563
rect 10523 21523 10643 24563
rect 11063 21523 11183 24563
rect 11287 21523 11407 24563
rect 12091 21523 12211 24563
rect 12315 21523 12435 24563
rect 13545 21477 13665 25015
rect 14059 22384 14179 25016
rect 15236 21477 15356 25015
rect 15750 22384 15870 25016
rect 16779 24633 16899 26901
rect 17003 24633 17123 26901
rect 17227 24633 17347 26901
rect 17451 24633 17571 26901
rect 17675 24633 17795 26901
rect 17899 24633 18019 26901
rect 18413 24633 18533 26901
rect 18637 24633 18757 26901
rect 18861 24633 18981 26901
rect 19085 24633 19205 26901
rect 19309 24633 19429 26901
rect 19533 24633 19653 26901
rect 20046 24633 20166 26901
rect 20270 24633 20390 26901
rect 20494 24633 20614 26901
rect 20718 24633 20838 26901
rect 20942 24633 21062 26901
rect 21166 24633 21286 26901
rect 21680 24633 21800 26901
rect 21904 24633 22024 26901
rect 22128 24633 22248 26901
rect 22352 24633 22472 26901
rect 22576 24633 22696 26901
rect 22800 24633 22920 26901
rect 16779 21911 16899 23997
rect 17003 21911 17123 23997
rect 17227 21911 17347 23997
rect 17451 21911 17571 23997
rect 17675 21911 17795 23997
rect 17899 21911 18019 23997
rect 18413 21911 18533 23997
rect 18637 21911 18757 23997
rect 18861 21911 18981 23997
rect 19085 21911 19205 23997
rect 19309 21911 19429 23997
rect 19533 21911 19653 23997
rect 20046 21911 20166 23997
rect 20270 21911 20390 23997
rect 20494 21911 20614 23997
rect 20718 21911 20838 23997
rect 20942 21911 21062 23997
rect 21166 21911 21286 23997
rect 21680 21911 21800 23997
rect 21904 21911 22024 23997
rect 22128 21911 22248 23997
rect 22352 21911 22472 23997
rect 22576 21911 22696 23997
rect 22800 21911 22920 23997
rect 24031 21881 24151 25147
rect 24545 21881 24665 25147
rect 25721 21881 25841 25147
rect 26235 21881 26355 25147
rect 27412 21881 27532 25147
rect 27926 21881 28046 25147
rect 2070 12585 2190 16585
rect 2518 12585 2638 16585
rect 2742 12585 2862 16585
rect 2966 12585 3086 16585
rect 3190 12585 3310 16585
rect 3638 12585 3758 16585
rect 3862 12585 3982 16585
rect 4086 12585 4206 16585
rect 4310 12585 4430 16585
rect 4758 12585 4878 16585
rect 4982 12585 5102 16585
rect 5206 12585 5326 16585
rect 5430 12585 5550 16585
rect 5878 12585 5998 16585
rect 6102 12585 6222 16585
rect 6326 12585 6446 16585
rect 6550 12585 6670 16585
rect 6998 12585 7118 16585
rect 7222 12585 7342 16585
rect 7446 12585 7566 16585
rect 7670 12585 7790 16585
rect 8118 12585 8238 16585
rect 8342 12585 8462 16585
rect 8566 12585 8686 16585
rect 8790 12585 8910 16585
rect 9238 12585 9358 16585
rect 9462 12585 9582 16585
rect 9686 12585 9806 16585
rect 9910 12585 10030 16585
rect 10358 12585 10478 16585
rect 10582 12585 10702 16585
rect 10806 12585 10926 16585
rect 11030 12585 11150 16585
rect 11478 12585 11598 16585
rect 11702 12585 11822 16585
rect 11926 12585 12046 16585
rect 12150 12585 12270 16585
rect 12598 12585 12718 16585
rect 12822 12585 12942 16585
rect 13046 12585 13166 16585
rect 13270 12585 13390 16585
rect 13718 12585 13838 16585
rect 13942 12585 14062 16585
rect 14166 12585 14286 16585
rect 14390 12585 14510 16585
rect 14838 12585 14958 16585
rect 15062 12585 15182 16585
rect 15286 12585 15406 16585
rect 15510 12585 15630 16585
rect 15958 12585 16078 16585
rect 16182 12585 16302 16585
rect 16406 12585 16526 16585
rect 16630 12585 16750 16585
rect 17078 12585 17198 16585
rect 17302 12585 17422 16585
rect 17526 12585 17646 16585
rect 17750 12585 17870 16585
rect 18198 12585 18318 16585
rect 18422 12585 18542 16585
rect 18646 12585 18766 16585
rect 18870 12585 18990 16585
rect 19318 12585 19438 16585
rect 19542 12585 19662 16585
rect 19766 12585 19886 16585
rect 2696 5255 2816 7977
rect 3210 5255 3330 7977
rect 4387 5255 4507 7977
rect 4901 5255 5021 7977
rect 6078 5255 6198 7977
rect 6592 5255 6712 7977
rect 7525 7132 7645 8286
rect 7749 7132 7869 8286
rect 7973 7132 8093 8286
rect 8197 7132 8317 8286
rect 8421 7132 8541 8286
rect 8645 7132 8765 8286
rect 9158 7132 9278 8286
rect 9382 7132 9502 8286
rect 9606 7132 9726 8286
rect 9830 7132 9950 8286
rect 10054 7132 10174 8286
rect 10278 7132 10398 8286
rect 10792 7132 10912 8286
rect 11016 7132 11136 8286
rect 11240 7132 11360 8286
rect 11464 7132 11584 8286
rect 11688 7132 11808 8286
rect 11912 7132 12032 8286
rect 12426 7132 12546 8286
rect 12650 7132 12770 8286
rect 12874 7132 12994 8286
rect 13098 7132 13218 8286
rect 13322 7132 13442 8286
rect 13546 7132 13666 8286
rect 7525 5285 7645 6419
rect 7749 5285 7869 6419
rect 7973 5285 8093 6419
rect 8197 5285 8317 6419
rect 8421 5285 8541 6419
rect 8645 5285 8765 6419
rect 9158 5285 9278 6419
rect 9382 5285 9502 6419
rect 9606 5285 9726 6419
rect 9830 5285 9950 6419
rect 10054 5285 10174 6419
rect 10278 5285 10398 6419
rect 10792 5285 10912 6419
rect 11016 5285 11136 6419
rect 11240 5285 11360 6419
rect 11464 5285 11584 6419
rect 11688 5285 11808 6419
rect 11912 5285 12032 6419
rect 12426 5285 12546 6419
rect 12650 5285 12770 6419
rect 12874 5285 12994 6419
rect 13098 5285 13218 6419
rect 13322 5285 13442 6419
rect 13546 5285 13666 6419
rect 7807 841 7927 1183
rect 8031 841 8151 1183
rect 8836 827 8956 1282
rect 9060 827 9180 1282
rect 9284 827 9404 1282
rect 9508 827 9628 1282
<< mvndiff >>
rect 1646 28640 1734 28653
rect 1646 28594 1659 28640
rect 1705 28594 1734 28640
rect 1646 28535 1734 28594
rect 1646 28489 1659 28535
rect 1705 28489 1734 28535
rect 1646 28430 1734 28489
rect 1646 28384 1659 28430
rect 1705 28384 1734 28430
rect 1646 28325 1734 28384
rect 1646 28279 1659 28325
rect 1705 28279 1734 28325
rect 1646 28220 1734 28279
rect 1646 28174 1659 28220
rect 1705 28174 1734 28220
rect 1646 28116 1734 28174
rect 1646 28070 1659 28116
rect 1705 28070 1734 28116
rect 1646 28012 1734 28070
rect 1646 27966 1659 28012
rect 1705 27966 1734 28012
rect 1646 27908 1734 27966
rect 1646 27862 1659 27908
rect 1705 27862 1734 27908
rect 1646 27804 1734 27862
rect 1646 27758 1659 27804
rect 1705 27758 1734 27804
rect 1646 27745 1734 27758
rect 1854 28640 1958 28653
rect 1854 28594 1883 28640
rect 1929 28594 1958 28640
rect 1854 28535 1958 28594
rect 1854 28489 1883 28535
rect 1929 28489 1958 28535
rect 1854 28430 1958 28489
rect 1854 28384 1883 28430
rect 1929 28384 1958 28430
rect 1854 28325 1958 28384
rect 1854 28279 1883 28325
rect 1929 28279 1958 28325
rect 1854 28220 1958 28279
rect 1854 28174 1883 28220
rect 1929 28174 1958 28220
rect 1854 28116 1958 28174
rect 1854 28070 1883 28116
rect 1929 28070 1958 28116
rect 1854 28012 1958 28070
rect 1854 27966 1883 28012
rect 1929 27966 1958 28012
rect 1854 27908 1958 27966
rect 1854 27862 1883 27908
rect 1929 27862 1958 27908
rect 1854 27804 1958 27862
rect 1854 27758 1883 27804
rect 1929 27758 1958 27804
rect 1854 27745 1958 27758
rect 2078 28640 2182 28653
rect 2078 28594 2107 28640
rect 2153 28594 2182 28640
rect 2078 28535 2182 28594
rect 2078 28489 2107 28535
rect 2153 28489 2182 28535
rect 2078 28430 2182 28489
rect 2078 28384 2107 28430
rect 2153 28384 2182 28430
rect 2078 28325 2182 28384
rect 2078 28279 2107 28325
rect 2153 28279 2182 28325
rect 2078 28220 2182 28279
rect 2078 28174 2107 28220
rect 2153 28174 2182 28220
rect 2078 28116 2182 28174
rect 2078 28070 2107 28116
rect 2153 28070 2182 28116
rect 2078 28012 2182 28070
rect 2078 27966 2107 28012
rect 2153 27966 2182 28012
rect 2078 27908 2182 27966
rect 2078 27862 2107 27908
rect 2153 27862 2182 27908
rect 2078 27804 2182 27862
rect 2078 27758 2107 27804
rect 2153 27758 2182 27804
rect 2078 27745 2182 27758
rect 2302 28640 2406 28653
rect 2302 28594 2331 28640
rect 2377 28594 2406 28640
rect 2302 28535 2406 28594
rect 2302 28489 2331 28535
rect 2377 28489 2406 28535
rect 2302 28430 2406 28489
rect 2302 28384 2331 28430
rect 2377 28384 2406 28430
rect 2302 28325 2406 28384
rect 2302 28279 2331 28325
rect 2377 28279 2406 28325
rect 2302 28220 2406 28279
rect 2302 28174 2331 28220
rect 2377 28174 2406 28220
rect 2302 28116 2406 28174
rect 2302 28070 2331 28116
rect 2377 28070 2406 28116
rect 2302 28012 2406 28070
rect 2302 27966 2331 28012
rect 2377 27966 2406 28012
rect 2302 27908 2406 27966
rect 2302 27862 2331 27908
rect 2377 27862 2406 27908
rect 2302 27804 2406 27862
rect 2302 27758 2331 27804
rect 2377 27758 2406 27804
rect 2302 27745 2406 27758
rect 2526 28640 2630 28653
rect 2526 28594 2555 28640
rect 2601 28594 2630 28640
rect 2526 28535 2630 28594
rect 2526 28489 2555 28535
rect 2601 28489 2630 28535
rect 2526 28430 2630 28489
rect 2526 28384 2555 28430
rect 2601 28384 2630 28430
rect 2526 28325 2630 28384
rect 2526 28279 2555 28325
rect 2601 28279 2630 28325
rect 2526 28220 2630 28279
rect 2526 28174 2555 28220
rect 2601 28174 2630 28220
rect 2526 28116 2630 28174
rect 2526 28070 2555 28116
rect 2601 28070 2630 28116
rect 2526 28012 2630 28070
rect 2526 27966 2555 28012
rect 2601 27966 2630 28012
rect 2526 27908 2630 27966
rect 2526 27862 2555 27908
rect 2601 27862 2630 27908
rect 2526 27804 2630 27862
rect 2526 27758 2555 27804
rect 2601 27758 2630 27804
rect 2526 27745 2630 27758
rect 2750 28640 2854 28653
rect 2750 28594 2779 28640
rect 2825 28594 2854 28640
rect 2750 28535 2854 28594
rect 2750 28489 2779 28535
rect 2825 28489 2854 28535
rect 2750 28430 2854 28489
rect 2750 28384 2779 28430
rect 2825 28384 2854 28430
rect 2750 28325 2854 28384
rect 2750 28279 2779 28325
rect 2825 28279 2854 28325
rect 2750 28220 2854 28279
rect 2750 28174 2779 28220
rect 2825 28174 2854 28220
rect 2750 28116 2854 28174
rect 2750 28070 2779 28116
rect 2825 28070 2854 28116
rect 2750 28012 2854 28070
rect 2750 27966 2779 28012
rect 2825 27966 2854 28012
rect 2750 27908 2854 27966
rect 2750 27862 2779 27908
rect 2825 27862 2854 27908
rect 2750 27804 2854 27862
rect 2750 27758 2779 27804
rect 2825 27758 2854 27804
rect 2750 27745 2854 27758
rect 2974 28640 3078 28653
rect 2974 28594 3003 28640
rect 3049 28594 3078 28640
rect 2974 28535 3078 28594
rect 2974 28489 3003 28535
rect 3049 28489 3078 28535
rect 2974 28430 3078 28489
rect 2974 28384 3003 28430
rect 3049 28384 3078 28430
rect 2974 28325 3078 28384
rect 2974 28279 3003 28325
rect 3049 28279 3078 28325
rect 2974 28220 3078 28279
rect 2974 28174 3003 28220
rect 3049 28174 3078 28220
rect 2974 28116 3078 28174
rect 2974 28070 3003 28116
rect 3049 28070 3078 28116
rect 2974 28012 3078 28070
rect 2974 27966 3003 28012
rect 3049 27966 3078 28012
rect 2974 27908 3078 27966
rect 2974 27862 3003 27908
rect 3049 27862 3078 27908
rect 2974 27804 3078 27862
rect 2974 27758 3003 27804
rect 3049 27758 3078 27804
rect 2974 27745 3078 27758
rect 3198 28640 3302 28653
rect 3198 28594 3227 28640
rect 3273 28594 3302 28640
rect 3198 28535 3302 28594
rect 3198 28489 3227 28535
rect 3273 28489 3302 28535
rect 3198 28430 3302 28489
rect 3198 28384 3227 28430
rect 3273 28384 3302 28430
rect 3198 28325 3302 28384
rect 3198 28279 3227 28325
rect 3273 28279 3302 28325
rect 3198 28220 3302 28279
rect 3198 28174 3227 28220
rect 3273 28174 3302 28220
rect 3198 28116 3302 28174
rect 3198 28070 3227 28116
rect 3273 28070 3302 28116
rect 3198 28012 3302 28070
rect 3198 27966 3227 28012
rect 3273 27966 3302 28012
rect 3198 27908 3302 27966
rect 3198 27862 3227 27908
rect 3273 27862 3302 27908
rect 3198 27804 3302 27862
rect 3198 27758 3227 27804
rect 3273 27758 3302 27804
rect 3198 27745 3302 27758
rect 3422 28640 3526 28653
rect 3422 28594 3451 28640
rect 3497 28594 3526 28640
rect 3422 28535 3526 28594
rect 3422 28489 3451 28535
rect 3497 28489 3526 28535
rect 3422 28430 3526 28489
rect 3422 28384 3451 28430
rect 3497 28384 3526 28430
rect 3422 28325 3526 28384
rect 3422 28279 3451 28325
rect 3497 28279 3526 28325
rect 3422 28220 3526 28279
rect 3422 28174 3451 28220
rect 3497 28174 3526 28220
rect 3422 28116 3526 28174
rect 3422 28070 3451 28116
rect 3497 28070 3526 28116
rect 3422 28012 3526 28070
rect 3422 27966 3451 28012
rect 3497 27966 3526 28012
rect 3422 27908 3526 27966
rect 3422 27862 3451 27908
rect 3497 27862 3526 27908
rect 3422 27804 3526 27862
rect 3422 27758 3451 27804
rect 3497 27758 3526 27804
rect 3422 27745 3526 27758
rect 3646 28640 3750 28653
rect 3646 28594 3675 28640
rect 3721 28594 3750 28640
rect 3646 28535 3750 28594
rect 3646 28489 3675 28535
rect 3721 28489 3750 28535
rect 3646 28430 3750 28489
rect 3646 28384 3675 28430
rect 3721 28384 3750 28430
rect 3646 28325 3750 28384
rect 3646 28279 3675 28325
rect 3721 28279 3750 28325
rect 3646 28220 3750 28279
rect 3646 28174 3675 28220
rect 3721 28174 3750 28220
rect 3646 28116 3750 28174
rect 3646 28070 3675 28116
rect 3721 28070 3750 28116
rect 3646 28012 3750 28070
rect 3646 27966 3675 28012
rect 3721 27966 3750 28012
rect 3646 27908 3750 27966
rect 3646 27862 3675 27908
rect 3721 27862 3750 27908
rect 3646 27804 3750 27862
rect 3646 27758 3675 27804
rect 3721 27758 3750 27804
rect 3646 27745 3750 27758
rect 3870 28640 3974 28653
rect 3870 28594 3899 28640
rect 3945 28594 3974 28640
rect 3870 28535 3974 28594
rect 3870 28489 3899 28535
rect 3945 28489 3974 28535
rect 3870 28430 3974 28489
rect 3870 28384 3899 28430
rect 3945 28384 3974 28430
rect 3870 28325 3974 28384
rect 3870 28279 3899 28325
rect 3945 28279 3974 28325
rect 3870 28220 3974 28279
rect 3870 28174 3899 28220
rect 3945 28174 3974 28220
rect 3870 28116 3974 28174
rect 3870 28070 3899 28116
rect 3945 28070 3974 28116
rect 3870 28012 3974 28070
rect 3870 27966 3899 28012
rect 3945 27966 3974 28012
rect 3870 27908 3974 27966
rect 3870 27862 3899 27908
rect 3945 27862 3974 27908
rect 3870 27804 3974 27862
rect 3870 27758 3899 27804
rect 3945 27758 3974 27804
rect 3870 27745 3974 27758
rect 4094 28640 4198 28653
rect 4094 28594 4123 28640
rect 4169 28594 4198 28640
rect 4094 28535 4198 28594
rect 4094 28489 4123 28535
rect 4169 28489 4198 28535
rect 4094 28430 4198 28489
rect 4094 28384 4123 28430
rect 4169 28384 4198 28430
rect 4094 28325 4198 28384
rect 4094 28279 4123 28325
rect 4169 28279 4198 28325
rect 4094 28220 4198 28279
rect 4094 28174 4123 28220
rect 4169 28174 4198 28220
rect 4094 28116 4198 28174
rect 4094 28070 4123 28116
rect 4169 28070 4198 28116
rect 4094 28012 4198 28070
rect 4094 27966 4123 28012
rect 4169 27966 4198 28012
rect 4094 27908 4198 27966
rect 4094 27862 4123 27908
rect 4169 27862 4198 27908
rect 4094 27804 4198 27862
rect 4094 27758 4123 27804
rect 4169 27758 4198 27804
rect 4094 27745 4198 27758
rect 4318 28640 4422 28653
rect 4318 28594 4347 28640
rect 4393 28594 4422 28640
rect 4318 28535 4422 28594
rect 4318 28489 4347 28535
rect 4393 28489 4422 28535
rect 4318 28430 4422 28489
rect 4318 28384 4347 28430
rect 4393 28384 4422 28430
rect 4318 28325 4422 28384
rect 4318 28279 4347 28325
rect 4393 28279 4422 28325
rect 4318 28220 4422 28279
rect 4318 28174 4347 28220
rect 4393 28174 4422 28220
rect 4318 28116 4422 28174
rect 4318 28070 4347 28116
rect 4393 28070 4422 28116
rect 4318 28012 4422 28070
rect 4318 27966 4347 28012
rect 4393 27966 4422 28012
rect 4318 27908 4422 27966
rect 4318 27862 4347 27908
rect 4393 27862 4422 27908
rect 4318 27804 4422 27862
rect 4318 27758 4347 27804
rect 4393 27758 4422 27804
rect 4318 27745 4422 27758
rect 4542 28640 4646 28653
rect 4542 28594 4571 28640
rect 4617 28594 4646 28640
rect 4542 28535 4646 28594
rect 4542 28489 4571 28535
rect 4617 28489 4646 28535
rect 4542 28430 4646 28489
rect 4542 28384 4571 28430
rect 4617 28384 4646 28430
rect 4542 28325 4646 28384
rect 4542 28279 4571 28325
rect 4617 28279 4646 28325
rect 4542 28220 4646 28279
rect 4542 28174 4571 28220
rect 4617 28174 4646 28220
rect 4542 28116 4646 28174
rect 4542 28070 4571 28116
rect 4617 28070 4646 28116
rect 4542 28012 4646 28070
rect 4542 27966 4571 28012
rect 4617 27966 4646 28012
rect 4542 27908 4646 27966
rect 4542 27862 4571 27908
rect 4617 27862 4646 27908
rect 4542 27804 4646 27862
rect 4542 27758 4571 27804
rect 4617 27758 4646 27804
rect 4542 27745 4646 27758
rect 4766 28640 4870 28653
rect 4766 28594 4795 28640
rect 4841 28594 4870 28640
rect 4766 28535 4870 28594
rect 4766 28489 4795 28535
rect 4841 28489 4870 28535
rect 4766 28430 4870 28489
rect 4766 28384 4795 28430
rect 4841 28384 4870 28430
rect 4766 28325 4870 28384
rect 4766 28279 4795 28325
rect 4841 28279 4870 28325
rect 4766 28220 4870 28279
rect 4766 28174 4795 28220
rect 4841 28174 4870 28220
rect 4766 28116 4870 28174
rect 4766 28070 4795 28116
rect 4841 28070 4870 28116
rect 4766 28012 4870 28070
rect 4766 27966 4795 28012
rect 4841 27966 4870 28012
rect 4766 27908 4870 27966
rect 4766 27862 4795 27908
rect 4841 27862 4870 27908
rect 4766 27804 4870 27862
rect 4766 27758 4795 27804
rect 4841 27758 4870 27804
rect 4766 27745 4870 27758
rect 4990 28640 5094 28653
rect 4990 28594 5019 28640
rect 5065 28594 5094 28640
rect 4990 28535 5094 28594
rect 4990 28489 5019 28535
rect 5065 28489 5094 28535
rect 4990 28430 5094 28489
rect 4990 28384 5019 28430
rect 5065 28384 5094 28430
rect 4990 28325 5094 28384
rect 4990 28279 5019 28325
rect 5065 28279 5094 28325
rect 4990 28220 5094 28279
rect 4990 28174 5019 28220
rect 5065 28174 5094 28220
rect 4990 28116 5094 28174
rect 4990 28070 5019 28116
rect 5065 28070 5094 28116
rect 4990 28012 5094 28070
rect 4990 27966 5019 28012
rect 5065 27966 5094 28012
rect 4990 27908 5094 27966
rect 4990 27862 5019 27908
rect 5065 27862 5094 27908
rect 4990 27804 5094 27862
rect 4990 27758 5019 27804
rect 5065 27758 5094 27804
rect 4990 27745 5094 27758
rect 5214 28640 5302 28653
rect 5214 28594 5243 28640
rect 5289 28594 5302 28640
rect 5214 28535 5302 28594
rect 5214 28489 5243 28535
rect 5289 28489 5302 28535
rect 5214 28430 5302 28489
rect 5214 28384 5243 28430
rect 5289 28384 5302 28430
rect 5214 28325 5302 28384
rect 5214 28279 5243 28325
rect 5289 28279 5302 28325
rect 5214 28220 5302 28279
rect 5214 28174 5243 28220
rect 5289 28174 5302 28220
rect 5214 28116 5302 28174
rect 9025 28640 9113 28653
rect 9025 28594 9038 28640
rect 9084 28594 9113 28640
rect 9025 28535 9113 28594
rect 9025 28489 9038 28535
rect 9084 28489 9113 28535
rect 9025 28430 9113 28489
rect 9025 28384 9038 28430
rect 9084 28384 9113 28430
rect 9025 28325 9113 28384
rect 9025 28279 9038 28325
rect 9084 28279 9113 28325
rect 9025 28220 9113 28279
rect 9025 28174 9038 28220
rect 9084 28174 9113 28220
rect 5214 28070 5243 28116
rect 5289 28070 5302 28116
rect 9025 28116 9113 28174
rect 5214 28012 5302 28070
rect 5214 27966 5243 28012
rect 5289 27966 5302 28012
rect 5214 27908 5302 27966
rect 5214 27862 5243 27908
rect 5289 27862 5302 27908
rect 5214 27804 5302 27862
rect 5920 28082 6008 28095
rect 5920 27834 5933 28082
rect 5979 27834 6008 28082
rect 5920 27821 6008 27834
rect 6128 28082 6232 28095
rect 6128 27834 6157 28082
rect 6203 27834 6232 28082
rect 6128 27821 6232 27834
rect 6352 28082 6440 28095
rect 6352 27834 6381 28082
rect 6427 27834 6440 28082
rect 6352 27821 6440 27834
rect 9025 28070 9038 28116
rect 9084 28070 9113 28116
rect 9025 28012 9113 28070
rect 5214 27758 5243 27804
rect 5289 27758 5302 27804
rect 5214 27745 5302 27758
rect 7514 27996 7602 28009
rect 7514 27950 7527 27996
rect 7573 27950 7602 27996
rect 7514 27876 7602 27950
rect 7514 27830 7527 27876
rect 7573 27830 7602 27876
rect 7514 27817 7602 27830
rect 7722 27996 7810 28009
rect 7722 27950 7751 27996
rect 7797 27950 7810 27996
rect 7722 27876 7810 27950
rect 7722 27830 7751 27876
rect 7797 27830 7810 27876
rect 7722 27817 7810 27830
rect 9025 27966 9038 28012
rect 9084 27966 9113 28012
rect 9025 27908 9113 27966
rect 9025 27862 9038 27908
rect 9084 27862 9113 27908
rect 9025 27804 9113 27862
rect 9025 27758 9038 27804
rect 9084 27758 9113 27804
rect 9025 27745 9113 27758
rect 9233 28640 9337 28653
rect 9233 28594 9262 28640
rect 9308 28594 9337 28640
rect 9233 28535 9337 28594
rect 9233 28489 9262 28535
rect 9308 28489 9337 28535
rect 9233 28430 9337 28489
rect 9233 28384 9262 28430
rect 9308 28384 9337 28430
rect 9233 28325 9337 28384
rect 9233 28279 9262 28325
rect 9308 28279 9337 28325
rect 9233 28220 9337 28279
rect 9233 28174 9262 28220
rect 9308 28174 9337 28220
rect 9233 28116 9337 28174
rect 9233 28070 9262 28116
rect 9308 28070 9337 28116
rect 9233 28012 9337 28070
rect 9233 27966 9262 28012
rect 9308 27966 9337 28012
rect 9233 27908 9337 27966
rect 9233 27862 9262 27908
rect 9308 27862 9337 27908
rect 9233 27804 9337 27862
rect 9233 27758 9262 27804
rect 9308 27758 9337 27804
rect 9233 27745 9337 27758
rect 9457 28640 9561 28653
rect 9457 28594 9486 28640
rect 9532 28594 9561 28640
rect 9457 28535 9561 28594
rect 9457 28489 9486 28535
rect 9532 28489 9561 28535
rect 9457 28430 9561 28489
rect 9457 28384 9486 28430
rect 9532 28384 9561 28430
rect 9457 28325 9561 28384
rect 9457 28279 9486 28325
rect 9532 28279 9561 28325
rect 9457 28220 9561 28279
rect 9457 28174 9486 28220
rect 9532 28174 9561 28220
rect 9457 28116 9561 28174
rect 9457 28070 9486 28116
rect 9532 28070 9561 28116
rect 9457 28012 9561 28070
rect 9457 27966 9486 28012
rect 9532 27966 9561 28012
rect 9457 27908 9561 27966
rect 9457 27862 9486 27908
rect 9532 27862 9561 27908
rect 9457 27804 9561 27862
rect 9457 27758 9486 27804
rect 9532 27758 9561 27804
rect 9457 27745 9561 27758
rect 9681 28640 9785 28653
rect 9681 28594 9710 28640
rect 9756 28594 9785 28640
rect 9681 28535 9785 28594
rect 9681 28489 9710 28535
rect 9756 28489 9785 28535
rect 9681 28430 9785 28489
rect 9681 28384 9710 28430
rect 9756 28384 9785 28430
rect 9681 28325 9785 28384
rect 9681 28279 9710 28325
rect 9756 28279 9785 28325
rect 9681 28220 9785 28279
rect 9681 28174 9710 28220
rect 9756 28174 9785 28220
rect 9681 28116 9785 28174
rect 9681 28070 9710 28116
rect 9756 28070 9785 28116
rect 9681 28012 9785 28070
rect 9681 27966 9710 28012
rect 9756 27966 9785 28012
rect 9681 27908 9785 27966
rect 9681 27862 9710 27908
rect 9756 27862 9785 27908
rect 9681 27804 9785 27862
rect 9681 27758 9710 27804
rect 9756 27758 9785 27804
rect 9681 27745 9785 27758
rect 9905 28640 10009 28653
rect 9905 28594 9934 28640
rect 9980 28594 10009 28640
rect 9905 28535 10009 28594
rect 9905 28489 9934 28535
rect 9980 28489 10009 28535
rect 9905 28430 10009 28489
rect 9905 28384 9934 28430
rect 9980 28384 10009 28430
rect 9905 28325 10009 28384
rect 9905 28279 9934 28325
rect 9980 28279 10009 28325
rect 9905 28220 10009 28279
rect 9905 28174 9934 28220
rect 9980 28174 10009 28220
rect 9905 28116 10009 28174
rect 9905 28070 9934 28116
rect 9980 28070 10009 28116
rect 9905 28012 10009 28070
rect 9905 27966 9934 28012
rect 9980 27966 10009 28012
rect 9905 27908 10009 27966
rect 9905 27862 9934 27908
rect 9980 27862 10009 27908
rect 9905 27804 10009 27862
rect 9905 27758 9934 27804
rect 9980 27758 10009 27804
rect 9905 27745 10009 27758
rect 10129 28640 10233 28653
rect 10129 28594 10158 28640
rect 10204 28594 10233 28640
rect 10129 28535 10233 28594
rect 10129 28489 10158 28535
rect 10204 28489 10233 28535
rect 10129 28430 10233 28489
rect 10129 28384 10158 28430
rect 10204 28384 10233 28430
rect 10129 28325 10233 28384
rect 10129 28279 10158 28325
rect 10204 28279 10233 28325
rect 10129 28220 10233 28279
rect 10129 28174 10158 28220
rect 10204 28174 10233 28220
rect 10129 28116 10233 28174
rect 10129 28070 10158 28116
rect 10204 28070 10233 28116
rect 10129 28012 10233 28070
rect 10129 27966 10158 28012
rect 10204 27966 10233 28012
rect 10129 27908 10233 27966
rect 10129 27862 10158 27908
rect 10204 27862 10233 27908
rect 10129 27804 10233 27862
rect 10129 27758 10158 27804
rect 10204 27758 10233 27804
rect 10129 27745 10233 27758
rect 10353 28640 10457 28653
rect 10353 28594 10382 28640
rect 10428 28594 10457 28640
rect 10353 28535 10457 28594
rect 10353 28489 10382 28535
rect 10428 28489 10457 28535
rect 10353 28430 10457 28489
rect 10353 28384 10382 28430
rect 10428 28384 10457 28430
rect 10353 28325 10457 28384
rect 10353 28279 10382 28325
rect 10428 28279 10457 28325
rect 10353 28220 10457 28279
rect 10353 28174 10382 28220
rect 10428 28174 10457 28220
rect 10353 28116 10457 28174
rect 10353 28070 10382 28116
rect 10428 28070 10457 28116
rect 10353 28012 10457 28070
rect 10353 27966 10382 28012
rect 10428 27966 10457 28012
rect 10353 27908 10457 27966
rect 10353 27862 10382 27908
rect 10428 27862 10457 27908
rect 10353 27804 10457 27862
rect 10353 27758 10382 27804
rect 10428 27758 10457 27804
rect 10353 27745 10457 27758
rect 10577 28640 10681 28653
rect 10577 28594 10606 28640
rect 10652 28594 10681 28640
rect 10577 28535 10681 28594
rect 10577 28489 10606 28535
rect 10652 28489 10681 28535
rect 10577 28430 10681 28489
rect 10577 28384 10606 28430
rect 10652 28384 10681 28430
rect 10577 28325 10681 28384
rect 10577 28279 10606 28325
rect 10652 28279 10681 28325
rect 10577 28220 10681 28279
rect 10577 28174 10606 28220
rect 10652 28174 10681 28220
rect 10577 28116 10681 28174
rect 10577 28070 10606 28116
rect 10652 28070 10681 28116
rect 10577 28012 10681 28070
rect 10577 27966 10606 28012
rect 10652 27966 10681 28012
rect 10577 27908 10681 27966
rect 10577 27862 10606 27908
rect 10652 27862 10681 27908
rect 10577 27804 10681 27862
rect 10577 27758 10606 27804
rect 10652 27758 10681 27804
rect 10577 27745 10681 27758
rect 10801 28640 10905 28653
rect 10801 28594 10830 28640
rect 10876 28594 10905 28640
rect 10801 28535 10905 28594
rect 10801 28489 10830 28535
rect 10876 28489 10905 28535
rect 10801 28430 10905 28489
rect 10801 28384 10830 28430
rect 10876 28384 10905 28430
rect 10801 28325 10905 28384
rect 10801 28279 10830 28325
rect 10876 28279 10905 28325
rect 10801 28220 10905 28279
rect 10801 28174 10830 28220
rect 10876 28174 10905 28220
rect 10801 28116 10905 28174
rect 10801 28070 10830 28116
rect 10876 28070 10905 28116
rect 10801 28012 10905 28070
rect 10801 27966 10830 28012
rect 10876 27966 10905 28012
rect 10801 27908 10905 27966
rect 10801 27862 10830 27908
rect 10876 27862 10905 27908
rect 10801 27804 10905 27862
rect 10801 27758 10830 27804
rect 10876 27758 10905 27804
rect 10801 27745 10905 27758
rect 11025 28640 11129 28653
rect 11025 28594 11054 28640
rect 11100 28594 11129 28640
rect 11025 28535 11129 28594
rect 11025 28489 11054 28535
rect 11100 28489 11129 28535
rect 11025 28430 11129 28489
rect 11025 28384 11054 28430
rect 11100 28384 11129 28430
rect 11025 28325 11129 28384
rect 11025 28279 11054 28325
rect 11100 28279 11129 28325
rect 11025 28220 11129 28279
rect 11025 28174 11054 28220
rect 11100 28174 11129 28220
rect 11025 28116 11129 28174
rect 11025 28070 11054 28116
rect 11100 28070 11129 28116
rect 11025 28012 11129 28070
rect 11025 27966 11054 28012
rect 11100 27966 11129 28012
rect 11025 27908 11129 27966
rect 11025 27862 11054 27908
rect 11100 27862 11129 27908
rect 11025 27804 11129 27862
rect 11025 27758 11054 27804
rect 11100 27758 11129 27804
rect 11025 27745 11129 27758
rect 11249 28640 11353 28653
rect 11249 28594 11278 28640
rect 11324 28594 11353 28640
rect 11249 28535 11353 28594
rect 11249 28489 11278 28535
rect 11324 28489 11353 28535
rect 11249 28430 11353 28489
rect 11249 28384 11278 28430
rect 11324 28384 11353 28430
rect 11249 28325 11353 28384
rect 11249 28279 11278 28325
rect 11324 28279 11353 28325
rect 11249 28220 11353 28279
rect 11249 28174 11278 28220
rect 11324 28174 11353 28220
rect 11249 28116 11353 28174
rect 11249 28070 11278 28116
rect 11324 28070 11353 28116
rect 11249 28012 11353 28070
rect 11249 27966 11278 28012
rect 11324 27966 11353 28012
rect 11249 27908 11353 27966
rect 11249 27862 11278 27908
rect 11324 27862 11353 27908
rect 11249 27804 11353 27862
rect 11249 27758 11278 27804
rect 11324 27758 11353 27804
rect 11249 27745 11353 27758
rect 11473 28640 11577 28653
rect 11473 28594 11502 28640
rect 11548 28594 11577 28640
rect 11473 28535 11577 28594
rect 11473 28489 11502 28535
rect 11548 28489 11577 28535
rect 11473 28430 11577 28489
rect 11473 28384 11502 28430
rect 11548 28384 11577 28430
rect 11473 28325 11577 28384
rect 11473 28279 11502 28325
rect 11548 28279 11577 28325
rect 11473 28220 11577 28279
rect 11473 28174 11502 28220
rect 11548 28174 11577 28220
rect 11473 28116 11577 28174
rect 11473 28070 11502 28116
rect 11548 28070 11577 28116
rect 11473 28012 11577 28070
rect 11473 27966 11502 28012
rect 11548 27966 11577 28012
rect 11473 27908 11577 27966
rect 11473 27862 11502 27908
rect 11548 27862 11577 27908
rect 11473 27804 11577 27862
rect 11473 27758 11502 27804
rect 11548 27758 11577 27804
rect 11473 27745 11577 27758
rect 11697 28640 11801 28653
rect 11697 28594 11726 28640
rect 11772 28594 11801 28640
rect 11697 28535 11801 28594
rect 11697 28489 11726 28535
rect 11772 28489 11801 28535
rect 11697 28430 11801 28489
rect 11697 28384 11726 28430
rect 11772 28384 11801 28430
rect 11697 28325 11801 28384
rect 11697 28279 11726 28325
rect 11772 28279 11801 28325
rect 11697 28220 11801 28279
rect 11697 28174 11726 28220
rect 11772 28174 11801 28220
rect 11697 28116 11801 28174
rect 11697 28070 11726 28116
rect 11772 28070 11801 28116
rect 11697 28012 11801 28070
rect 11697 27966 11726 28012
rect 11772 27966 11801 28012
rect 11697 27908 11801 27966
rect 11697 27862 11726 27908
rect 11772 27862 11801 27908
rect 11697 27804 11801 27862
rect 11697 27758 11726 27804
rect 11772 27758 11801 27804
rect 11697 27745 11801 27758
rect 11921 28640 12025 28653
rect 11921 28594 11950 28640
rect 11996 28594 12025 28640
rect 11921 28535 12025 28594
rect 11921 28489 11950 28535
rect 11996 28489 12025 28535
rect 11921 28430 12025 28489
rect 11921 28384 11950 28430
rect 11996 28384 12025 28430
rect 11921 28325 12025 28384
rect 11921 28279 11950 28325
rect 11996 28279 12025 28325
rect 11921 28220 12025 28279
rect 11921 28174 11950 28220
rect 11996 28174 12025 28220
rect 11921 28116 12025 28174
rect 11921 28070 11950 28116
rect 11996 28070 12025 28116
rect 11921 28012 12025 28070
rect 11921 27966 11950 28012
rect 11996 27966 12025 28012
rect 11921 27908 12025 27966
rect 11921 27862 11950 27908
rect 11996 27862 12025 27908
rect 11921 27804 12025 27862
rect 11921 27758 11950 27804
rect 11996 27758 12025 27804
rect 11921 27745 12025 27758
rect 12145 28640 12249 28653
rect 12145 28594 12174 28640
rect 12220 28594 12249 28640
rect 12145 28535 12249 28594
rect 12145 28489 12174 28535
rect 12220 28489 12249 28535
rect 12145 28430 12249 28489
rect 12145 28384 12174 28430
rect 12220 28384 12249 28430
rect 12145 28325 12249 28384
rect 12145 28279 12174 28325
rect 12220 28279 12249 28325
rect 12145 28220 12249 28279
rect 12145 28174 12174 28220
rect 12220 28174 12249 28220
rect 12145 28116 12249 28174
rect 12145 28070 12174 28116
rect 12220 28070 12249 28116
rect 12145 28012 12249 28070
rect 12145 27966 12174 28012
rect 12220 27966 12249 28012
rect 12145 27908 12249 27966
rect 12145 27862 12174 27908
rect 12220 27862 12249 27908
rect 12145 27804 12249 27862
rect 12145 27758 12174 27804
rect 12220 27758 12249 27804
rect 12145 27745 12249 27758
rect 12369 28640 12473 28653
rect 12369 28594 12398 28640
rect 12444 28594 12473 28640
rect 12369 28535 12473 28594
rect 12369 28489 12398 28535
rect 12444 28489 12473 28535
rect 12369 28430 12473 28489
rect 12369 28384 12398 28430
rect 12444 28384 12473 28430
rect 12369 28325 12473 28384
rect 12369 28279 12398 28325
rect 12444 28279 12473 28325
rect 12369 28220 12473 28279
rect 12369 28174 12398 28220
rect 12444 28174 12473 28220
rect 12369 28116 12473 28174
rect 12369 28070 12398 28116
rect 12444 28070 12473 28116
rect 12369 28012 12473 28070
rect 12369 27966 12398 28012
rect 12444 27966 12473 28012
rect 12369 27908 12473 27966
rect 12369 27862 12398 27908
rect 12444 27862 12473 27908
rect 12369 27804 12473 27862
rect 12369 27758 12398 27804
rect 12444 27758 12473 27804
rect 12369 27745 12473 27758
rect 12593 28640 12681 28653
rect 12593 28594 12622 28640
rect 12668 28594 12681 28640
rect 12593 28535 12681 28594
rect 12593 28489 12622 28535
rect 12668 28489 12681 28535
rect 12593 28430 12681 28489
rect 12593 28384 12622 28430
rect 12668 28384 12681 28430
rect 12593 28325 12681 28384
rect 12593 28279 12622 28325
rect 12668 28279 12681 28325
rect 12593 28220 12681 28279
rect 12593 28174 12622 28220
rect 12668 28174 12681 28220
rect 12593 28116 12681 28174
rect 23784 28190 23872 28203
rect 12593 28070 12622 28116
rect 12668 28070 12681 28116
rect 23784 28144 23797 28190
rect 23843 28144 23872 28190
rect 12593 28012 12681 28070
rect 12593 27966 12622 28012
rect 12668 27966 12681 28012
rect 12593 27908 12681 27966
rect 12593 27862 12622 27908
rect 12668 27862 12681 27908
rect 12593 27804 12681 27862
rect 13299 28082 13387 28095
rect 13299 27834 13312 28082
rect 13358 27834 13387 28082
rect 13299 27821 13387 27834
rect 13507 28082 13611 28095
rect 13507 27834 13536 28082
rect 13582 27834 13611 28082
rect 13507 27821 13611 27834
rect 13731 28082 13819 28095
rect 13731 27834 13760 28082
rect 13806 27834 13819 28082
rect 13731 27821 13819 27834
rect 16691 28076 16779 28089
rect 16691 28030 16704 28076
rect 16750 28030 16779 28076
rect 12593 27758 12622 27804
rect 12668 27758 12681 27804
rect 12593 27745 12681 27758
rect 14893 27996 14981 28009
rect 14893 27950 14906 27996
rect 14952 27950 14981 27996
rect 14893 27876 14981 27950
rect 14893 27830 14906 27876
rect 14952 27830 14981 27876
rect 14893 27817 14981 27830
rect 15101 27996 15189 28009
rect 15101 27950 15130 27996
rect 15176 27950 15189 27996
rect 15101 27876 15189 27950
rect 15101 27830 15130 27876
rect 15176 27830 15189 27876
rect 15101 27817 15189 27830
rect 16691 27971 16779 28030
rect 16691 27925 16704 27971
rect 16750 27925 16779 27971
rect 16691 27866 16779 27925
rect 16691 27820 16704 27866
rect 16750 27820 16779 27866
rect 6078 26731 6166 26744
rect 6078 26379 6091 26731
rect 6137 26379 6166 26731
rect 6078 26322 6166 26379
rect 6078 26276 6091 26322
rect 6137 26276 6166 26322
rect 6078 26219 6166 26276
rect 6078 26173 6091 26219
rect 6137 26173 6166 26219
rect 6078 26116 6166 26173
rect 6078 26070 6091 26116
rect 6137 26070 6166 26116
rect 6078 26013 6166 26070
rect 6078 25967 6091 26013
rect 6137 25967 6166 26013
rect 6078 25910 6166 25967
rect 6078 25864 6091 25910
rect 6137 25864 6166 25910
rect 6078 25807 6166 25864
rect 6078 25761 6091 25807
rect 6137 25761 6166 25807
rect 6078 25704 6166 25761
rect 6078 25658 6091 25704
rect 6137 25658 6166 25704
rect 6078 25601 6166 25658
rect 6078 25555 6091 25601
rect 6137 25555 6166 25601
rect 6078 25498 6166 25555
rect 6078 25452 6091 25498
rect 6137 25452 6166 25498
rect 6078 25395 6166 25452
rect 6078 25349 6091 25395
rect 6137 25349 6166 25395
rect 6078 25336 6166 25349
rect 6286 26731 6374 26744
rect 6286 26379 6315 26731
rect 6361 26379 6374 26731
rect 7769 26731 7857 26744
rect 6286 26322 6374 26379
rect 6286 26276 6315 26322
rect 6361 26276 6374 26322
rect 6286 26219 6374 26276
rect 6286 26173 6315 26219
rect 6361 26173 6374 26219
rect 6286 26116 6374 26173
rect 6286 26070 6315 26116
rect 6361 26070 6374 26116
rect 6286 26013 6374 26070
rect 6286 25967 6315 26013
rect 6361 25967 6374 26013
rect 6286 25910 6374 25967
rect 6286 25864 6315 25910
rect 6361 25864 6374 25910
rect 6286 25807 6374 25864
rect 6286 25761 6315 25807
rect 6361 25761 6374 25807
rect 6286 25704 6374 25761
rect 6286 25658 6315 25704
rect 6361 25658 6374 25704
rect 6286 25601 6374 25658
rect 6286 25555 6315 25601
rect 6361 25555 6374 25601
rect 6286 25498 6374 25555
rect 6286 25452 6315 25498
rect 6361 25452 6374 25498
rect 6286 25395 6374 25452
rect 6592 26446 6680 26459
rect 6592 26400 6605 26446
rect 6651 26400 6680 26446
rect 6592 26338 6680 26400
rect 6592 26292 6605 26338
rect 6651 26292 6680 26338
rect 6592 26230 6680 26292
rect 6592 26184 6605 26230
rect 6651 26184 6680 26230
rect 6592 26122 6680 26184
rect 6592 26076 6605 26122
rect 6651 26076 6680 26122
rect 6592 26014 6680 26076
rect 6592 25968 6605 26014
rect 6651 25968 6680 26014
rect 6592 25906 6680 25968
rect 6592 25860 6605 25906
rect 6651 25860 6680 25906
rect 6592 25798 6680 25860
rect 6592 25752 6605 25798
rect 6651 25752 6680 25798
rect 6592 25690 6680 25752
rect 6592 25644 6605 25690
rect 6651 25644 6680 25690
rect 6592 25582 6680 25644
rect 6592 25536 6605 25582
rect 6651 25536 6680 25582
rect 6592 25474 6680 25536
rect 6592 25428 6605 25474
rect 6651 25428 6680 25474
rect 6592 25415 6680 25428
rect 6800 26446 6888 26459
rect 6800 26400 6829 26446
rect 6875 26400 6888 26446
rect 6800 26338 6888 26400
rect 6800 26292 6829 26338
rect 6875 26292 6888 26338
rect 6800 26230 6888 26292
rect 6800 26184 6829 26230
rect 6875 26184 6888 26230
rect 6800 26122 6888 26184
rect 6800 26076 6829 26122
rect 6875 26076 6888 26122
rect 6800 26014 6888 26076
rect 6800 25968 6829 26014
rect 6875 25968 6888 26014
rect 6800 25906 6888 25968
rect 6800 25860 6829 25906
rect 6875 25860 6888 25906
rect 6800 25798 6888 25860
rect 6800 25752 6829 25798
rect 6875 25752 6888 25798
rect 6800 25690 6888 25752
rect 6800 25644 6829 25690
rect 6875 25644 6888 25690
rect 6800 25582 6888 25644
rect 6800 25536 6829 25582
rect 6875 25536 6888 25582
rect 6800 25474 6888 25536
rect 6800 25428 6829 25474
rect 6875 25428 6888 25474
rect 7769 26379 7782 26731
rect 7828 26379 7857 26731
rect 7769 26322 7857 26379
rect 7769 26276 7782 26322
rect 7828 26276 7857 26322
rect 7769 26219 7857 26276
rect 7769 26173 7782 26219
rect 7828 26173 7857 26219
rect 7769 26116 7857 26173
rect 7769 26070 7782 26116
rect 7828 26070 7857 26116
rect 7769 26013 7857 26070
rect 7769 25967 7782 26013
rect 7828 25967 7857 26013
rect 7769 25910 7857 25967
rect 7769 25864 7782 25910
rect 7828 25864 7857 25910
rect 7769 25807 7857 25864
rect 7769 25761 7782 25807
rect 7828 25761 7857 25807
rect 7769 25704 7857 25761
rect 7769 25658 7782 25704
rect 7828 25658 7857 25704
rect 7769 25601 7857 25658
rect 7769 25555 7782 25601
rect 7828 25555 7857 25601
rect 7769 25498 7857 25555
rect 6800 25415 6888 25428
rect 7769 25452 7782 25498
rect 7828 25452 7857 25498
rect 6286 25349 6315 25395
rect 6361 25349 6374 25395
rect 6286 25336 6374 25349
rect 7769 25395 7857 25452
rect 7769 25349 7782 25395
rect 7828 25349 7857 25395
rect 7769 25336 7857 25349
rect 7977 26731 8065 26744
rect 7977 26379 8006 26731
rect 8052 26379 8065 26731
rect 7977 26322 8065 26379
rect 7977 26276 8006 26322
rect 8052 26276 8065 26322
rect 7977 26219 8065 26276
rect 7977 26173 8006 26219
rect 8052 26173 8065 26219
rect 7977 26116 8065 26173
rect 7977 26070 8006 26116
rect 8052 26070 8065 26116
rect 7977 26013 8065 26070
rect 7977 25967 8006 26013
rect 8052 25967 8065 26013
rect 7977 25910 8065 25967
rect 7977 25864 8006 25910
rect 8052 25864 8065 25910
rect 7977 25807 8065 25864
rect 7977 25761 8006 25807
rect 8052 25761 8065 25807
rect 7977 25704 8065 25761
rect 7977 25658 8006 25704
rect 8052 25658 8065 25704
rect 7977 25601 8065 25658
rect 7977 25555 8006 25601
rect 8052 25555 8065 25601
rect 7977 25498 8065 25555
rect 7977 25452 8006 25498
rect 8052 25452 8065 25498
rect 7977 25395 8065 25452
rect 8283 26446 8371 26459
rect 8283 26400 8296 26446
rect 8342 26400 8371 26446
rect 8283 26338 8371 26400
rect 8283 26292 8296 26338
rect 8342 26292 8371 26338
rect 8283 26230 8371 26292
rect 8283 26184 8296 26230
rect 8342 26184 8371 26230
rect 8283 26122 8371 26184
rect 8283 26076 8296 26122
rect 8342 26076 8371 26122
rect 8283 26014 8371 26076
rect 8283 25968 8296 26014
rect 8342 25968 8371 26014
rect 8283 25906 8371 25968
rect 8283 25860 8296 25906
rect 8342 25860 8371 25906
rect 8283 25798 8371 25860
rect 8283 25752 8296 25798
rect 8342 25752 8371 25798
rect 8283 25690 8371 25752
rect 8283 25644 8296 25690
rect 8342 25644 8371 25690
rect 8283 25582 8371 25644
rect 8283 25536 8296 25582
rect 8342 25536 8371 25582
rect 8283 25474 8371 25536
rect 8283 25428 8296 25474
rect 8342 25428 8371 25474
rect 8283 25415 8371 25428
rect 8491 26446 8579 26459
rect 8491 26400 8520 26446
rect 8566 26400 8579 26446
rect 8491 26338 8579 26400
rect 8491 26292 8520 26338
rect 8566 26292 8579 26338
rect 8491 26230 8579 26292
rect 8491 26184 8520 26230
rect 8566 26184 8579 26230
rect 8491 26122 8579 26184
rect 8491 26076 8520 26122
rect 8566 26076 8579 26122
rect 8491 26014 8579 26076
rect 8491 25968 8520 26014
rect 8566 25968 8579 26014
rect 8491 25906 8579 25968
rect 8491 25860 8520 25906
rect 8566 25860 8579 25906
rect 8491 25798 8579 25860
rect 8491 25752 8520 25798
rect 8566 25752 8579 25798
rect 8491 25690 8579 25752
rect 8491 25644 8520 25690
rect 8566 25644 8579 25690
rect 8491 25582 8579 25644
rect 8491 25536 8520 25582
rect 8566 25536 8579 25582
rect 8491 25474 8579 25536
rect 8491 25428 8520 25474
rect 8566 25428 8579 25474
rect 8491 25415 8579 25428
rect 7977 25349 8006 25395
rect 8052 25349 8065 25395
rect 7977 25336 8065 25349
rect 16691 27761 16779 27820
rect 16691 27715 16704 27761
rect 16750 27715 16779 27761
rect 16691 27656 16779 27715
rect 16691 27610 16704 27656
rect 16750 27610 16779 27656
rect 16691 27552 16779 27610
rect 16691 27506 16704 27552
rect 16750 27506 16779 27552
rect 16691 27448 16779 27506
rect 16691 27402 16704 27448
rect 16750 27402 16779 27448
rect 16691 27344 16779 27402
rect 16691 27298 16704 27344
rect 16750 27298 16779 27344
rect 16691 27240 16779 27298
rect 16691 27194 16704 27240
rect 16750 27194 16779 27240
rect 16691 27181 16779 27194
rect 16899 28076 17003 28089
rect 16899 28030 16928 28076
rect 16974 28030 17003 28076
rect 16899 27971 17003 28030
rect 16899 27925 16928 27971
rect 16974 27925 17003 27971
rect 16899 27866 17003 27925
rect 16899 27820 16928 27866
rect 16974 27820 17003 27866
rect 16899 27761 17003 27820
rect 16899 27715 16928 27761
rect 16974 27715 17003 27761
rect 16899 27656 17003 27715
rect 16899 27610 16928 27656
rect 16974 27610 17003 27656
rect 16899 27552 17003 27610
rect 16899 27506 16928 27552
rect 16974 27506 17003 27552
rect 16899 27448 17003 27506
rect 16899 27402 16928 27448
rect 16974 27402 17003 27448
rect 16899 27344 17003 27402
rect 16899 27298 16928 27344
rect 16974 27298 17003 27344
rect 16899 27240 17003 27298
rect 16899 27194 16928 27240
rect 16974 27194 17003 27240
rect 16899 27181 17003 27194
rect 17123 28076 17227 28089
rect 17123 28030 17152 28076
rect 17198 28030 17227 28076
rect 17123 27971 17227 28030
rect 17123 27925 17152 27971
rect 17198 27925 17227 27971
rect 17123 27866 17227 27925
rect 17123 27820 17152 27866
rect 17198 27820 17227 27866
rect 17123 27761 17227 27820
rect 17123 27715 17152 27761
rect 17198 27715 17227 27761
rect 17123 27656 17227 27715
rect 17123 27610 17152 27656
rect 17198 27610 17227 27656
rect 17123 27552 17227 27610
rect 17123 27506 17152 27552
rect 17198 27506 17227 27552
rect 17123 27448 17227 27506
rect 17123 27402 17152 27448
rect 17198 27402 17227 27448
rect 17123 27344 17227 27402
rect 17123 27298 17152 27344
rect 17198 27298 17227 27344
rect 17123 27240 17227 27298
rect 17123 27194 17152 27240
rect 17198 27194 17227 27240
rect 17123 27181 17227 27194
rect 17347 28076 17451 28089
rect 17347 28030 17376 28076
rect 17422 28030 17451 28076
rect 17347 27971 17451 28030
rect 17347 27925 17376 27971
rect 17422 27925 17451 27971
rect 17347 27866 17451 27925
rect 17347 27820 17376 27866
rect 17422 27820 17451 27866
rect 17347 27761 17451 27820
rect 17347 27715 17376 27761
rect 17422 27715 17451 27761
rect 17347 27656 17451 27715
rect 17347 27610 17376 27656
rect 17422 27610 17451 27656
rect 17347 27552 17451 27610
rect 17347 27506 17376 27552
rect 17422 27506 17451 27552
rect 17347 27448 17451 27506
rect 17347 27402 17376 27448
rect 17422 27402 17451 27448
rect 17347 27344 17451 27402
rect 17347 27298 17376 27344
rect 17422 27298 17451 27344
rect 17347 27240 17451 27298
rect 17347 27194 17376 27240
rect 17422 27194 17451 27240
rect 17347 27181 17451 27194
rect 17571 28076 17675 28089
rect 17571 28030 17600 28076
rect 17646 28030 17675 28076
rect 17571 27971 17675 28030
rect 17571 27925 17600 27971
rect 17646 27925 17675 27971
rect 17571 27866 17675 27925
rect 17571 27820 17600 27866
rect 17646 27820 17675 27866
rect 17571 27761 17675 27820
rect 17571 27715 17600 27761
rect 17646 27715 17675 27761
rect 17571 27656 17675 27715
rect 17571 27610 17600 27656
rect 17646 27610 17675 27656
rect 17571 27552 17675 27610
rect 17571 27506 17600 27552
rect 17646 27506 17675 27552
rect 17571 27448 17675 27506
rect 17571 27402 17600 27448
rect 17646 27402 17675 27448
rect 17571 27344 17675 27402
rect 17571 27298 17600 27344
rect 17646 27298 17675 27344
rect 17571 27240 17675 27298
rect 17571 27194 17600 27240
rect 17646 27194 17675 27240
rect 17571 27181 17675 27194
rect 17795 28076 17899 28089
rect 17795 28030 17824 28076
rect 17870 28030 17899 28076
rect 17795 27971 17899 28030
rect 17795 27925 17824 27971
rect 17870 27925 17899 27971
rect 17795 27866 17899 27925
rect 17795 27820 17824 27866
rect 17870 27820 17899 27866
rect 17795 27761 17899 27820
rect 17795 27715 17824 27761
rect 17870 27715 17899 27761
rect 17795 27656 17899 27715
rect 17795 27610 17824 27656
rect 17870 27610 17899 27656
rect 17795 27552 17899 27610
rect 17795 27506 17824 27552
rect 17870 27506 17899 27552
rect 17795 27448 17899 27506
rect 17795 27402 17824 27448
rect 17870 27402 17899 27448
rect 17795 27344 17899 27402
rect 17795 27298 17824 27344
rect 17870 27298 17899 27344
rect 17795 27240 17899 27298
rect 17795 27194 17824 27240
rect 17870 27194 17899 27240
rect 17795 27181 17899 27194
rect 18019 28076 18107 28089
rect 18019 28030 18048 28076
rect 18094 28030 18107 28076
rect 18019 27971 18107 28030
rect 18019 27925 18048 27971
rect 18094 27925 18107 27971
rect 18019 27866 18107 27925
rect 18019 27820 18048 27866
rect 18094 27820 18107 27866
rect 18019 27761 18107 27820
rect 18019 27715 18048 27761
rect 18094 27715 18107 27761
rect 18019 27656 18107 27715
rect 18019 27610 18048 27656
rect 18094 27610 18107 27656
rect 18019 27552 18107 27610
rect 18019 27506 18048 27552
rect 18094 27506 18107 27552
rect 18019 27448 18107 27506
rect 18019 27402 18048 27448
rect 18094 27402 18107 27448
rect 18019 27344 18107 27402
rect 18019 27298 18048 27344
rect 18094 27298 18107 27344
rect 18019 27240 18107 27298
rect 18019 27194 18048 27240
rect 18094 27194 18107 27240
rect 18019 27181 18107 27194
rect 18325 28076 18413 28089
rect 18325 28030 18338 28076
rect 18384 28030 18413 28076
rect 18325 27971 18413 28030
rect 18325 27925 18338 27971
rect 18384 27925 18413 27971
rect 18325 27866 18413 27925
rect 18325 27820 18338 27866
rect 18384 27820 18413 27866
rect 18325 27761 18413 27820
rect 18325 27715 18338 27761
rect 18384 27715 18413 27761
rect 18325 27656 18413 27715
rect 18325 27610 18338 27656
rect 18384 27610 18413 27656
rect 18325 27552 18413 27610
rect 18325 27506 18338 27552
rect 18384 27506 18413 27552
rect 18325 27448 18413 27506
rect 18325 27402 18338 27448
rect 18384 27402 18413 27448
rect 18325 27344 18413 27402
rect 18325 27298 18338 27344
rect 18384 27298 18413 27344
rect 18325 27240 18413 27298
rect 18325 27194 18338 27240
rect 18384 27194 18413 27240
rect 18325 27181 18413 27194
rect 18533 28076 18637 28089
rect 18533 28030 18562 28076
rect 18608 28030 18637 28076
rect 18533 27971 18637 28030
rect 18533 27925 18562 27971
rect 18608 27925 18637 27971
rect 18533 27866 18637 27925
rect 18533 27820 18562 27866
rect 18608 27820 18637 27866
rect 18533 27761 18637 27820
rect 18533 27715 18562 27761
rect 18608 27715 18637 27761
rect 18533 27656 18637 27715
rect 18533 27610 18562 27656
rect 18608 27610 18637 27656
rect 18533 27552 18637 27610
rect 18533 27506 18562 27552
rect 18608 27506 18637 27552
rect 18533 27448 18637 27506
rect 18533 27402 18562 27448
rect 18608 27402 18637 27448
rect 18533 27344 18637 27402
rect 18533 27298 18562 27344
rect 18608 27298 18637 27344
rect 18533 27240 18637 27298
rect 18533 27194 18562 27240
rect 18608 27194 18637 27240
rect 18533 27181 18637 27194
rect 18757 28076 18861 28089
rect 18757 28030 18786 28076
rect 18832 28030 18861 28076
rect 18757 27971 18861 28030
rect 18757 27925 18786 27971
rect 18832 27925 18861 27971
rect 18757 27866 18861 27925
rect 18757 27820 18786 27866
rect 18832 27820 18861 27866
rect 18757 27761 18861 27820
rect 18757 27715 18786 27761
rect 18832 27715 18861 27761
rect 18757 27656 18861 27715
rect 18757 27610 18786 27656
rect 18832 27610 18861 27656
rect 18757 27552 18861 27610
rect 18757 27506 18786 27552
rect 18832 27506 18861 27552
rect 18757 27448 18861 27506
rect 18757 27402 18786 27448
rect 18832 27402 18861 27448
rect 18757 27344 18861 27402
rect 18757 27298 18786 27344
rect 18832 27298 18861 27344
rect 18757 27240 18861 27298
rect 18757 27194 18786 27240
rect 18832 27194 18861 27240
rect 18757 27181 18861 27194
rect 18981 28076 19085 28089
rect 18981 28030 19010 28076
rect 19056 28030 19085 28076
rect 18981 27971 19085 28030
rect 18981 27925 19010 27971
rect 19056 27925 19085 27971
rect 18981 27866 19085 27925
rect 18981 27820 19010 27866
rect 19056 27820 19085 27866
rect 18981 27761 19085 27820
rect 18981 27715 19010 27761
rect 19056 27715 19085 27761
rect 18981 27656 19085 27715
rect 18981 27610 19010 27656
rect 19056 27610 19085 27656
rect 18981 27552 19085 27610
rect 18981 27506 19010 27552
rect 19056 27506 19085 27552
rect 18981 27448 19085 27506
rect 18981 27402 19010 27448
rect 19056 27402 19085 27448
rect 18981 27344 19085 27402
rect 18981 27298 19010 27344
rect 19056 27298 19085 27344
rect 18981 27240 19085 27298
rect 18981 27194 19010 27240
rect 19056 27194 19085 27240
rect 18981 27181 19085 27194
rect 19205 28076 19309 28089
rect 19205 28030 19234 28076
rect 19280 28030 19309 28076
rect 19205 27971 19309 28030
rect 19205 27925 19234 27971
rect 19280 27925 19309 27971
rect 19205 27866 19309 27925
rect 19205 27820 19234 27866
rect 19280 27820 19309 27866
rect 19205 27761 19309 27820
rect 19205 27715 19234 27761
rect 19280 27715 19309 27761
rect 19205 27656 19309 27715
rect 19205 27610 19234 27656
rect 19280 27610 19309 27656
rect 19205 27552 19309 27610
rect 19205 27506 19234 27552
rect 19280 27506 19309 27552
rect 19205 27448 19309 27506
rect 19205 27402 19234 27448
rect 19280 27402 19309 27448
rect 19205 27344 19309 27402
rect 19205 27298 19234 27344
rect 19280 27298 19309 27344
rect 19205 27240 19309 27298
rect 19205 27194 19234 27240
rect 19280 27194 19309 27240
rect 19205 27181 19309 27194
rect 19429 28076 19533 28089
rect 19429 28030 19458 28076
rect 19504 28030 19533 28076
rect 19429 27971 19533 28030
rect 19429 27925 19458 27971
rect 19504 27925 19533 27971
rect 19429 27866 19533 27925
rect 19429 27820 19458 27866
rect 19504 27820 19533 27866
rect 19429 27761 19533 27820
rect 19429 27715 19458 27761
rect 19504 27715 19533 27761
rect 19429 27656 19533 27715
rect 19429 27610 19458 27656
rect 19504 27610 19533 27656
rect 19429 27552 19533 27610
rect 19429 27506 19458 27552
rect 19504 27506 19533 27552
rect 19429 27448 19533 27506
rect 19429 27402 19458 27448
rect 19504 27402 19533 27448
rect 19429 27344 19533 27402
rect 19429 27298 19458 27344
rect 19504 27298 19533 27344
rect 19429 27240 19533 27298
rect 19429 27194 19458 27240
rect 19504 27194 19533 27240
rect 19429 27181 19533 27194
rect 19653 28076 19741 28089
rect 19653 28030 19682 28076
rect 19728 28030 19741 28076
rect 19653 27971 19741 28030
rect 19653 27925 19682 27971
rect 19728 27925 19741 27971
rect 19653 27866 19741 27925
rect 19653 27820 19682 27866
rect 19728 27820 19741 27866
rect 19653 27761 19741 27820
rect 19653 27715 19682 27761
rect 19728 27715 19741 27761
rect 19653 27656 19741 27715
rect 19653 27610 19682 27656
rect 19728 27610 19741 27656
rect 19653 27552 19741 27610
rect 19653 27506 19682 27552
rect 19728 27506 19741 27552
rect 19653 27448 19741 27506
rect 19653 27402 19682 27448
rect 19728 27402 19741 27448
rect 19653 27344 19741 27402
rect 19653 27298 19682 27344
rect 19728 27298 19741 27344
rect 19653 27240 19741 27298
rect 19653 27194 19682 27240
rect 19728 27194 19741 27240
rect 19653 27181 19741 27194
rect 19958 28076 20046 28089
rect 19958 28030 19971 28076
rect 20017 28030 20046 28076
rect 19958 27971 20046 28030
rect 19958 27925 19971 27971
rect 20017 27925 20046 27971
rect 19958 27866 20046 27925
rect 19958 27820 19971 27866
rect 20017 27820 20046 27866
rect 19958 27761 20046 27820
rect 19958 27715 19971 27761
rect 20017 27715 20046 27761
rect 19958 27656 20046 27715
rect 19958 27610 19971 27656
rect 20017 27610 20046 27656
rect 19958 27552 20046 27610
rect 19958 27506 19971 27552
rect 20017 27506 20046 27552
rect 19958 27448 20046 27506
rect 19958 27402 19971 27448
rect 20017 27402 20046 27448
rect 19958 27344 20046 27402
rect 19958 27298 19971 27344
rect 20017 27298 20046 27344
rect 19958 27240 20046 27298
rect 19958 27194 19971 27240
rect 20017 27194 20046 27240
rect 19958 27181 20046 27194
rect 20166 28076 20270 28089
rect 20166 28030 20195 28076
rect 20241 28030 20270 28076
rect 20166 27971 20270 28030
rect 20166 27925 20195 27971
rect 20241 27925 20270 27971
rect 20166 27866 20270 27925
rect 20166 27820 20195 27866
rect 20241 27820 20270 27866
rect 20166 27761 20270 27820
rect 20166 27715 20195 27761
rect 20241 27715 20270 27761
rect 20166 27656 20270 27715
rect 20166 27610 20195 27656
rect 20241 27610 20270 27656
rect 20166 27552 20270 27610
rect 20166 27506 20195 27552
rect 20241 27506 20270 27552
rect 20166 27448 20270 27506
rect 20166 27402 20195 27448
rect 20241 27402 20270 27448
rect 20166 27344 20270 27402
rect 20166 27298 20195 27344
rect 20241 27298 20270 27344
rect 20166 27240 20270 27298
rect 20166 27194 20195 27240
rect 20241 27194 20270 27240
rect 20166 27181 20270 27194
rect 20390 28076 20494 28089
rect 20390 28030 20419 28076
rect 20465 28030 20494 28076
rect 20390 27971 20494 28030
rect 20390 27925 20419 27971
rect 20465 27925 20494 27971
rect 20390 27866 20494 27925
rect 20390 27820 20419 27866
rect 20465 27820 20494 27866
rect 20390 27761 20494 27820
rect 20390 27715 20419 27761
rect 20465 27715 20494 27761
rect 20390 27656 20494 27715
rect 20390 27610 20419 27656
rect 20465 27610 20494 27656
rect 20390 27552 20494 27610
rect 20390 27506 20419 27552
rect 20465 27506 20494 27552
rect 20390 27448 20494 27506
rect 20390 27402 20419 27448
rect 20465 27402 20494 27448
rect 20390 27344 20494 27402
rect 20390 27298 20419 27344
rect 20465 27298 20494 27344
rect 20390 27240 20494 27298
rect 20390 27194 20419 27240
rect 20465 27194 20494 27240
rect 20390 27181 20494 27194
rect 20614 28076 20718 28089
rect 20614 28030 20643 28076
rect 20689 28030 20718 28076
rect 20614 27971 20718 28030
rect 20614 27925 20643 27971
rect 20689 27925 20718 27971
rect 20614 27866 20718 27925
rect 20614 27820 20643 27866
rect 20689 27820 20718 27866
rect 20614 27761 20718 27820
rect 20614 27715 20643 27761
rect 20689 27715 20718 27761
rect 20614 27656 20718 27715
rect 20614 27610 20643 27656
rect 20689 27610 20718 27656
rect 20614 27552 20718 27610
rect 20614 27506 20643 27552
rect 20689 27506 20718 27552
rect 20614 27448 20718 27506
rect 20614 27402 20643 27448
rect 20689 27402 20718 27448
rect 20614 27344 20718 27402
rect 20614 27298 20643 27344
rect 20689 27298 20718 27344
rect 20614 27240 20718 27298
rect 20614 27194 20643 27240
rect 20689 27194 20718 27240
rect 20614 27181 20718 27194
rect 20838 28076 20942 28089
rect 20838 28030 20867 28076
rect 20913 28030 20942 28076
rect 20838 27971 20942 28030
rect 20838 27925 20867 27971
rect 20913 27925 20942 27971
rect 20838 27866 20942 27925
rect 20838 27820 20867 27866
rect 20913 27820 20942 27866
rect 20838 27761 20942 27820
rect 20838 27715 20867 27761
rect 20913 27715 20942 27761
rect 20838 27656 20942 27715
rect 20838 27610 20867 27656
rect 20913 27610 20942 27656
rect 20838 27552 20942 27610
rect 20838 27506 20867 27552
rect 20913 27506 20942 27552
rect 20838 27448 20942 27506
rect 20838 27402 20867 27448
rect 20913 27402 20942 27448
rect 20838 27344 20942 27402
rect 20838 27298 20867 27344
rect 20913 27298 20942 27344
rect 20838 27240 20942 27298
rect 20838 27194 20867 27240
rect 20913 27194 20942 27240
rect 20838 27181 20942 27194
rect 21062 28076 21166 28089
rect 21062 28030 21091 28076
rect 21137 28030 21166 28076
rect 21062 27971 21166 28030
rect 21062 27925 21091 27971
rect 21137 27925 21166 27971
rect 21062 27866 21166 27925
rect 21062 27820 21091 27866
rect 21137 27820 21166 27866
rect 21062 27761 21166 27820
rect 21062 27715 21091 27761
rect 21137 27715 21166 27761
rect 21062 27656 21166 27715
rect 21062 27610 21091 27656
rect 21137 27610 21166 27656
rect 21062 27552 21166 27610
rect 21062 27506 21091 27552
rect 21137 27506 21166 27552
rect 21062 27448 21166 27506
rect 21062 27402 21091 27448
rect 21137 27402 21166 27448
rect 21062 27344 21166 27402
rect 21062 27298 21091 27344
rect 21137 27298 21166 27344
rect 21062 27240 21166 27298
rect 21062 27194 21091 27240
rect 21137 27194 21166 27240
rect 21062 27181 21166 27194
rect 21286 28076 21374 28089
rect 21286 28030 21315 28076
rect 21361 28030 21374 28076
rect 21286 27971 21374 28030
rect 21286 27925 21315 27971
rect 21361 27925 21374 27971
rect 21286 27866 21374 27925
rect 21286 27820 21315 27866
rect 21361 27820 21374 27866
rect 21286 27761 21374 27820
rect 21286 27715 21315 27761
rect 21361 27715 21374 27761
rect 21286 27656 21374 27715
rect 21286 27610 21315 27656
rect 21361 27610 21374 27656
rect 21286 27552 21374 27610
rect 21286 27506 21315 27552
rect 21361 27506 21374 27552
rect 21286 27448 21374 27506
rect 21286 27402 21315 27448
rect 21361 27402 21374 27448
rect 21286 27344 21374 27402
rect 21286 27298 21315 27344
rect 21361 27298 21374 27344
rect 21286 27240 21374 27298
rect 21286 27194 21315 27240
rect 21361 27194 21374 27240
rect 21286 27181 21374 27194
rect 21592 28076 21680 28089
rect 21592 28030 21605 28076
rect 21651 28030 21680 28076
rect 21592 27971 21680 28030
rect 21592 27925 21605 27971
rect 21651 27925 21680 27971
rect 21592 27866 21680 27925
rect 21592 27820 21605 27866
rect 21651 27820 21680 27866
rect 21592 27761 21680 27820
rect 21592 27715 21605 27761
rect 21651 27715 21680 27761
rect 21592 27656 21680 27715
rect 21592 27610 21605 27656
rect 21651 27610 21680 27656
rect 21592 27552 21680 27610
rect 21592 27506 21605 27552
rect 21651 27506 21680 27552
rect 21592 27448 21680 27506
rect 21592 27402 21605 27448
rect 21651 27402 21680 27448
rect 21592 27344 21680 27402
rect 21592 27298 21605 27344
rect 21651 27298 21680 27344
rect 21592 27240 21680 27298
rect 21592 27194 21605 27240
rect 21651 27194 21680 27240
rect 21592 27181 21680 27194
rect 21800 28076 21904 28089
rect 21800 28030 21829 28076
rect 21875 28030 21904 28076
rect 21800 27971 21904 28030
rect 21800 27925 21829 27971
rect 21875 27925 21904 27971
rect 21800 27866 21904 27925
rect 21800 27820 21829 27866
rect 21875 27820 21904 27866
rect 21800 27761 21904 27820
rect 21800 27715 21829 27761
rect 21875 27715 21904 27761
rect 21800 27656 21904 27715
rect 21800 27610 21829 27656
rect 21875 27610 21904 27656
rect 21800 27552 21904 27610
rect 21800 27506 21829 27552
rect 21875 27506 21904 27552
rect 21800 27448 21904 27506
rect 21800 27402 21829 27448
rect 21875 27402 21904 27448
rect 21800 27344 21904 27402
rect 21800 27298 21829 27344
rect 21875 27298 21904 27344
rect 21800 27240 21904 27298
rect 21800 27194 21829 27240
rect 21875 27194 21904 27240
rect 21800 27181 21904 27194
rect 22024 28076 22128 28089
rect 22024 28030 22053 28076
rect 22099 28030 22128 28076
rect 22024 27971 22128 28030
rect 22024 27925 22053 27971
rect 22099 27925 22128 27971
rect 22024 27866 22128 27925
rect 22024 27820 22053 27866
rect 22099 27820 22128 27866
rect 22024 27761 22128 27820
rect 22024 27715 22053 27761
rect 22099 27715 22128 27761
rect 22024 27656 22128 27715
rect 22024 27610 22053 27656
rect 22099 27610 22128 27656
rect 22024 27552 22128 27610
rect 22024 27506 22053 27552
rect 22099 27506 22128 27552
rect 22024 27448 22128 27506
rect 22024 27402 22053 27448
rect 22099 27402 22128 27448
rect 22024 27344 22128 27402
rect 22024 27298 22053 27344
rect 22099 27298 22128 27344
rect 22024 27240 22128 27298
rect 22024 27194 22053 27240
rect 22099 27194 22128 27240
rect 22024 27181 22128 27194
rect 22248 28076 22352 28089
rect 22248 28030 22277 28076
rect 22323 28030 22352 28076
rect 22248 27971 22352 28030
rect 22248 27925 22277 27971
rect 22323 27925 22352 27971
rect 22248 27866 22352 27925
rect 22248 27820 22277 27866
rect 22323 27820 22352 27866
rect 22248 27761 22352 27820
rect 22248 27715 22277 27761
rect 22323 27715 22352 27761
rect 22248 27656 22352 27715
rect 22248 27610 22277 27656
rect 22323 27610 22352 27656
rect 22248 27552 22352 27610
rect 22248 27506 22277 27552
rect 22323 27506 22352 27552
rect 22248 27448 22352 27506
rect 22248 27402 22277 27448
rect 22323 27402 22352 27448
rect 22248 27344 22352 27402
rect 22248 27298 22277 27344
rect 22323 27298 22352 27344
rect 22248 27240 22352 27298
rect 22248 27194 22277 27240
rect 22323 27194 22352 27240
rect 22248 27181 22352 27194
rect 22472 28076 22576 28089
rect 22472 28030 22501 28076
rect 22547 28030 22576 28076
rect 22472 27971 22576 28030
rect 22472 27925 22501 27971
rect 22547 27925 22576 27971
rect 22472 27866 22576 27925
rect 22472 27820 22501 27866
rect 22547 27820 22576 27866
rect 22472 27761 22576 27820
rect 22472 27715 22501 27761
rect 22547 27715 22576 27761
rect 22472 27656 22576 27715
rect 22472 27610 22501 27656
rect 22547 27610 22576 27656
rect 22472 27552 22576 27610
rect 22472 27506 22501 27552
rect 22547 27506 22576 27552
rect 22472 27448 22576 27506
rect 22472 27402 22501 27448
rect 22547 27402 22576 27448
rect 22472 27344 22576 27402
rect 22472 27298 22501 27344
rect 22547 27298 22576 27344
rect 22472 27240 22576 27298
rect 22472 27194 22501 27240
rect 22547 27194 22576 27240
rect 22472 27181 22576 27194
rect 22696 28076 22800 28089
rect 22696 28030 22725 28076
rect 22771 28030 22800 28076
rect 22696 27971 22800 28030
rect 22696 27925 22725 27971
rect 22771 27925 22800 27971
rect 22696 27866 22800 27925
rect 22696 27820 22725 27866
rect 22771 27820 22800 27866
rect 22696 27761 22800 27820
rect 22696 27715 22725 27761
rect 22771 27715 22800 27761
rect 22696 27656 22800 27715
rect 22696 27610 22725 27656
rect 22771 27610 22800 27656
rect 22696 27552 22800 27610
rect 22696 27506 22725 27552
rect 22771 27506 22800 27552
rect 22696 27448 22800 27506
rect 22696 27402 22725 27448
rect 22771 27402 22800 27448
rect 22696 27344 22800 27402
rect 22696 27298 22725 27344
rect 22771 27298 22800 27344
rect 22696 27240 22800 27298
rect 22696 27194 22725 27240
rect 22771 27194 22800 27240
rect 22696 27181 22800 27194
rect 22920 28076 23008 28089
rect 22920 28030 22949 28076
rect 22995 28030 23008 28076
rect 22920 27971 23008 28030
rect 22920 27925 22949 27971
rect 22995 27925 23008 27971
rect 22920 27866 23008 27925
rect 22920 27820 22949 27866
rect 22995 27820 23008 27866
rect 23784 28087 23872 28144
rect 23784 28041 23797 28087
rect 23843 28041 23872 28087
rect 23784 27984 23872 28041
rect 23784 27938 23797 27984
rect 23843 27938 23872 27984
rect 23784 27880 23872 27938
rect 23784 27834 23797 27880
rect 23843 27834 23872 27880
rect 23784 27821 23872 27834
rect 23992 28190 24096 28203
rect 23992 28144 24021 28190
rect 24067 28144 24096 28190
rect 23992 28087 24096 28144
rect 23992 28041 24021 28087
rect 24067 28041 24096 28087
rect 23992 27984 24096 28041
rect 23992 27938 24021 27984
rect 24067 27938 24096 27984
rect 23992 27880 24096 27938
rect 23992 27834 24021 27880
rect 24067 27834 24096 27880
rect 23992 27821 24096 27834
rect 24216 28190 24304 28203
rect 24216 28144 24245 28190
rect 24291 28144 24304 28190
rect 24216 28087 24304 28144
rect 24216 28041 24245 28087
rect 24291 28041 24304 28087
rect 25379 28076 25467 28089
rect 24216 27984 24304 28041
rect 24216 27938 24245 27984
rect 24291 27938 24304 27984
rect 24216 27880 24304 27938
rect 24216 27834 24245 27880
rect 24291 27834 24304 27880
rect 24216 27821 24304 27834
rect 22920 27761 23008 27820
rect 22920 27715 22949 27761
rect 22995 27715 23008 27761
rect 22920 27656 23008 27715
rect 22920 27610 22949 27656
rect 22995 27610 23008 27656
rect 22920 27552 23008 27610
rect 22920 27506 22949 27552
rect 22995 27506 23008 27552
rect 25379 27830 25392 28076
rect 25438 27830 25467 28076
rect 25379 27817 25467 27830
rect 25587 28076 25675 28089
rect 25587 27830 25616 28076
rect 25662 27830 25675 28076
rect 25587 27817 25675 27830
rect 22920 27448 23008 27506
rect 22920 27402 22949 27448
rect 22995 27402 23008 27448
rect 22920 27344 23008 27402
rect 22920 27298 22949 27344
rect 22995 27298 23008 27344
rect 22920 27240 23008 27298
rect 22920 27194 22949 27240
rect 22995 27194 23008 27240
rect 22920 27181 23008 27194
rect 13457 26731 13545 26744
rect 13457 26379 13470 26731
rect 13516 26379 13545 26731
rect 13457 26322 13545 26379
rect 13457 26276 13470 26322
rect 13516 26276 13545 26322
rect 13457 26219 13545 26276
rect 13457 26173 13470 26219
rect 13516 26173 13545 26219
rect 13457 26116 13545 26173
rect 13457 26070 13470 26116
rect 13516 26070 13545 26116
rect 13457 26013 13545 26070
rect 13457 25967 13470 26013
rect 13516 25967 13545 26013
rect 13457 25910 13545 25967
rect 13457 25864 13470 25910
rect 13516 25864 13545 25910
rect 13457 25807 13545 25864
rect 13457 25761 13470 25807
rect 13516 25761 13545 25807
rect 13457 25704 13545 25761
rect 13457 25658 13470 25704
rect 13516 25658 13545 25704
rect 13457 25601 13545 25658
rect 13457 25555 13470 25601
rect 13516 25555 13545 25601
rect 13457 25498 13545 25555
rect 13457 25452 13470 25498
rect 13516 25452 13545 25498
rect 13457 25395 13545 25452
rect 13457 25349 13470 25395
rect 13516 25349 13545 25395
rect 13457 25336 13545 25349
rect 13665 26731 13753 26744
rect 13665 26379 13694 26731
rect 13740 26379 13753 26731
rect 15148 26731 15236 26744
rect 13665 26322 13753 26379
rect 13665 26276 13694 26322
rect 13740 26276 13753 26322
rect 13665 26219 13753 26276
rect 13665 26173 13694 26219
rect 13740 26173 13753 26219
rect 13665 26116 13753 26173
rect 13665 26070 13694 26116
rect 13740 26070 13753 26116
rect 13665 26013 13753 26070
rect 13665 25967 13694 26013
rect 13740 25967 13753 26013
rect 13665 25910 13753 25967
rect 13665 25864 13694 25910
rect 13740 25864 13753 25910
rect 13665 25807 13753 25864
rect 13665 25761 13694 25807
rect 13740 25761 13753 25807
rect 13665 25704 13753 25761
rect 13665 25658 13694 25704
rect 13740 25658 13753 25704
rect 13665 25601 13753 25658
rect 13665 25555 13694 25601
rect 13740 25555 13753 25601
rect 13665 25498 13753 25555
rect 13665 25452 13694 25498
rect 13740 25452 13753 25498
rect 13665 25395 13753 25452
rect 13971 26446 14059 26459
rect 13971 26400 13984 26446
rect 14030 26400 14059 26446
rect 13971 26338 14059 26400
rect 13971 26292 13984 26338
rect 14030 26292 14059 26338
rect 13971 26230 14059 26292
rect 13971 26184 13984 26230
rect 14030 26184 14059 26230
rect 13971 26122 14059 26184
rect 13971 26076 13984 26122
rect 14030 26076 14059 26122
rect 13971 26014 14059 26076
rect 13971 25968 13984 26014
rect 14030 25968 14059 26014
rect 13971 25906 14059 25968
rect 13971 25860 13984 25906
rect 14030 25860 14059 25906
rect 13971 25798 14059 25860
rect 13971 25752 13984 25798
rect 14030 25752 14059 25798
rect 13971 25690 14059 25752
rect 13971 25644 13984 25690
rect 14030 25644 14059 25690
rect 13971 25582 14059 25644
rect 13971 25536 13984 25582
rect 14030 25536 14059 25582
rect 13971 25474 14059 25536
rect 13971 25428 13984 25474
rect 14030 25428 14059 25474
rect 13971 25415 14059 25428
rect 14179 26446 14267 26459
rect 14179 26400 14208 26446
rect 14254 26400 14267 26446
rect 14179 26338 14267 26400
rect 14179 26292 14208 26338
rect 14254 26292 14267 26338
rect 14179 26230 14267 26292
rect 14179 26184 14208 26230
rect 14254 26184 14267 26230
rect 14179 26122 14267 26184
rect 14179 26076 14208 26122
rect 14254 26076 14267 26122
rect 14179 26014 14267 26076
rect 14179 25968 14208 26014
rect 14254 25968 14267 26014
rect 14179 25906 14267 25968
rect 14179 25860 14208 25906
rect 14254 25860 14267 25906
rect 14179 25798 14267 25860
rect 14179 25752 14208 25798
rect 14254 25752 14267 25798
rect 14179 25690 14267 25752
rect 14179 25644 14208 25690
rect 14254 25644 14267 25690
rect 14179 25582 14267 25644
rect 14179 25536 14208 25582
rect 14254 25536 14267 25582
rect 14179 25474 14267 25536
rect 14179 25428 14208 25474
rect 14254 25428 14267 25474
rect 15148 26379 15161 26731
rect 15207 26379 15236 26731
rect 15148 26322 15236 26379
rect 15148 26276 15161 26322
rect 15207 26276 15236 26322
rect 15148 26219 15236 26276
rect 15148 26173 15161 26219
rect 15207 26173 15236 26219
rect 15148 26116 15236 26173
rect 15148 26070 15161 26116
rect 15207 26070 15236 26116
rect 15148 26013 15236 26070
rect 15148 25967 15161 26013
rect 15207 25967 15236 26013
rect 15148 25910 15236 25967
rect 15148 25864 15161 25910
rect 15207 25864 15236 25910
rect 15148 25807 15236 25864
rect 15148 25761 15161 25807
rect 15207 25761 15236 25807
rect 15148 25704 15236 25761
rect 15148 25658 15161 25704
rect 15207 25658 15236 25704
rect 15148 25601 15236 25658
rect 15148 25555 15161 25601
rect 15207 25555 15236 25601
rect 15148 25498 15236 25555
rect 14179 25415 14267 25428
rect 15148 25452 15161 25498
rect 15207 25452 15236 25498
rect 13665 25349 13694 25395
rect 13740 25349 13753 25395
rect 13665 25336 13753 25349
rect 15148 25395 15236 25452
rect 15148 25349 15161 25395
rect 15207 25349 15236 25395
rect 15148 25336 15236 25349
rect 15356 26731 15444 26744
rect 15356 26379 15385 26731
rect 15431 26379 15444 26731
rect 15356 26322 15444 26379
rect 15356 26276 15385 26322
rect 15431 26276 15444 26322
rect 15356 26219 15444 26276
rect 15356 26173 15385 26219
rect 15431 26173 15444 26219
rect 15356 26116 15444 26173
rect 15356 26070 15385 26116
rect 15431 26070 15444 26116
rect 15356 26013 15444 26070
rect 15356 25967 15385 26013
rect 15431 25967 15444 26013
rect 15356 25910 15444 25967
rect 15356 25864 15385 25910
rect 15431 25864 15444 25910
rect 15356 25807 15444 25864
rect 15356 25761 15385 25807
rect 15431 25761 15444 25807
rect 15356 25704 15444 25761
rect 15356 25658 15385 25704
rect 15431 25658 15444 25704
rect 15356 25601 15444 25658
rect 15356 25555 15385 25601
rect 15431 25555 15444 25601
rect 15356 25498 15444 25555
rect 15356 25452 15385 25498
rect 15431 25452 15444 25498
rect 15356 25395 15444 25452
rect 15662 26446 15750 26459
rect 15662 26400 15675 26446
rect 15721 26400 15750 26446
rect 15662 26338 15750 26400
rect 15662 26292 15675 26338
rect 15721 26292 15750 26338
rect 15662 26230 15750 26292
rect 15662 26184 15675 26230
rect 15721 26184 15750 26230
rect 15662 26122 15750 26184
rect 15662 26076 15675 26122
rect 15721 26076 15750 26122
rect 15662 26014 15750 26076
rect 15662 25968 15675 26014
rect 15721 25968 15750 26014
rect 15662 25906 15750 25968
rect 15662 25860 15675 25906
rect 15721 25860 15750 25906
rect 15662 25798 15750 25860
rect 15662 25752 15675 25798
rect 15721 25752 15750 25798
rect 15662 25690 15750 25752
rect 15662 25644 15675 25690
rect 15721 25644 15750 25690
rect 15662 25582 15750 25644
rect 15662 25536 15675 25582
rect 15721 25536 15750 25582
rect 15662 25474 15750 25536
rect 15662 25428 15675 25474
rect 15721 25428 15750 25474
rect 15662 25415 15750 25428
rect 15870 26446 15958 26459
rect 15870 26400 15899 26446
rect 15945 26400 15958 26446
rect 15870 26338 15958 26400
rect 15870 26292 15899 26338
rect 15945 26292 15958 26338
rect 15870 26230 15958 26292
rect 15870 26184 15899 26230
rect 15945 26184 15958 26230
rect 15870 26122 15958 26184
rect 15870 26076 15899 26122
rect 15945 26076 15958 26122
rect 15870 26014 15958 26076
rect 15870 25968 15899 26014
rect 15945 25968 15958 26014
rect 15870 25906 15958 25968
rect 15870 25860 15899 25906
rect 15945 25860 15958 25906
rect 15870 25798 15958 25860
rect 15870 25752 15899 25798
rect 15945 25752 15958 25798
rect 15870 25690 15958 25752
rect 15870 25644 15899 25690
rect 15945 25644 15958 25690
rect 15870 25582 15958 25644
rect 15870 25536 15899 25582
rect 15945 25536 15958 25582
rect 15870 25474 15958 25536
rect 15870 25428 15899 25474
rect 15945 25428 15958 25474
rect 15870 25415 15958 25428
rect 15356 25349 15385 25395
rect 15431 25349 15444 25395
rect 15356 25336 15444 25349
rect 23943 26730 24031 26743
rect 23943 26684 23956 26730
rect 24002 26684 24031 26730
rect 23943 26627 24031 26684
rect 23943 26581 23956 26627
rect 24002 26581 24031 26627
rect 23943 26524 24031 26581
rect 23943 26478 23956 26524
rect 24002 26478 24031 26524
rect 23943 26421 24031 26478
rect 23943 26375 23956 26421
rect 24002 26375 24031 26421
rect 23943 26318 24031 26375
rect 23943 26272 23956 26318
rect 24002 26272 24031 26318
rect 23943 26214 24031 26272
rect 23943 26168 23956 26214
rect 24002 26168 24031 26214
rect 23943 26110 24031 26168
rect 23943 26064 23956 26110
rect 24002 26064 24031 26110
rect 23943 26006 24031 26064
rect 23943 25960 23956 26006
rect 24002 25960 24031 26006
rect 23943 25902 24031 25960
rect 23943 25856 23956 25902
rect 24002 25856 24031 25902
rect 23943 25798 24031 25856
rect 23943 25752 23956 25798
rect 24002 25752 24031 25798
rect 23943 25694 24031 25752
rect 23943 25648 23956 25694
rect 24002 25648 24031 25694
rect 23943 25590 24031 25648
rect 23943 25544 23956 25590
rect 24002 25544 24031 25590
rect 23943 25486 24031 25544
rect 23943 25440 23956 25486
rect 24002 25440 24031 25486
rect 23943 25427 24031 25440
rect 24151 26730 24239 26743
rect 24151 26684 24180 26730
rect 24226 26684 24239 26730
rect 24151 26627 24239 26684
rect 24151 26581 24180 26627
rect 24226 26581 24239 26627
rect 24151 26524 24239 26581
rect 24151 26478 24180 26524
rect 24226 26478 24239 26524
rect 24151 26421 24239 26478
rect 24151 26375 24180 26421
rect 24226 26375 24239 26421
rect 24151 26318 24239 26375
rect 24151 26272 24180 26318
rect 24226 26272 24239 26318
rect 24151 26214 24239 26272
rect 24151 26168 24180 26214
rect 24226 26168 24239 26214
rect 24151 26110 24239 26168
rect 24151 26064 24180 26110
rect 24226 26064 24239 26110
rect 24151 26006 24239 26064
rect 24151 25960 24180 26006
rect 24226 25960 24239 26006
rect 24151 25902 24239 25960
rect 24151 25856 24180 25902
rect 24226 25856 24239 25902
rect 24151 25798 24239 25856
rect 24151 25752 24180 25798
rect 24226 25752 24239 25798
rect 24151 25694 24239 25752
rect 24151 25648 24180 25694
rect 24226 25648 24239 25694
rect 24151 25590 24239 25648
rect 24151 25544 24180 25590
rect 24226 25544 24239 25590
rect 24151 25486 24239 25544
rect 24151 25440 24180 25486
rect 24226 25440 24239 25486
rect 24151 25427 24239 25440
rect 24457 26730 24545 26743
rect 24457 26684 24470 26730
rect 24516 26684 24545 26730
rect 24457 26627 24545 26684
rect 24457 26581 24470 26627
rect 24516 26581 24545 26627
rect 24457 26524 24545 26581
rect 24457 26478 24470 26524
rect 24516 26478 24545 26524
rect 24457 26421 24545 26478
rect 24457 26375 24470 26421
rect 24516 26375 24545 26421
rect 24457 26318 24545 26375
rect 24457 26272 24470 26318
rect 24516 26272 24545 26318
rect 24457 26214 24545 26272
rect 24457 26168 24470 26214
rect 24516 26168 24545 26214
rect 24457 26110 24545 26168
rect 24457 26064 24470 26110
rect 24516 26064 24545 26110
rect 24457 26006 24545 26064
rect 24457 25960 24470 26006
rect 24516 25960 24545 26006
rect 24457 25902 24545 25960
rect 24457 25856 24470 25902
rect 24516 25856 24545 25902
rect 24457 25798 24545 25856
rect 24457 25752 24470 25798
rect 24516 25752 24545 25798
rect 24457 25694 24545 25752
rect 24457 25648 24470 25694
rect 24516 25648 24545 25694
rect 24457 25590 24545 25648
rect 24457 25544 24470 25590
rect 24516 25544 24545 25590
rect 24457 25486 24545 25544
rect 24457 25440 24470 25486
rect 24516 25440 24545 25486
rect 24457 25427 24545 25440
rect 24665 26730 24753 26743
rect 24665 26684 24694 26730
rect 24740 26684 24753 26730
rect 25633 26730 25721 26743
rect 24665 26627 24753 26684
rect 24665 26581 24694 26627
rect 24740 26581 24753 26627
rect 24665 26524 24753 26581
rect 24665 26478 24694 26524
rect 24740 26478 24753 26524
rect 24665 26421 24753 26478
rect 24665 26375 24694 26421
rect 24740 26375 24753 26421
rect 24665 26318 24753 26375
rect 24665 26272 24694 26318
rect 24740 26272 24753 26318
rect 24665 26214 24753 26272
rect 24665 26168 24694 26214
rect 24740 26168 24753 26214
rect 24665 26110 24753 26168
rect 24665 26064 24694 26110
rect 24740 26064 24753 26110
rect 24665 26006 24753 26064
rect 24665 25960 24694 26006
rect 24740 25960 24753 26006
rect 24665 25902 24753 25960
rect 24665 25856 24694 25902
rect 24740 25856 24753 25902
rect 24665 25798 24753 25856
rect 24665 25752 24694 25798
rect 24740 25752 24753 25798
rect 24665 25694 24753 25752
rect 24665 25648 24694 25694
rect 24740 25648 24753 25694
rect 24665 25590 24753 25648
rect 24665 25544 24694 25590
rect 24740 25544 24753 25590
rect 25633 26684 25646 26730
rect 25692 26684 25721 26730
rect 25633 26627 25721 26684
rect 25633 26581 25646 26627
rect 25692 26581 25721 26627
rect 25633 26524 25721 26581
rect 25633 26478 25646 26524
rect 25692 26478 25721 26524
rect 25633 26421 25721 26478
rect 25633 26375 25646 26421
rect 25692 26375 25721 26421
rect 25633 26318 25721 26375
rect 25633 26272 25646 26318
rect 25692 26272 25721 26318
rect 25633 26214 25721 26272
rect 25633 26168 25646 26214
rect 25692 26168 25721 26214
rect 25633 26110 25721 26168
rect 25633 26064 25646 26110
rect 25692 26064 25721 26110
rect 25633 26006 25721 26064
rect 25633 25960 25646 26006
rect 25692 25960 25721 26006
rect 25633 25902 25721 25960
rect 25633 25856 25646 25902
rect 25692 25856 25721 25902
rect 25633 25798 25721 25856
rect 25633 25752 25646 25798
rect 25692 25752 25721 25798
rect 25633 25694 25721 25752
rect 25633 25648 25646 25694
rect 25692 25648 25721 25694
rect 25633 25590 25721 25648
rect 24665 25486 24753 25544
rect 24665 25440 24694 25486
rect 24740 25440 24753 25486
rect 24665 25427 24753 25440
rect 25633 25544 25646 25590
rect 25692 25544 25721 25590
rect 25633 25486 25721 25544
rect 25633 25440 25646 25486
rect 25692 25440 25721 25486
rect 25633 25427 25721 25440
rect 25841 26730 25929 26743
rect 25841 26684 25870 26730
rect 25916 26684 25929 26730
rect 25841 26627 25929 26684
rect 25841 26581 25870 26627
rect 25916 26581 25929 26627
rect 25841 26524 25929 26581
rect 25841 26478 25870 26524
rect 25916 26478 25929 26524
rect 25841 26421 25929 26478
rect 25841 26375 25870 26421
rect 25916 26375 25929 26421
rect 25841 26318 25929 26375
rect 25841 26272 25870 26318
rect 25916 26272 25929 26318
rect 25841 26214 25929 26272
rect 25841 26168 25870 26214
rect 25916 26168 25929 26214
rect 25841 26110 25929 26168
rect 25841 26064 25870 26110
rect 25916 26064 25929 26110
rect 25841 26006 25929 26064
rect 25841 25960 25870 26006
rect 25916 25960 25929 26006
rect 25841 25902 25929 25960
rect 25841 25856 25870 25902
rect 25916 25856 25929 25902
rect 25841 25798 25929 25856
rect 25841 25752 25870 25798
rect 25916 25752 25929 25798
rect 25841 25694 25929 25752
rect 25841 25648 25870 25694
rect 25916 25648 25929 25694
rect 25841 25590 25929 25648
rect 25841 25544 25870 25590
rect 25916 25544 25929 25590
rect 25841 25486 25929 25544
rect 25841 25440 25870 25486
rect 25916 25440 25929 25486
rect 25841 25427 25929 25440
rect 26147 26730 26235 26743
rect 26147 26684 26160 26730
rect 26206 26684 26235 26730
rect 26147 26627 26235 26684
rect 26147 26581 26160 26627
rect 26206 26581 26235 26627
rect 26147 26524 26235 26581
rect 26147 26478 26160 26524
rect 26206 26478 26235 26524
rect 26147 26421 26235 26478
rect 26147 26375 26160 26421
rect 26206 26375 26235 26421
rect 26147 26318 26235 26375
rect 26147 26272 26160 26318
rect 26206 26272 26235 26318
rect 26147 26214 26235 26272
rect 26147 26168 26160 26214
rect 26206 26168 26235 26214
rect 26147 26110 26235 26168
rect 26147 26064 26160 26110
rect 26206 26064 26235 26110
rect 26147 26006 26235 26064
rect 26147 25960 26160 26006
rect 26206 25960 26235 26006
rect 26147 25902 26235 25960
rect 26147 25856 26160 25902
rect 26206 25856 26235 25902
rect 26147 25798 26235 25856
rect 26147 25752 26160 25798
rect 26206 25752 26235 25798
rect 26147 25694 26235 25752
rect 26147 25648 26160 25694
rect 26206 25648 26235 25694
rect 26147 25590 26235 25648
rect 26147 25544 26160 25590
rect 26206 25544 26235 25590
rect 26147 25486 26235 25544
rect 26147 25440 26160 25486
rect 26206 25440 26235 25486
rect 26147 25427 26235 25440
rect 26355 26730 26443 26743
rect 26355 26684 26384 26730
rect 26430 26684 26443 26730
rect 27324 26730 27412 26743
rect 26355 26627 26443 26684
rect 26355 26581 26384 26627
rect 26430 26581 26443 26627
rect 26355 26524 26443 26581
rect 26355 26478 26384 26524
rect 26430 26478 26443 26524
rect 26355 26421 26443 26478
rect 26355 26375 26384 26421
rect 26430 26375 26443 26421
rect 26355 26318 26443 26375
rect 26355 26272 26384 26318
rect 26430 26272 26443 26318
rect 26355 26214 26443 26272
rect 26355 26168 26384 26214
rect 26430 26168 26443 26214
rect 26355 26110 26443 26168
rect 26355 26064 26384 26110
rect 26430 26064 26443 26110
rect 26355 26006 26443 26064
rect 26355 25960 26384 26006
rect 26430 25960 26443 26006
rect 26355 25902 26443 25960
rect 26355 25856 26384 25902
rect 26430 25856 26443 25902
rect 26355 25798 26443 25856
rect 26355 25752 26384 25798
rect 26430 25752 26443 25798
rect 26355 25694 26443 25752
rect 26355 25648 26384 25694
rect 26430 25648 26443 25694
rect 26355 25590 26443 25648
rect 26355 25544 26384 25590
rect 26430 25544 26443 25590
rect 27324 26684 27337 26730
rect 27383 26684 27412 26730
rect 27324 26627 27412 26684
rect 27324 26581 27337 26627
rect 27383 26581 27412 26627
rect 27324 26524 27412 26581
rect 27324 26478 27337 26524
rect 27383 26478 27412 26524
rect 27324 26421 27412 26478
rect 27324 26375 27337 26421
rect 27383 26375 27412 26421
rect 27324 26318 27412 26375
rect 27324 26272 27337 26318
rect 27383 26272 27412 26318
rect 27324 26214 27412 26272
rect 27324 26168 27337 26214
rect 27383 26168 27412 26214
rect 27324 26110 27412 26168
rect 27324 26064 27337 26110
rect 27383 26064 27412 26110
rect 27324 26006 27412 26064
rect 27324 25960 27337 26006
rect 27383 25960 27412 26006
rect 27324 25902 27412 25960
rect 27324 25856 27337 25902
rect 27383 25856 27412 25902
rect 27324 25798 27412 25856
rect 27324 25752 27337 25798
rect 27383 25752 27412 25798
rect 27324 25694 27412 25752
rect 27324 25648 27337 25694
rect 27383 25648 27412 25694
rect 27324 25590 27412 25648
rect 26355 25486 26443 25544
rect 26355 25440 26384 25486
rect 26430 25440 26443 25486
rect 26355 25427 26443 25440
rect 27324 25544 27337 25590
rect 27383 25544 27412 25590
rect 27324 25486 27412 25544
rect 27324 25440 27337 25486
rect 27383 25440 27412 25486
rect 27324 25427 27412 25440
rect 27532 26730 27620 26743
rect 27532 26684 27561 26730
rect 27607 26684 27620 26730
rect 27532 26627 27620 26684
rect 27532 26581 27561 26627
rect 27607 26581 27620 26627
rect 27532 26524 27620 26581
rect 27532 26478 27561 26524
rect 27607 26478 27620 26524
rect 27532 26421 27620 26478
rect 27532 26375 27561 26421
rect 27607 26375 27620 26421
rect 27532 26318 27620 26375
rect 27532 26272 27561 26318
rect 27607 26272 27620 26318
rect 27532 26214 27620 26272
rect 27532 26168 27561 26214
rect 27607 26168 27620 26214
rect 27532 26110 27620 26168
rect 27532 26064 27561 26110
rect 27607 26064 27620 26110
rect 27532 26006 27620 26064
rect 27532 25960 27561 26006
rect 27607 25960 27620 26006
rect 27532 25902 27620 25960
rect 27532 25856 27561 25902
rect 27607 25856 27620 25902
rect 27532 25798 27620 25856
rect 27532 25752 27561 25798
rect 27607 25752 27620 25798
rect 27532 25694 27620 25752
rect 27532 25648 27561 25694
rect 27607 25648 27620 25694
rect 27532 25590 27620 25648
rect 27532 25544 27561 25590
rect 27607 25544 27620 25590
rect 27532 25486 27620 25544
rect 27532 25440 27561 25486
rect 27607 25440 27620 25486
rect 27532 25427 27620 25440
rect 27838 26730 27926 26743
rect 27838 26684 27851 26730
rect 27897 26684 27926 26730
rect 27838 26627 27926 26684
rect 27838 26581 27851 26627
rect 27897 26581 27926 26627
rect 27838 26524 27926 26581
rect 27838 26478 27851 26524
rect 27897 26478 27926 26524
rect 27838 26421 27926 26478
rect 27838 26375 27851 26421
rect 27897 26375 27926 26421
rect 27838 26318 27926 26375
rect 27838 26272 27851 26318
rect 27897 26272 27926 26318
rect 27838 26214 27926 26272
rect 27838 26168 27851 26214
rect 27897 26168 27926 26214
rect 27838 26110 27926 26168
rect 27838 26064 27851 26110
rect 27897 26064 27926 26110
rect 27838 26006 27926 26064
rect 27838 25960 27851 26006
rect 27897 25960 27926 26006
rect 27838 25902 27926 25960
rect 27838 25856 27851 25902
rect 27897 25856 27926 25902
rect 27838 25798 27926 25856
rect 27838 25752 27851 25798
rect 27897 25752 27926 25798
rect 27838 25694 27926 25752
rect 27838 25648 27851 25694
rect 27897 25648 27926 25694
rect 27838 25590 27926 25648
rect 27838 25544 27851 25590
rect 27897 25544 27926 25590
rect 27838 25486 27926 25544
rect 27838 25440 27851 25486
rect 27897 25440 27926 25486
rect 27838 25427 27926 25440
rect 28046 26730 28134 26743
rect 28046 26684 28075 26730
rect 28121 26684 28134 26730
rect 28046 26627 28134 26684
rect 28046 26581 28075 26627
rect 28121 26581 28134 26627
rect 28046 26524 28134 26581
rect 28046 26478 28075 26524
rect 28121 26478 28134 26524
rect 28046 26421 28134 26478
rect 28046 26375 28075 26421
rect 28121 26375 28134 26421
rect 28046 26318 28134 26375
rect 28046 26272 28075 26318
rect 28121 26272 28134 26318
rect 28046 26214 28134 26272
rect 28046 26168 28075 26214
rect 28121 26168 28134 26214
rect 28046 26110 28134 26168
rect 28046 26064 28075 26110
rect 28121 26064 28134 26110
rect 28046 26006 28134 26064
rect 28046 25960 28075 26006
rect 28121 25960 28134 26006
rect 28046 25902 28134 25960
rect 28046 25856 28075 25902
rect 28121 25856 28134 25902
rect 28046 25798 28134 25856
rect 28046 25752 28075 25798
rect 28121 25752 28134 25798
rect 28046 25694 28134 25752
rect 28046 25648 28075 25694
rect 28121 25648 28134 25694
rect 28046 25590 28134 25648
rect 28046 25544 28075 25590
rect 28121 25544 28134 25590
rect 28046 25486 28134 25544
rect 28046 25440 28075 25486
rect 28121 25440 28134 25486
rect 28046 25427 28134 25440
rect 1774 20506 1892 20551
rect 1774 20460 1817 20506
rect 1863 20460 1892 20506
rect 1774 20338 1892 20460
rect 1774 20292 1817 20338
rect 1863 20292 1892 20338
rect 1774 20171 1892 20292
rect 1774 20125 1817 20171
rect 1863 20125 1892 20171
rect 1774 20003 1892 20125
rect 1774 19957 1817 20003
rect 1863 19957 1892 20003
rect 1774 19835 1892 19957
rect 1774 19789 1817 19835
rect 1863 19789 1892 19835
rect 1774 19667 1892 19789
rect 1774 19621 1817 19667
rect 1863 19621 1892 19667
rect 1774 19499 1892 19621
rect 1774 19453 1817 19499
rect 1863 19453 1892 19499
rect 1774 19332 1892 19453
rect 1774 19286 1817 19332
rect 1863 19286 1892 19332
rect 1774 19164 1892 19286
rect 1774 19118 1817 19164
rect 1863 19118 1892 19164
rect 1774 18996 1892 19118
rect 1774 18950 1817 18996
rect 1863 18950 1892 18996
rect 1774 18828 1892 18950
rect 1774 18782 1817 18828
rect 1863 18782 1892 18828
rect 1774 18658 1892 18782
rect 1774 18612 1817 18658
rect 1863 18612 1892 18658
rect 1774 18488 1892 18612
rect 1774 18442 1817 18488
rect 1863 18442 1892 18488
rect 1774 18318 1892 18442
rect 1774 18272 1817 18318
rect 1863 18272 1892 18318
rect 1774 18101 1892 18272
rect 2012 18101 2116 20551
rect 2236 20506 2355 20551
rect 2236 20460 2266 20506
rect 2312 20460 2355 20506
rect 2236 20338 2355 20460
rect 2236 20292 2266 20338
rect 2312 20292 2355 20338
rect 2236 20171 2355 20292
rect 2236 20125 2266 20171
rect 2312 20125 2355 20171
rect 2236 20003 2355 20125
rect 2236 19957 2266 20003
rect 2312 19957 2355 20003
rect 2236 19835 2355 19957
rect 2236 19789 2266 19835
rect 2312 19789 2355 19835
rect 2236 19667 2355 19789
rect 2236 19621 2266 19667
rect 2312 19621 2355 19667
rect 2236 19499 2355 19621
rect 2236 19453 2266 19499
rect 2312 19453 2355 19499
rect 2236 19332 2355 19453
rect 2236 19286 2266 19332
rect 2312 19286 2355 19332
rect 2236 19164 2355 19286
rect 2236 19118 2266 19164
rect 2312 19118 2355 19164
rect 2236 18996 2355 19118
rect 2236 18950 2266 18996
rect 2312 18950 2355 18996
rect 2236 18828 2355 18950
rect 2236 18782 2266 18828
rect 2312 18782 2355 18828
rect 2236 18658 2355 18782
rect 2236 18612 2266 18658
rect 2312 18612 2355 18658
rect 2236 18488 2355 18612
rect 2236 18442 2266 18488
rect 2312 18442 2355 18488
rect 2236 18318 2355 18442
rect 2236 18272 2266 18318
rect 2312 18272 2355 18318
rect 2236 18101 2355 18272
rect 2801 20506 2920 20551
rect 2801 20460 2844 20506
rect 2890 20460 2920 20506
rect 2801 20338 2920 20460
rect 2801 20292 2844 20338
rect 2890 20292 2920 20338
rect 2801 20171 2920 20292
rect 2801 20125 2844 20171
rect 2890 20125 2920 20171
rect 2801 20003 2920 20125
rect 2801 19957 2844 20003
rect 2890 19957 2920 20003
rect 2801 19835 2920 19957
rect 2801 19789 2844 19835
rect 2890 19789 2920 19835
rect 2801 19667 2920 19789
rect 2801 19621 2844 19667
rect 2890 19621 2920 19667
rect 2801 19499 2920 19621
rect 2801 19453 2844 19499
rect 2890 19453 2920 19499
rect 2801 19332 2920 19453
rect 2801 19286 2844 19332
rect 2890 19286 2920 19332
rect 2801 19164 2920 19286
rect 2801 19118 2844 19164
rect 2890 19118 2920 19164
rect 2801 18996 2920 19118
rect 2801 18950 2844 18996
rect 2890 18950 2920 18996
rect 2801 18828 2920 18950
rect 2801 18782 2844 18828
rect 2890 18782 2920 18828
rect 2801 18658 2920 18782
rect 2801 18612 2844 18658
rect 2890 18612 2920 18658
rect 2801 18488 2920 18612
rect 2801 18442 2844 18488
rect 2890 18442 2920 18488
rect 2801 18318 2920 18442
rect 2801 18272 2844 18318
rect 2890 18272 2920 18318
rect 2801 18101 2920 18272
rect 3040 18101 3144 20551
rect 3264 20506 3382 20551
rect 3264 20460 3293 20506
rect 3339 20460 3382 20506
rect 3264 20338 3382 20460
rect 3264 20292 3293 20338
rect 3339 20292 3382 20338
rect 3264 20171 3382 20292
rect 3264 20125 3293 20171
rect 3339 20125 3382 20171
rect 3264 20003 3382 20125
rect 3264 19957 3293 20003
rect 3339 19957 3382 20003
rect 3264 19835 3382 19957
rect 3264 19789 3293 19835
rect 3339 19789 3382 19835
rect 3264 19667 3382 19789
rect 3264 19621 3293 19667
rect 3339 19621 3382 19667
rect 3264 19499 3382 19621
rect 3264 19453 3293 19499
rect 3339 19453 3382 19499
rect 3264 19332 3382 19453
rect 3264 19286 3293 19332
rect 3339 19286 3382 19332
rect 3264 19164 3382 19286
rect 3264 19118 3293 19164
rect 3339 19118 3382 19164
rect 3264 18996 3382 19118
rect 3264 18950 3293 18996
rect 3339 18950 3382 18996
rect 3264 18828 3382 18950
rect 3264 18782 3293 18828
rect 3339 18782 3382 18828
rect 3264 18658 3382 18782
rect 3264 18612 3293 18658
rect 3339 18612 3382 18658
rect 3264 18488 3382 18612
rect 3264 18442 3293 18488
rect 3339 18442 3382 18488
rect 3264 18318 3382 18442
rect 3264 18272 3293 18318
rect 3339 18272 3382 18318
rect 3264 18101 3382 18272
rect 3566 20506 3684 20551
rect 3566 20460 3609 20506
rect 3655 20460 3684 20506
rect 3566 20338 3684 20460
rect 3566 20292 3609 20338
rect 3655 20292 3684 20338
rect 3566 20171 3684 20292
rect 3566 20125 3609 20171
rect 3655 20125 3684 20171
rect 3566 20003 3684 20125
rect 3566 19957 3609 20003
rect 3655 19957 3684 20003
rect 3566 19835 3684 19957
rect 3566 19789 3609 19835
rect 3655 19789 3684 19835
rect 3566 19667 3684 19789
rect 3566 19621 3609 19667
rect 3655 19621 3684 19667
rect 3566 19499 3684 19621
rect 3566 19453 3609 19499
rect 3655 19453 3684 19499
rect 3566 19332 3684 19453
rect 3566 19286 3609 19332
rect 3655 19286 3684 19332
rect 3566 19164 3684 19286
rect 3566 19118 3609 19164
rect 3655 19118 3684 19164
rect 3566 18996 3684 19118
rect 3566 18950 3609 18996
rect 3655 18950 3684 18996
rect 3566 18828 3684 18950
rect 3566 18782 3609 18828
rect 3655 18782 3684 18828
rect 3566 18658 3684 18782
rect 3566 18612 3609 18658
rect 3655 18612 3684 18658
rect 3566 18488 3684 18612
rect 3566 18442 3609 18488
rect 3655 18442 3684 18488
rect 3566 18318 3684 18442
rect 3566 18272 3609 18318
rect 3655 18272 3684 18318
rect 3566 18101 3684 18272
rect 3804 18101 3908 20551
rect 4028 20506 4147 20551
rect 4028 20460 4058 20506
rect 4104 20460 4147 20506
rect 4028 20338 4147 20460
rect 4028 20292 4058 20338
rect 4104 20292 4147 20338
rect 4028 20171 4147 20292
rect 4028 20125 4058 20171
rect 4104 20125 4147 20171
rect 4028 20003 4147 20125
rect 4028 19957 4058 20003
rect 4104 19957 4147 20003
rect 4028 19835 4147 19957
rect 4028 19789 4058 19835
rect 4104 19789 4147 19835
rect 4028 19667 4147 19789
rect 4028 19621 4058 19667
rect 4104 19621 4147 19667
rect 4028 19499 4147 19621
rect 4028 19453 4058 19499
rect 4104 19453 4147 19499
rect 4028 19332 4147 19453
rect 4028 19286 4058 19332
rect 4104 19286 4147 19332
rect 4028 19164 4147 19286
rect 4028 19118 4058 19164
rect 4104 19118 4147 19164
rect 4028 18996 4147 19118
rect 4028 18950 4058 18996
rect 4104 18950 4147 18996
rect 4028 18828 4147 18950
rect 4028 18782 4058 18828
rect 4104 18782 4147 18828
rect 4028 18658 4147 18782
rect 4028 18612 4058 18658
rect 4104 18612 4147 18658
rect 4028 18488 4147 18612
rect 4028 18442 4058 18488
rect 4104 18442 4147 18488
rect 4028 18318 4147 18442
rect 4028 18272 4058 18318
rect 4104 18272 4147 18318
rect 4028 18101 4147 18272
rect 4593 20506 4712 20551
rect 4593 20460 4636 20506
rect 4682 20460 4712 20506
rect 4593 20338 4712 20460
rect 4593 20292 4636 20338
rect 4682 20292 4712 20338
rect 4593 20171 4712 20292
rect 4593 20125 4636 20171
rect 4682 20125 4712 20171
rect 4593 20003 4712 20125
rect 4593 19957 4636 20003
rect 4682 19957 4712 20003
rect 4593 19835 4712 19957
rect 4593 19789 4636 19835
rect 4682 19789 4712 19835
rect 4593 19667 4712 19789
rect 4593 19621 4636 19667
rect 4682 19621 4712 19667
rect 4593 19499 4712 19621
rect 4593 19453 4636 19499
rect 4682 19453 4712 19499
rect 4593 19332 4712 19453
rect 4593 19286 4636 19332
rect 4682 19286 4712 19332
rect 4593 19164 4712 19286
rect 4593 19118 4636 19164
rect 4682 19118 4712 19164
rect 4593 18996 4712 19118
rect 4593 18950 4636 18996
rect 4682 18950 4712 18996
rect 4593 18828 4712 18950
rect 4593 18782 4636 18828
rect 4682 18782 4712 18828
rect 4593 18658 4712 18782
rect 4593 18612 4636 18658
rect 4682 18612 4712 18658
rect 4593 18488 4712 18612
rect 4593 18442 4636 18488
rect 4682 18442 4712 18488
rect 4593 18318 4712 18442
rect 4593 18272 4636 18318
rect 4682 18272 4712 18318
rect 4593 18101 4712 18272
rect 4832 18101 4936 20551
rect 5056 20506 5174 20551
rect 5056 20460 5085 20506
rect 5131 20460 5174 20506
rect 5056 20338 5174 20460
rect 5056 20292 5085 20338
rect 5131 20292 5174 20338
rect 5056 20171 5174 20292
rect 5056 20125 5085 20171
rect 5131 20125 5174 20171
rect 5056 20003 5174 20125
rect 5056 19957 5085 20003
rect 5131 19957 5174 20003
rect 5056 19835 5174 19957
rect 5056 19789 5085 19835
rect 5131 19789 5174 19835
rect 5056 19667 5174 19789
rect 5056 19621 5085 19667
rect 5131 19621 5174 19667
rect 5056 19499 5174 19621
rect 5056 19453 5085 19499
rect 5131 19453 5174 19499
rect 5056 19332 5174 19453
rect 5056 19286 5085 19332
rect 5131 19286 5174 19332
rect 5056 19164 5174 19286
rect 5056 19118 5085 19164
rect 5131 19118 5174 19164
rect 5056 18996 5174 19118
rect 5056 18950 5085 18996
rect 5131 18950 5174 18996
rect 5056 18828 5174 18950
rect 5056 18782 5085 18828
rect 5131 18782 5174 18828
rect 5056 18658 5174 18782
rect 5056 18612 5085 18658
rect 5131 18612 5174 18658
rect 5056 18488 5174 18612
rect 5056 18442 5085 18488
rect 5131 18442 5174 18488
rect 5056 18318 5174 18442
rect 5056 18272 5085 18318
rect 5131 18272 5174 18318
rect 5056 18101 5174 18272
rect 9153 20506 9271 20551
rect 9153 20460 9196 20506
rect 9242 20460 9271 20506
rect 9153 20338 9271 20460
rect 9153 20292 9196 20338
rect 9242 20292 9271 20338
rect 9153 20171 9271 20292
rect 9153 20125 9196 20171
rect 9242 20125 9271 20171
rect 9153 20003 9271 20125
rect 9153 19957 9196 20003
rect 9242 19957 9271 20003
rect 9153 19835 9271 19957
rect 9153 19789 9196 19835
rect 9242 19789 9271 19835
rect 9153 19667 9271 19789
rect 9153 19621 9196 19667
rect 9242 19621 9271 19667
rect 9153 19499 9271 19621
rect 9153 19453 9196 19499
rect 9242 19453 9271 19499
rect 9153 19332 9271 19453
rect 9153 19286 9196 19332
rect 9242 19286 9271 19332
rect 9153 19164 9271 19286
rect 9153 19118 9196 19164
rect 9242 19118 9271 19164
rect 9153 18996 9271 19118
rect 9153 18950 9196 18996
rect 9242 18950 9271 18996
rect 9153 18828 9271 18950
rect 9153 18782 9196 18828
rect 9242 18782 9271 18828
rect 9153 18658 9271 18782
rect 9153 18612 9196 18658
rect 9242 18612 9271 18658
rect 9153 18488 9271 18612
rect 9153 18442 9196 18488
rect 9242 18442 9271 18488
rect 9153 18318 9271 18442
rect 9153 18272 9196 18318
rect 9242 18272 9271 18318
rect 9153 18101 9271 18272
rect 9391 18101 9495 20551
rect 9615 20506 9734 20551
rect 9615 20460 9645 20506
rect 9691 20460 9734 20506
rect 9615 20338 9734 20460
rect 9615 20292 9645 20338
rect 9691 20292 9734 20338
rect 9615 20171 9734 20292
rect 9615 20125 9645 20171
rect 9691 20125 9734 20171
rect 9615 20003 9734 20125
rect 9615 19957 9645 20003
rect 9691 19957 9734 20003
rect 9615 19835 9734 19957
rect 9615 19789 9645 19835
rect 9691 19789 9734 19835
rect 9615 19667 9734 19789
rect 9615 19621 9645 19667
rect 9691 19621 9734 19667
rect 9615 19499 9734 19621
rect 9615 19453 9645 19499
rect 9691 19453 9734 19499
rect 9615 19332 9734 19453
rect 9615 19286 9645 19332
rect 9691 19286 9734 19332
rect 9615 19164 9734 19286
rect 9615 19118 9645 19164
rect 9691 19118 9734 19164
rect 9615 18996 9734 19118
rect 9615 18950 9645 18996
rect 9691 18950 9734 18996
rect 9615 18828 9734 18950
rect 9615 18782 9645 18828
rect 9691 18782 9734 18828
rect 9615 18658 9734 18782
rect 9615 18612 9645 18658
rect 9691 18612 9734 18658
rect 9615 18488 9734 18612
rect 9615 18442 9645 18488
rect 9691 18442 9734 18488
rect 9615 18318 9734 18442
rect 9615 18272 9645 18318
rect 9691 18272 9734 18318
rect 9615 18101 9734 18272
rect 10180 20506 10299 20551
rect 10180 20460 10223 20506
rect 10269 20460 10299 20506
rect 10180 20338 10299 20460
rect 10180 20292 10223 20338
rect 10269 20292 10299 20338
rect 10180 20171 10299 20292
rect 10180 20125 10223 20171
rect 10269 20125 10299 20171
rect 10180 20003 10299 20125
rect 10180 19957 10223 20003
rect 10269 19957 10299 20003
rect 10180 19835 10299 19957
rect 10180 19789 10223 19835
rect 10269 19789 10299 19835
rect 10180 19667 10299 19789
rect 10180 19621 10223 19667
rect 10269 19621 10299 19667
rect 10180 19499 10299 19621
rect 10180 19453 10223 19499
rect 10269 19453 10299 19499
rect 10180 19332 10299 19453
rect 10180 19286 10223 19332
rect 10269 19286 10299 19332
rect 10180 19164 10299 19286
rect 10180 19118 10223 19164
rect 10269 19118 10299 19164
rect 10180 18996 10299 19118
rect 10180 18950 10223 18996
rect 10269 18950 10299 18996
rect 10180 18828 10299 18950
rect 10180 18782 10223 18828
rect 10269 18782 10299 18828
rect 10180 18658 10299 18782
rect 10180 18612 10223 18658
rect 10269 18612 10299 18658
rect 10180 18488 10299 18612
rect 10180 18442 10223 18488
rect 10269 18442 10299 18488
rect 10180 18318 10299 18442
rect 10180 18272 10223 18318
rect 10269 18272 10299 18318
rect 10180 18101 10299 18272
rect 10419 18101 10523 20551
rect 10643 20506 10761 20551
rect 10643 20460 10672 20506
rect 10718 20460 10761 20506
rect 10643 20338 10761 20460
rect 10643 20292 10672 20338
rect 10718 20292 10761 20338
rect 10643 20171 10761 20292
rect 10643 20125 10672 20171
rect 10718 20125 10761 20171
rect 10643 20003 10761 20125
rect 10643 19957 10672 20003
rect 10718 19957 10761 20003
rect 10643 19835 10761 19957
rect 10643 19789 10672 19835
rect 10718 19789 10761 19835
rect 10643 19667 10761 19789
rect 10643 19621 10672 19667
rect 10718 19621 10761 19667
rect 10643 19499 10761 19621
rect 10643 19453 10672 19499
rect 10718 19453 10761 19499
rect 10643 19332 10761 19453
rect 10643 19286 10672 19332
rect 10718 19286 10761 19332
rect 10643 19164 10761 19286
rect 10643 19118 10672 19164
rect 10718 19118 10761 19164
rect 10643 18996 10761 19118
rect 10643 18950 10672 18996
rect 10718 18950 10761 18996
rect 10643 18828 10761 18950
rect 10643 18782 10672 18828
rect 10718 18782 10761 18828
rect 10643 18658 10761 18782
rect 10643 18612 10672 18658
rect 10718 18612 10761 18658
rect 10643 18488 10761 18612
rect 10643 18442 10672 18488
rect 10718 18442 10761 18488
rect 10643 18318 10761 18442
rect 10643 18272 10672 18318
rect 10718 18272 10761 18318
rect 10643 18101 10761 18272
rect 10945 20506 11063 20551
rect 10945 20460 10988 20506
rect 11034 20460 11063 20506
rect 10945 20338 11063 20460
rect 10945 20292 10988 20338
rect 11034 20292 11063 20338
rect 10945 20171 11063 20292
rect 10945 20125 10988 20171
rect 11034 20125 11063 20171
rect 10945 20003 11063 20125
rect 10945 19957 10988 20003
rect 11034 19957 11063 20003
rect 10945 19835 11063 19957
rect 10945 19789 10988 19835
rect 11034 19789 11063 19835
rect 10945 19667 11063 19789
rect 10945 19621 10988 19667
rect 11034 19621 11063 19667
rect 10945 19499 11063 19621
rect 10945 19453 10988 19499
rect 11034 19453 11063 19499
rect 10945 19332 11063 19453
rect 10945 19286 10988 19332
rect 11034 19286 11063 19332
rect 10945 19164 11063 19286
rect 10945 19118 10988 19164
rect 11034 19118 11063 19164
rect 10945 18996 11063 19118
rect 10945 18950 10988 18996
rect 11034 18950 11063 18996
rect 10945 18828 11063 18950
rect 10945 18782 10988 18828
rect 11034 18782 11063 18828
rect 10945 18658 11063 18782
rect 10945 18612 10988 18658
rect 11034 18612 11063 18658
rect 10945 18488 11063 18612
rect 10945 18442 10988 18488
rect 11034 18442 11063 18488
rect 10945 18318 11063 18442
rect 10945 18272 10988 18318
rect 11034 18272 11063 18318
rect 10945 18101 11063 18272
rect 11183 18101 11287 20551
rect 11407 20506 11526 20551
rect 11407 20460 11437 20506
rect 11483 20460 11526 20506
rect 11407 20338 11526 20460
rect 11407 20292 11437 20338
rect 11483 20292 11526 20338
rect 11407 20171 11526 20292
rect 11407 20125 11437 20171
rect 11483 20125 11526 20171
rect 11407 20003 11526 20125
rect 11407 19957 11437 20003
rect 11483 19957 11526 20003
rect 11407 19835 11526 19957
rect 11407 19789 11437 19835
rect 11483 19789 11526 19835
rect 11407 19667 11526 19789
rect 11407 19621 11437 19667
rect 11483 19621 11526 19667
rect 11407 19499 11526 19621
rect 11407 19453 11437 19499
rect 11483 19453 11526 19499
rect 11407 19332 11526 19453
rect 11407 19286 11437 19332
rect 11483 19286 11526 19332
rect 11407 19164 11526 19286
rect 11407 19118 11437 19164
rect 11483 19118 11526 19164
rect 11407 18996 11526 19118
rect 11407 18950 11437 18996
rect 11483 18950 11526 18996
rect 11407 18828 11526 18950
rect 11407 18782 11437 18828
rect 11483 18782 11526 18828
rect 11407 18658 11526 18782
rect 11407 18612 11437 18658
rect 11483 18612 11526 18658
rect 11407 18488 11526 18612
rect 11407 18442 11437 18488
rect 11483 18442 11526 18488
rect 11407 18318 11526 18442
rect 11407 18272 11437 18318
rect 11483 18272 11526 18318
rect 11407 18101 11526 18272
rect 11972 20506 12091 20551
rect 11972 20460 12015 20506
rect 12061 20460 12091 20506
rect 11972 20338 12091 20460
rect 11972 20292 12015 20338
rect 12061 20292 12091 20338
rect 11972 20171 12091 20292
rect 11972 20125 12015 20171
rect 12061 20125 12091 20171
rect 11972 20003 12091 20125
rect 11972 19957 12015 20003
rect 12061 19957 12091 20003
rect 11972 19835 12091 19957
rect 11972 19789 12015 19835
rect 12061 19789 12091 19835
rect 11972 19667 12091 19789
rect 11972 19621 12015 19667
rect 12061 19621 12091 19667
rect 11972 19499 12091 19621
rect 11972 19453 12015 19499
rect 12061 19453 12091 19499
rect 11972 19332 12091 19453
rect 11972 19286 12015 19332
rect 12061 19286 12091 19332
rect 11972 19164 12091 19286
rect 11972 19118 12015 19164
rect 12061 19118 12091 19164
rect 11972 18996 12091 19118
rect 11972 18950 12015 18996
rect 12061 18950 12091 18996
rect 11972 18828 12091 18950
rect 11972 18782 12015 18828
rect 12061 18782 12091 18828
rect 11972 18658 12091 18782
rect 11972 18612 12015 18658
rect 12061 18612 12091 18658
rect 11972 18488 12091 18612
rect 11972 18442 12015 18488
rect 12061 18442 12091 18488
rect 11972 18318 12091 18442
rect 11972 18272 12015 18318
rect 12061 18272 12091 18318
rect 11972 18101 12091 18272
rect 12211 18101 12315 20551
rect 12435 20506 12553 20551
rect 12435 20460 12464 20506
rect 12510 20460 12553 20506
rect 12435 20338 12553 20460
rect 12435 20292 12464 20338
rect 12510 20292 12553 20338
rect 12435 20171 12553 20292
rect 12435 20125 12464 20171
rect 12510 20125 12553 20171
rect 12435 20003 12553 20125
rect 12435 19957 12464 20003
rect 12510 19957 12553 20003
rect 12435 19835 12553 19957
rect 12435 19789 12464 19835
rect 12510 19789 12553 19835
rect 12435 19667 12553 19789
rect 12435 19621 12464 19667
rect 12510 19621 12553 19667
rect 12435 19499 12553 19621
rect 12435 19453 12464 19499
rect 12510 19453 12553 19499
rect 12435 19332 12553 19453
rect 12435 19286 12464 19332
rect 12510 19286 12553 19332
rect 12435 19164 12553 19286
rect 12435 19118 12464 19164
rect 12510 19118 12553 19164
rect 12435 18996 12553 19118
rect 12435 18950 12464 18996
rect 12510 18950 12553 18996
rect 12435 18828 12553 18950
rect 12435 18782 12464 18828
rect 12510 18782 12553 18828
rect 12435 18658 12553 18782
rect 12435 18612 12464 18658
rect 12510 18612 12553 18658
rect 12435 18488 12553 18612
rect 12435 18442 12464 18488
rect 12510 18442 12553 18488
rect 12435 18318 12553 18442
rect 12435 18272 12464 18318
rect 12510 18272 12553 18318
rect 12435 18101 12553 18272
rect 16661 20492 16779 20538
rect 16661 20446 16704 20492
rect 16750 20446 16779 20492
rect 16661 20325 16779 20446
rect 16661 20279 16704 20325
rect 16750 20279 16779 20325
rect 16661 20157 16779 20279
rect 16661 20111 16704 20157
rect 16750 20111 16779 20157
rect 16661 19989 16779 20111
rect 16661 19943 16704 19989
rect 16750 19943 16779 19989
rect 16661 19821 16779 19943
rect 16661 19775 16704 19821
rect 16750 19775 16779 19821
rect 16661 19654 16779 19775
rect 16661 19608 16704 19654
rect 16750 19608 16779 19654
rect 16661 19486 16779 19608
rect 16661 19440 16704 19486
rect 16750 19440 16779 19486
rect 16661 19318 16779 19440
rect 16661 19272 16704 19318
rect 16750 19272 16779 19318
rect 16661 19150 16779 19272
rect 16661 19104 16704 19150
rect 16750 19104 16779 19150
rect 16661 18982 16779 19104
rect 16661 18936 16704 18982
rect 16750 18936 16779 18982
rect 16661 18815 16779 18936
rect 16661 18769 16704 18815
rect 16750 18769 16779 18815
rect 16661 18645 16779 18769
rect 16661 18599 16704 18645
rect 16750 18599 16779 18645
rect 16661 18475 16779 18599
rect 16661 18429 16704 18475
rect 16750 18429 16779 18475
rect 16661 18305 16779 18429
rect 16661 18259 16704 18305
rect 16750 18259 16779 18305
rect 16661 18135 16779 18259
rect 16661 18089 16704 18135
rect 16750 18089 16779 18135
rect 16661 18043 16779 18089
rect 16899 18043 17003 20538
rect 17123 18043 17227 20538
rect 17347 20492 17451 20538
rect 17347 20446 17376 20492
rect 17422 20446 17451 20492
rect 17347 20325 17451 20446
rect 17347 20279 17376 20325
rect 17422 20279 17451 20325
rect 17347 20157 17451 20279
rect 17347 20111 17376 20157
rect 17422 20111 17451 20157
rect 17347 19989 17451 20111
rect 17347 19943 17376 19989
rect 17422 19943 17451 19989
rect 17347 19821 17451 19943
rect 17347 19775 17376 19821
rect 17422 19775 17451 19821
rect 17347 19654 17451 19775
rect 17347 19608 17376 19654
rect 17422 19608 17451 19654
rect 17347 19486 17451 19608
rect 17347 19440 17376 19486
rect 17422 19440 17451 19486
rect 17347 19318 17451 19440
rect 17347 19272 17376 19318
rect 17422 19272 17451 19318
rect 17347 19150 17451 19272
rect 17347 19104 17376 19150
rect 17422 19104 17451 19150
rect 17347 18982 17451 19104
rect 17347 18936 17376 18982
rect 17422 18936 17451 18982
rect 17347 18815 17451 18936
rect 17347 18769 17376 18815
rect 17422 18769 17451 18815
rect 17347 18645 17451 18769
rect 17347 18599 17376 18645
rect 17422 18599 17451 18645
rect 17347 18475 17451 18599
rect 17347 18429 17376 18475
rect 17422 18429 17451 18475
rect 17347 18305 17451 18429
rect 17347 18259 17376 18305
rect 17422 18259 17451 18305
rect 17347 18135 17451 18259
rect 17347 18089 17376 18135
rect 17422 18089 17451 18135
rect 17347 18043 17451 18089
rect 17571 18043 17675 20538
rect 17795 18043 17899 20538
rect 18019 20492 18137 20538
rect 18019 20446 18048 20492
rect 18094 20446 18137 20492
rect 18019 20325 18137 20446
rect 18019 20279 18048 20325
rect 18094 20279 18137 20325
rect 18019 20157 18137 20279
rect 18019 20111 18048 20157
rect 18094 20111 18137 20157
rect 18019 19989 18137 20111
rect 18019 19943 18048 19989
rect 18094 19943 18137 19989
rect 18019 19821 18137 19943
rect 18019 19775 18048 19821
rect 18094 19775 18137 19821
rect 18019 19654 18137 19775
rect 18019 19608 18048 19654
rect 18094 19608 18137 19654
rect 18019 19486 18137 19608
rect 18019 19440 18048 19486
rect 18094 19440 18137 19486
rect 18019 19318 18137 19440
rect 18019 19272 18048 19318
rect 18094 19272 18137 19318
rect 18019 19150 18137 19272
rect 18019 19104 18048 19150
rect 18094 19104 18137 19150
rect 18019 18982 18137 19104
rect 18019 18936 18048 18982
rect 18094 18936 18137 18982
rect 18019 18815 18137 18936
rect 18019 18769 18048 18815
rect 18094 18769 18137 18815
rect 18019 18645 18137 18769
rect 18019 18599 18048 18645
rect 18094 18599 18137 18645
rect 18019 18475 18137 18599
rect 18019 18429 18048 18475
rect 18094 18429 18137 18475
rect 18019 18305 18137 18429
rect 18019 18259 18048 18305
rect 18094 18259 18137 18305
rect 18019 18135 18137 18259
rect 18019 18089 18048 18135
rect 18094 18089 18137 18135
rect 18019 18043 18137 18089
rect 18295 20492 18413 20538
rect 18295 20446 18338 20492
rect 18384 20446 18413 20492
rect 18295 20325 18413 20446
rect 18295 20279 18338 20325
rect 18384 20279 18413 20325
rect 18295 20157 18413 20279
rect 18295 20111 18338 20157
rect 18384 20111 18413 20157
rect 18295 19989 18413 20111
rect 18295 19943 18338 19989
rect 18384 19943 18413 19989
rect 18295 19821 18413 19943
rect 18295 19775 18338 19821
rect 18384 19775 18413 19821
rect 18295 19654 18413 19775
rect 18295 19608 18338 19654
rect 18384 19608 18413 19654
rect 18295 19486 18413 19608
rect 18295 19440 18338 19486
rect 18384 19440 18413 19486
rect 18295 19318 18413 19440
rect 18295 19272 18338 19318
rect 18384 19272 18413 19318
rect 18295 19150 18413 19272
rect 18295 19104 18338 19150
rect 18384 19104 18413 19150
rect 18295 18982 18413 19104
rect 18295 18936 18338 18982
rect 18384 18936 18413 18982
rect 18295 18815 18413 18936
rect 18295 18769 18338 18815
rect 18384 18769 18413 18815
rect 18295 18645 18413 18769
rect 18295 18599 18338 18645
rect 18384 18599 18413 18645
rect 18295 18475 18413 18599
rect 18295 18429 18338 18475
rect 18384 18429 18413 18475
rect 18295 18305 18413 18429
rect 18295 18259 18338 18305
rect 18384 18259 18413 18305
rect 18295 18135 18413 18259
rect 18295 18089 18338 18135
rect 18384 18089 18413 18135
rect 18295 18043 18413 18089
rect 18533 18043 18637 20538
rect 18757 18043 18861 20538
rect 18981 20492 19085 20538
rect 18981 20446 19010 20492
rect 19056 20446 19085 20492
rect 18981 20325 19085 20446
rect 18981 20279 19010 20325
rect 19056 20279 19085 20325
rect 18981 20157 19085 20279
rect 18981 20111 19010 20157
rect 19056 20111 19085 20157
rect 18981 19989 19085 20111
rect 18981 19943 19010 19989
rect 19056 19943 19085 19989
rect 18981 19821 19085 19943
rect 18981 19775 19010 19821
rect 19056 19775 19085 19821
rect 18981 19654 19085 19775
rect 18981 19608 19010 19654
rect 19056 19608 19085 19654
rect 18981 19486 19085 19608
rect 18981 19440 19010 19486
rect 19056 19440 19085 19486
rect 18981 19318 19085 19440
rect 18981 19272 19010 19318
rect 19056 19272 19085 19318
rect 18981 19150 19085 19272
rect 18981 19104 19010 19150
rect 19056 19104 19085 19150
rect 18981 18982 19085 19104
rect 18981 18936 19010 18982
rect 19056 18936 19085 18982
rect 18981 18815 19085 18936
rect 18981 18769 19010 18815
rect 19056 18769 19085 18815
rect 18981 18645 19085 18769
rect 18981 18599 19010 18645
rect 19056 18599 19085 18645
rect 18981 18475 19085 18599
rect 18981 18429 19010 18475
rect 19056 18429 19085 18475
rect 18981 18305 19085 18429
rect 18981 18259 19010 18305
rect 19056 18259 19085 18305
rect 18981 18135 19085 18259
rect 18981 18089 19010 18135
rect 19056 18089 19085 18135
rect 18981 18043 19085 18089
rect 19205 18043 19309 20538
rect 19429 18043 19533 20538
rect 19653 20492 19771 20538
rect 19653 20446 19682 20492
rect 19728 20446 19771 20492
rect 19653 20325 19771 20446
rect 19653 20279 19682 20325
rect 19728 20279 19771 20325
rect 19653 20157 19771 20279
rect 19653 20111 19682 20157
rect 19728 20111 19771 20157
rect 19653 19989 19771 20111
rect 19653 19943 19682 19989
rect 19728 19943 19771 19989
rect 19653 19821 19771 19943
rect 19653 19775 19682 19821
rect 19728 19775 19771 19821
rect 19653 19654 19771 19775
rect 19653 19608 19682 19654
rect 19728 19608 19771 19654
rect 19653 19486 19771 19608
rect 19653 19440 19682 19486
rect 19728 19440 19771 19486
rect 19653 19318 19771 19440
rect 19653 19272 19682 19318
rect 19728 19272 19771 19318
rect 19653 19150 19771 19272
rect 19653 19104 19682 19150
rect 19728 19104 19771 19150
rect 19653 18982 19771 19104
rect 19653 18936 19682 18982
rect 19728 18936 19771 18982
rect 19653 18815 19771 18936
rect 19653 18769 19682 18815
rect 19728 18769 19771 18815
rect 19653 18645 19771 18769
rect 19653 18599 19682 18645
rect 19728 18599 19771 18645
rect 19653 18475 19771 18599
rect 19653 18429 19682 18475
rect 19728 18429 19771 18475
rect 19653 18305 19771 18429
rect 19653 18259 19682 18305
rect 19728 18259 19771 18305
rect 19653 18135 19771 18259
rect 19653 18089 19682 18135
rect 19728 18089 19771 18135
rect 19653 18043 19771 18089
rect 19928 20492 20046 20538
rect 19928 20446 19971 20492
rect 20017 20446 20046 20492
rect 19928 20325 20046 20446
rect 19928 20279 19971 20325
rect 20017 20279 20046 20325
rect 19928 20157 20046 20279
rect 19928 20111 19971 20157
rect 20017 20111 20046 20157
rect 19928 19989 20046 20111
rect 19928 19943 19971 19989
rect 20017 19943 20046 19989
rect 19928 19821 20046 19943
rect 19928 19775 19971 19821
rect 20017 19775 20046 19821
rect 19928 19654 20046 19775
rect 19928 19608 19971 19654
rect 20017 19608 20046 19654
rect 19928 19486 20046 19608
rect 19928 19440 19971 19486
rect 20017 19440 20046 19486
rect 19928 19318 20046 19440
rect 19928 19272 19971 19318
rect 20017 19272 20046 19318
rect 19928 19150 20046 19272
rect 19928 19104 19971 19150
rect 20017 19104 20046 19150
rect 19928 18982 20046 19104
rect 19928 18936 19971 18982
rect 20017 18936 20046 18982
rect 19928 18815 20046 18936
rect 19928 18769 19971 18815
rect 20017 18769 20046 18815
rect 19928 18645 20046 18769
rect 19928 18599 19971 18645
rect 20017 18599 20046 18645
rect 19928 18475 20046 18599
rect 19928 18429 19971 18475
rect 20017 18429 20046 18475
rect 19928 18305 20046 18429
rect 19928 18259 19971 18305
rect 20017 18259 20046 18305
rect 19928 18135 20046 18259
rect 19928 18089 19971 18135
rect 20017 18089 20046 18135
rect 19928 18043 20046 18089
rect 20166 18043 20270 20538
rect 20390 18043 20494 20538
rect 20614 20492 20718 20538
rect 20614 20446 20643 20492
rect 20689 20446 20718 20492
rect 20614 20325 20718 20446
rect 20614 20279 20643 20325
rect 20689 20279 20718 20325
rect 20614 20157 20718 20279
rect 20614 20111 20643 20157
rect 20689 20111 20718 20157
rect 20614 19989 20718 20111
rect 20614 19943 20643 19989
rect 20689 19943 20718 19989
rect 20614 19821 20718 19943
rect 20614 19775 20643 19821
rect 20689 19775 20718 19821
rect 20614 19654 20718 19775
rect 20614 19608 20643 19654
rect 20689 19608 20718 19654
rect 20614 19486 20718 19608
rect 20614 19440 20643 19486
rect 20689 19440 20718 19486
rect 20614 19318 20718 19440
rect 20614 19272 20643 19318
rect 20689 19272 20718 19318
rect 20614 19150 20718 19272
rect 20614 19104 20643 19150
rect 20689 19104 20718 19150
rect 20614 18982 20718 19104
rect 20614 18936 20643 18982
rect 20689 18936 20718 18982
rect 20614 18815 20718 18936
rect 20614 18769 20643 18815
rect 20689 18769 20718 18815
rect 20614 18645 20718 18769
rect 20614 18599 20643 18645
rect 20689 18599 20718 18645
rect 20614 18475 20718 18599
rect 20614 18429 20643 18475
rect 20689 18429 20718 18475
rect 20614 18305 20718 18429
rect 20614 18259 20643 18305
rect 20689 18259 20718 18305
rect 20614 18135 20718 18259
rect 20614 18089 20643 18135
rect 20689 18089 20718 18135
rect 20614 18043 20718 18089
rect 20838 18043 20942 20538
rect 21062 18043 21166 20538
rect 21286 20492 21404 20538
rect 21286 20446 21315 20492
rect 21361 20446 21404 20492
rect 21286 20325 21404 20446
rect 21286 20279 21315 20325
rect 21361 20279 21404 20325
rect 21286 20157 21404 20279
rect 21286 20111 21315 20157
rect 21361 20111 21404 20157
rect 21286 19989 21404 20111
rect 21286 19943 21315 19989
rect 21361 19943 21404 19989
rect 21286 19821 21404 19943
rect 21286 19775 21315 19821
rect 21361 19775 21404 19821
rect 21286 19654 21404 19775
rect 21286 19608 21315 19654
rect 21361 19608 21404 19654
rect 21286 19486 21404 19608
rect 21286 19440 21315 19486
rect 21361 19440 21404 19486
rect 21286 19318 21404 19440
rect 21286 19272 21315 19318
rect 21361 19272 21404 19318
rect 21286 19150 21404 19272
rect 21286 19104 21315 19150
rect 21361 19104 21404 19150
rect 21286 18982 21404 19104
rect 21286 18936 21315 18982
rect 21361 18936 21404 18982
rect 21286 18815 21404 18936
rect 21286 18769 21315 18815
rect 21361 18769 21404 18815
rect 21286 18645 21404 18769
rect 21286 18599 21315 18645
rect 21361 18599 21404 18645
rect 21286 18475 21404 18599
rect 21286 18429 21315 18475
rect 21361 18429 21404 18475
rect 21286 18305 21404 18429
rect 21286 18259 21315 18305
rect 21361 18259 21404 18305
rect 21286 18135 21404 18259
rect 21286 18089 21315 18135
rect 21361 18089 21404 18135
rect 21286 18043 21404 18089
rect 21562 20492 21680 20538
rect 21562 20446 21605 20492
rect 21651 20446 21680 20492
rect 21562 20325 21680 20446
rect 21562 20279 21605 20325
rect 21651 20279 21680 20325
rect 21562 20157 21680 20279
rect 21562 20111 21605 20157
rect 21651 20111 21680 20157
rect 21562 19989 21680 20111
rect 21562 19943 21605 19989
rect 21651 19943 21680 19989
rect 21562 19821 21680 19943
rect 21562 19775 21605 19821
rect 21651 19775 21680 19821
rect 21562 19654 21680 19775
rect 21562 19608 21605 19654
rect 21651 19608 21680 19654
rect 21562 19486 21680 19608
rect 21562 19440 21605 19486
rect 21651 19440 21680 19486
rect 21562 19318 21680 19440
rect 21562 19272 21605 19318
rect 21651 19272 21680 19318
rect 21562 19150 21680 19272
rect 21562 19104 21605 19150
rect 21651 19104 21680 19150
rect 21562 18982 21680 19104
rect 21562 18936 21605 18982
rect 21651 18936 21680 18982
rect 21562 18815 21680 18936
rect 21562 18769 21605 18815
rect 21651 18769 21680 18815
rect 21562 18645 21680 18769
rect 21562 18599 21605 18645
rect 21651 18599 21680 18645
rect 21562 18475 21680 18599
rect 21562 18429 21605 18475
rect 21651 18429 21680 18475
rect 21562 18305 21680 18429
rect 21562 18259 21605 18305
rect 21651 18259 21680 18305
rect 21562 18135 21680 18259
rect 21562 18089 21605 18135
rect 21651 18089 21680 18135
rect 21562 18043 21680 18089
rect 21800 18043 21904 20538
rect 22024 18043 22128 20538
rect 22248 20492 22352 20538
rect 22248 20446 22277 20492
rect 22323 20446 22352 20492
rect 22248 20325 22352 20446
rect 22248 20279 22277 20325
rect 22323 20279 22352 20325
rect 22248 20157 22352 20279
rect 22248 20111 22277 20157
rect 22323 20111 22352 20157
rect 22248 19989 22352 20111
rect 22248 19943 22277 19989
rect 22323 19943 22352 19989
rect 22248 19821 22352 19943
rect 22248 19775 22277 19821
rect 22323 19775 22352 19821
rect 22248 19654 22352 19775
rect 22248 19608 22277 19654
rect 22323 19608 22352 19654
rect 22248 19486 22352 19608
rect 22248 19440 22277 19486
rect 22323 19440 22352 19486
rect 22248 19318 22352 19440
rect 22248 19272 22277 19318
rect 22323 19272 22352 19318
rect 22248 19150 22352 19272
rect 22248 19104 22277 19150
rect 22323 19104 22352 19150
rect 22248 18982 22352 19104
rect 22248 18936 22277 18982
rect 22323 18936 22352 18982
rect 22248 18815 22352 18936
rect 22248 18769 22277 18815
rect 22323 18769 22352 18815
rect 22248 18645 22352 18769
rect 22248 18599 22277 18645
rect 22323 18599 22352 18645
rect 22248 18475 22352 18599
rect 22248 18429 22277 18475
rect 22323 18429 22352 18475
rect 22248 18305 22352 18429
rect 22248 18259 22277 18305
rect 22323 18259 22352 18305
rect 22248 18135 22352 18259
rect 22248 18089 22277 18135
rect 22323 18089 22352 18135
rect 22248 18043 22352 18089
rect 22472 18043 22576 20538
rect 22696 18043 22800 20538
rect 22920 20492 23038 20538
rect 22920 20446 22949 20492
rect 22995 20446 23038 20492
rect 22920 20325 23038 20446
rect 22920 20279 22949 20325
rect 22995 20279 23038 20325
rect 22920 20157 23038 20279
rect 22920 20111 22949 20157
rect 22995 20111 23038 20157
rect 22920 19989 23038 20111
rect 22920 19943 22949 19989
rect 22995 19943 23038 19989
rect 22920 19821 23038 19943
rect 22920 19775 22949 19821
rect 22995 19775 23038 19821
rect 22920 19654 23038 19775
rect 22920 19608 22949 19654
rect 22995 19608 23038 19654
rect 22920 19486 23038 19608
rect 22920 19440 22949 19486
rect 22995 19440 23038 19486
rect 22920 19318 23038 19440
rect 22920 19272 22949 19318
rect 22995 19272 23038 19318
rect 22920 19150 23038 19272
rect 22920 19104 22949 19150
rect 22995 19104 23038 19150
rect 22920 18982 23038 19104
rect 22920 18936 22949 18982
rect 22995 18936 23038 18982
rect 22920 18815 23038 18936
rect 22920 18769 22949 18815
rect 22995 18769 23038 18815
rect 22920 18645 23038 18769
rect 22920 18599 22949 18645
rect 22995 18599 23038 18645
rect 22920 18475 23038 18599
rect 22920 18429 22949 18475
rect 22995 18429 23038 18475
rect 22920 18305 23038 18429
rect 22920 18259 22949 18305
rect 22995 18259 23038 18305
rect 22920 18135 23038 18259
rect 22920 18089 22949 18135
rect 22995 18089 23038 18135
rect 22920 18043 23038 18089
rect 1982 11757 2070 11770
rect 1982 10997 1995 11757
rect 2041 10997 2070 11757
rect 1982 10940 2070 10997
rect 1982 10894 1995 10940
rect 2041 10894 2070 10940
rect 1982 10837 2070 10894
rect 1982 10791 1995 10837
rect 2041 10791 2070 10837
rect 1982 10734 2070 10791
rect 1982 10688 1995 10734
rect 2041 10688 2070 10734
rect 1982 10631 2070 10688
rect 1982 10585 1995 10631
rect 2041 10585 2070 10631
rect 1982 10528 2070 10585
rect 1982 10482 1995 10528
rect 2041 10482 2070 10528
rect 1982 10425 2070 10482
rect 1982 10379 1995 10425
rect 2041 10379 2070 10425
rect 1982 10322 2070 10379
rect 1982 10276 1995 10322
rect 2041 10276 2070 10322
rect 1982 10219 2070 10276
rect 1982 10173 1995 10219
rect 2041 10173 2070 10219
rect 1982 10116 2070 10173
rect 1982 10070 1995 10116
rect 2041 10070 2070 10116
rect 1982 10013 2070 10070
rect 1982 9967 1995 10013
rect 2041 9967 2070 10013
rect 1982 9954 2070 9967
rect 2190 11757 2278 11770
rect 2190 10997 2219 11757
rect 2265 10997 2278 11757
rect 2190 10940 2278 10997
rect 2190 10894 2219 10940
rect 2265 10894 2278 10940
rect 2190 10837 2278 10894
rect 2190 10791 2219 10837
rect 2265 10791 2278 10837
rect 2190 10734 2278 10791
rect 2190 10688 2219 10734
rect 2265 10688 2278 10734
rect 2190 10631 2278 10688
rect 2190 10585 2219 10631
rect 2265 10585 2278 10631
rect 2190 10528 2278 10585
rect 2190 10482 2219 10528
rect 2265 10482 2278 10528
rect 2190 10425 2278 10482
rect 2190 10379 2219 10425
rect 2265 10379 2278 10425
rect 2190 10322 2278 10379
rect 2190 10276 2219 10322
rect 2265 10276 2278 10322
rect 2190 10219 2278 10276
rect 2190 10173 2219 10219
rect 2265 10173 2278 10219
rect 2190 10116 2278 10173
rect 2190 10070 2219 10116
rect 2265 10070 2278 10116
rect 2190 10013 2278 10070
rect 2190 9967 2219 10013
rect 2265 9967 2278 10013
rect 2190 9954 2278 9967
rect 2430 11757 2518 11770
rect 2430 10997 2443 11757
rect 2489 10997 2518 11757
rect 2430 10940 2518 10997
rect 2430 10894 2443 10940
rect 2489 10894 2518 10940
rect 2430 10837 2518 10894
rect 2430 10791 2443 10837
rect 2489 10791 2518 10837
rect 2430 10734 2518 10791
rect 2430 10688 2443 10734
rect 2489 10688 2518 10734
rect 2430 10631 2518 10688
rect 2430 10585 2443 10631
rect 2489 10585 2518 10631
rect 2430 10528 2518 10585
rect 2430 10482 2443 10528
rect 2489 10482 2518 10528
rect 2430 10425 2518 10482
rect 2430 10379 2443 10425
rect 2489 10379 2518 10425
rect 2430 10322 2518 10379
rect 2430 10276 2443 10322
rect 2489 10276 2518 10322
rect 2430 10219 2518 10276
rect 2430 10173 2443 10219
rect 2489 10173 2518 10219
rect 2430 10116 2518 10173
rect 2430 10070 2443 10116
rect 2489 10070 2518 10116
rect 2430 10013 2518 10070
rect 2430 9967 2443 10013
rect 2489 9967 2518 10013
rect 2430 9954 2518 9967
rect 2638 11757 2742 11770
rect 2638 10997 2667 11757
rect 2713 10997 2742 11757
rect 2638 10940 2742 10997
rect 2638 10894 2667 10940
rect 2713 10894 2742 10940
rect 2638 10837 2742 10894
rect 2638 10791 2667 10837
rect 2713 10791 2742 10837
rect 2638 10734 2742 10791
rect 2638 10688 2667 10734
rect 2713 10688 2742 10734
rect 2638 10631 2742 10688
rect 2638 10585 2667 10631
rect 2713 10585 2742 10631
rect 2638 10528 2742 10585
rect 2638 10482 2667 10528
rect 2713 10482 2742 10528
rect 2638 10425 2742 10482
rect 2638 10379 2667 10425
rect 2713 10379 2742 10425
rect 2638 10322 2742 10379
rect 2638 10276 2667 10322
rect 2713 10276 2742 10322
rect 2638 10219 2742 10276
rect 2638 10173 2667 10219
rect 2713 10173 2742 10219
rect 2638 10116 2742 10173
rect 2638 10070 2667 10116
rect 2713 10070 2742 10116
rect 2638 10013 2742 10070
rect 2638 9967 2667 10013
rect 2713 9967 2742 10013
rect 2638 9954 2742 9967
rect 2862 11757 2966 11770
rect 2862 10997 2891 11757
rect 2937 10997 2966 11757
rect 2862 10940 2966 10997
rect 2862 10894 2891 10940
rect 2937 10894 2966 10940
rect 2862 10837 2966 10894
rect 2862 10791 2891 10837
rect 2937 10791 2966 10837
rect 2862 10734 2966 10791
rect 2862 10688 2891 10734
rect 2937 10688 2966 10734
rect 2862 10631 2966 10688
rect 2862 10585 2891 10631
rect 2937 10585 2966 10631
rect 2862 10528 2966 10585
rect 2862 10482 2891 10528
rect 2937 10482 2966 10528
rect 2862 10425 2966 10482
rect 2862 10379 2891 10425
rect 2937 10379 2966 10425
rect 2862 10322 2966 10379
rect 2862 10276 2891 10322
rect 2937 10276 2966 10322
rect 2862 10219 2966 10276
rect 2862 10173 2891 10219
rect 2937 10173 2966 10219
rect 2862 10116 2966 10173
rect 2862 10070 2891 10116
rect 2937 10070 2966 10116
rect 2862 10013 2966 10070
rect 2862 9967 2891 10013
rect 2937 9967 2966 10013
rect 2862 9954 2966 9967
rect 3086 11757 3190 11770
rect 3086 10997 3115 11757
rect 3161 10997 3190 11757
rect 3086 10940 3190 10997
rect 3086 10894 3115 10940
rect 3161 10894 3190 10940
rect 3086 10837 3190 10894
rect 3086 10791 3115 10837
rect 3161 10791 3190 10837
rect 3086 10734 3190 10791
rect 3086 10688 3115 10734
rect 3161 10688 3190 10734
rect 3086 10631 3190 10688
rect 3086 10585 3115 10631
rect 3161 10585 3190 10631
rect 3086 10528 3190 10585
rect 3086 10482 3115 10528
rect 3161 10482 3190 10528
rect 3086 10425 3190 10482
rect 3086 10379 3115 10425
rect 3161 10379 3190 10425
rect 3086 10322 3190 10379
rect 3086 10276 3115 10322
rect 3161 10276 3190 10322
rect 3086 10219 3190 10276
rect 3086 10173 3115 10219
rect 3161 10173 3190 10219
rect 3086 10116 3190 10173
rect 3086 10070 3115 10116
rect 3161 10070 3190 10116
rect 3086 10013 3190 10070
rect 3086 9967 3115 10013
rect 3161 9967 3190 10013
rect 3086 9954 3190 9967
rect 3310 11757 3398 11770
rect 3310 10997 3339 11757
rect 3385 10997 3398 11757
rect 3310 10940 3398 10997
rect 3310 10894 3339 10940
rect 3385 10894 3398 10940
rect 3310 10837 3398 10894
rect 3310 10791 3339 10837
rect 3385 10791 3398 10837
rect 3310 10734 3398 10791
rect 3310 10688 3339 10734
rect 3385 10688 3398 10734
rect 3310 10631 3398 10688
rect 3310 10585 3339 10631
rect 3385 10585 3398 10631
rect 3310 10528 3398 10585
rect 3310 10482 3339 10528
rect 3385 10482 3398 10528
rect 3310 10425 3398 10482
rect 3310 10379 3339 10425
rect 3385 10379 3398 10425
rect 3310 10322 3398 10379
rect 3310 10276 3339 10322
rect 3385 10276 3398 10322
rect 3310 10219 3398 10276
rect 3310 10173 3339 10219
rect 3385 10173 3398 10219
rect 3310 10116 3398 10173
rect 3310 10070 3339 10116
rect 3385 10070 3398 10116
rect 3310 10013 3398 10070
rect 3310 9967 3339 10013
rect 3385 9967 3398 10013
rect 3310 9954 3398 9967
rect 3550 11757 3638 11770
rect 3550 10997 3563 11757
rect 3609 10997 3638 11757
rect 3550 10940 3638 10997
rect 3550 10894 3563 10940
rect 3609 10894 3638 10940
rect 3550 10837 3638 10894
rect 3550 10791 3563 10837
rect 3609 10791 3638 10837
rect 3550 10734 3638 10791
rect 3550 10688 3563 10734
rect 3609 10688 3638 10734
rect 3550 10631 3638 10688
rect 3550 10585 3563 10631
rect 3609 10585 3638 10631
rect 3550 10528 3638 10585
rect 3550 10482 3563 10528
rect 3609 10482 3638 10528
rect 3550 10425 3638 10482
rect 3550 10379 3563 10425
rect 3609 10379 3638 10425
rect 3550 10322 3638 10379
rect 3550 10276 3563 10322
rect 3609 10276 3638 10322
rect 3550 10219 3638 10276
rect 3550 10173 3563 10219
rect 3609 10173 3638 10219
rect 3550 10116 3638 10173
rect 3550 10070 3563 10116
rect 3609 10070 3638 10116
rect 3550 10013 3638 10070
rect 3550 9967 3563 10013
rect 3609 9967 3638 10013
rect 3550 9954 3638 9967
rect 3758 11757 3862 11770
rect 3758 10997 3787 11757
rect 3833 10997 3862 11757
rect 3758 10940 3862 10997
rect 3758 10894 3787 10940
rect 3833 10894 3862 10940
rect 3758 10837 3862 10894
rect 3758 10791 3787 10837
rect 3833 10791 3862 10837
rect 3758 10734 3862 10791
rect 3758 10688 3787 10734
rect 3833 10688 3862 10734
rect 3758 10631 3862 10688
rect 3758 10585 3787 10631
rect 3833 10585 3862 10631
rect 3758 10528 3862 10585
rect 3758 10482 3787 10528
rect 3833 10482 3862 10528
rect 3758 10425 3862 10482
rect 3758 10379 3787 10425
rect 3833 10379 3862 10425
rect 3758 10322 3862 10379
rect 3758 10276 3787 10322
rect 3833 10276 3862 10322
rect 3758 10219 3862 10276
rect 3758 10173 3787 10219
rect 3833 10173 3862 10219
rect 3758 10116 3862 10173
rect 3758 10070 3787 10116
rect 3833 10070 3862 10116
rect 3758 10013 3862 10070
rect 3758 9967 3787 10013
rect 3833 9967 3862 10013
rect 3758 9954 3862 9967
rect 3982 11757 4086 11770
rect 3982 10997 4011 11757
rect 4057 10997 4086 11757
rect 3982 10940 4086 10997
rect 3982 10894 4011 10940
rect 4057 10894 4086 10940
rect 3982 10837 4086 10894
rect 3982 10791 4011 10837
rect 4057 10791 4086 10837
rect 3982 10734 4086 10791
rect 3982 10688 4011 10734
rect 4057 10688 4086 10734
rect 3982 10631 4086 10688
rect 3982 10585 4011 10631
rect 4057 10585 4086 10631
rect 3982 10528 4086 10585
rect 3982 10482 4011 10528
rect 4057 10482 4086 10528
rect 3982 10425 4086 10482
rect 3982 10379 4011 10425
rect 4057 10379 4086 10425
rect 3982 10322 4086 10379
rect 3982 10276 4011 10322
rect 4057 10276 4086 10322
rect 3982 10219 4086 10276
rect 3982 10173 4011 10219
rect 4057 10173 4086 10219
rect 3982 10116 4086 10173
rect 3982 10070 4011 10116
rect 4057 10070 4086 10116
rect 3982 10013 4086 10070
rect 3982 9967 4011 10013
rect 4057 9967 4086 10013
rect 3982 9954 4086 9967
rect 4206 11757 4310 11770
rect 4206 10997 4235 11757
rect 4281 10997 4310 11757
rect 4206 10940 4310 10997
rect 4206 10894 4235 10940
rect 4281 10894 4310 10940
rect 4206 10837 4310 10894
rect 4206 10791 4235 10837
rect 4281 10791 4310 10837
rect 4206 10734 4310 10791
rect 4206 10688 4235 10734
rect 4281 10688 4310 10734
rect 4206 10631 4310 10688
rect 4206 10585 4235 10631
rect 4281 10585 4310 10631
rect 4206 10528 4310 10585
rect 4206 10482 4235 10528
rect 4281 10482 4310 10528
rect 4206 10425 4310 10482
rect 4206 10379 4235 10425
rect 4281 10379 4310 10425
rect 4206 10322 4310 10379
rect 4206 10276 4235 10322
rect 4281 10276 4310 10322
rect 4206 10219 4310 10276
rect 4206 10173 4235 10219
rect 4281 10173 4310 10219
rect 4206 10116 4310 10173
rect 4206 10070 4235 10116
rect 4281 10070 4310 10116
rect 4206 10013 4310 10070
rect 4206 9967 4235 10013
rect 4281 9967 4310 10013
rect 4206 9954 4310 9967
rect 4430 11757 4518 11770
rect 4430 10997 4459 11757
rect 4505 10997 4518 11757
rect 4430 10940 4518 10997
rect 4430 10894 4459 10940
rect 4505 10894 4518 10940
rect 4430 10837 4518 10894
rect 4430 10791 4459 10837
rect 4505 10791 4518 10837
rect 4430 10734 4518 10791
rect 4430 10688 4459 10734
rect 4505 10688 4518 10734
rect 4430 10631 4518 10688
rect 4430 10585 4459 10631
rect 4505 10585 4518 10631
rect 4430 10528 4518 10585
rect 4430 10482 4459 10528
rect 4505 10482 4518 10528
rect 4430 10425 4518 10482
rect 4430 10379 4459 10425
rect 4505 10379 4518 10425
rect 4430 10322 4518 10379
rect 4430 10276 4459 10322
rect 4505 10276 4518 10322
rect 4430 10219 4518 10276
rect 4430 10173 4459 10219
rect 4505 10173 4518 10219
rect 4430 10116 4518 10173
rect 4430 10070 4459 10116
rect 4505 10070 4518 10116
rect 4430 10013 4518 10070
rect 4430 9967 4459 10013
rect 4505 9967 4518 10013
rect 4430 9954 4518 9967
rect 4670 11757 4758 11770
rect 4670 10997 4683 11757
rect 4729 10997 4758 11757
rect 4670 10940 4758 10997
rect 4670 10894 4683 10940
rect 4729 10894 4758 10940
rect 4670 10837 4758 10894
rect 4670 10791 4683 10837
rect 4729 10791 4758 10837
rect 4670 10734 4758 10791
rect 4670 10688 4683 10734
rect 4729 10688 4758 10734
rect 4670 10631 4758 10688
rect 4670 10585 4683 10631
rect 4729 10585 4758 10631
rect 4670 10528 4758 10585
rect 4670 10482 4683 10528
rect 4729 10482 4758 10528
rect 4670 10425 4758 10482
rect 4670 10379 4683 10425
rect 4729 10379 4758 10425
rect 4670 10322 4758 10379
rect 4670 10276 4683 10322
rect 4729 10276 4758 10322
rect 4670 10219 4758 10276
rect 4670 10173 4683 10219
rect 4729 10173 4758 10219
rect 4670 10116 4758 10173
rect 4670 10070 4683 10116
rect 4729 10070 4758 10116
rect 4670 10013 4758 10070
rect 4670 9967 4683 10013
rect 4729 9967 4758 10013
rect 4670 9954 4758 9967
rect 4878 11757 4982 11770
rect 4878 10997 4907 11757
rect 4953 10997 4982 11757
rect 4878 10940 4982 10997
rect 4878 10894 4907 10940
rect 4953 10894 4982 10940
rect 4878 10837 4982 10894
rect 4878 10791 4907 10837
rect 4953 10791 4982 10837
rect 4878 10734 4982 10791
rect 4878 10688 4907 10734
rect 4953 10688 4982 10734
rect 4878 10631 4982 10688
rect 4878 10585 4907 10631
rect 4953 10585 4982 10631
rect 4878 10528 4982 10585
rect 4878 10482 4907 10528
rect 4953 10482 4982 10528
rect 4878 10425 4982 10482
rect 4878 10379 4907 10425
rect 4953 10379 4982 10425
rect 4878 10322 4982 10379
rect 4878 10276 4907 10322
rect 4953 10276 4982 10322
rect 4878 10219 4982 10276
rect 4878 10173 4907 10219
rect 4953 10173 4982 10219
rect 4878 10116 4982 10173
rect 4878 10070 4907 10116
rect 4953 10070 4982 10116
rect 4878 10013 4982 10070
rect 4878 9967 4907 10013
rect 4953 9967 4982 10013
rect 4878 9954 4982 9967
rect 5102 11757 5206 11770
rect 5102 10997 5131 11757
rect 5177 10997 5206 11757
rect 5102 10940 5206 10997
rect 5102 10894 5131 10940
rect 5177 10894 5206 10940
rect 5102 10837 5206 10894
rect 5102 10791 5131 10837
rect 5177 10791 5206 10837
rect 5102 10734 5206 10791
rect 5102 10688 5131 10734
rect 5177 10688 5206 10734
rect 5102 10631 5206 10688
rect 5102 10585 5131 10631
rect 5177 10585 5206 10631
rect 5102 10528 5206 10585
rect 5102 10482 5131 10528
rect 5177 10482 5206 10528
rect 5102 10425 5206 10482
rect 5102 10379 5131 10425
rect 5177 10379 5206 10425
rect 5102 10322 5206 10379
rect 5102 10276 5131 10322
rect 5177 10276 5206 10322
rect 5102 10219 5206 10276
rect 5102 10173 5131 10219
rect 5177 10173 5206 10219
rect 5102 10116 5206 10173
rect 5102 10070 5131 10116
rect 5177 10070 5206 10116
rect 5102 10013 5206 10070
rect 5102 9967 5131 10013
rect 5177 9967 5206 10013
rect 5102 9954 5206 9967
rect 5326 11757 5430 11770
rect 5326 10997 5355 11757
rect 5401 10997 5430 11757
rect 5326 10940 5430 10997
rect 5326 10894 5355 10940
rect 5401 10894 5430 10940
rect 5326 10837 5430 10894
rect 5326 10791 5355 10837
rect 5401 10791 5430 10837
rect 5326 10734 5430 10791
rect 5326 10688 5355 10734
rect 5401 10688 5430 10734
rect 5326 10631 5430 10688
rect 5326 10585 5355 10631
rect 5401 10585 5430 10631
rect 5326 10528 5430 10585
rect 5326 10482 5355 10528
rect 5401 10482 5430 10528
rect 5326 10425 5430 10482
rect 5326 10379 5355 10425
rect 5401 10379 5430 10425
rect 5326 10322 5430 10379
rect 5326 10276 5355 10322
rect 5401 10276 5430 10322
rect 5326 10219 5430 10276
rect 5326 10173 5355 10219
rect 5401 10173 5430 10219
rect 5326 10116 5430 10173
rect 5326 10070 5355 10116
rect 5401 10070 5430 10116
rect 5326 10013 5430 10070
rect 5326 9967 5355 10013
rect 5401 9967 5430 10013
rect 5326 9954 5430 9967
rect 5550 11757 5638 11770
rect 5550 10997 5579 11757
rect 5625 10997 5638 11757
rect 5550 10940 5638 10997
rect 5550 10894 5579 10940
rect 5625 10894 5638 10940
rect 5550 10837 5638 10894
rect 5550 10791 5579 10837
rect 5625 10791 5638 10837
rect 5550 10734 5638 10791
rect 5550 10688 5579 10734
rect 5625 10688 5638 10734
rect 5550 10631 5638 10688
rect 5550 10585 5579 10631
rect 5625 10585 5638 10631
rect 5550 10528 5638 10585
rect 5550 10482 5579 10528
rect 5625 10482 5638 10528
rect 5550 10425 5638 10482
rect 5550 10379 5579 10425
rect 5625 10379 5638 10425
rect 5550 10322 5638 10379
rect 5550 10276 5579 10322
rect 5625 10276 5638 10322
rect 5550 10219 5638 10276
rect 5550 10173 5579 10219
rect 5625 10173 5638 10219
rect 5550 10116 5638 10173
rect 5550 10070 5579 10116
rect 5625 10070 5638 10116
rect 5550 10013 5638 10070
rect 5550 9967 5579 10013
rect 5625 9967 5638 10013
rect 5550 9954 5638 9967
rect 5790 11757 5878 11770
rect 5790 10997 5803 11757
rect 5849 10997 5878 11757
rect 5790 10940 5878 10997
rect 5790 10894 5803 10940
rect 5849 10894 5878 10940
rect 5790 10837 5878 10894
rect 5790 10791 5803 10837
rect 5849 10791 5878 10837
rect 5790 10734 5878 10791
rect 5790 10688 5803 10734
rect 5849 10688 5878 10734
rect 5790 10631 5878 10688
rect 5790 10585 5803 10631
rect 5849 10585 5878 10631
rect 5790 10528 5878 10585
rect 5790 10482 5803 10528
rect 5849 10482 5878 10528
rect 5790 10425 5878 10482
rect 5790 10379 5803 10425
rect 5849 10379 5878 10425
rect 5790 10322 5878 10379
rect 5790 10276 5803 10322
rect 5849 10276 5878 10322
rect 5790 10219 5878 10276
rect 5790 10173 5803 10219
rect 5849 10173 5878 10219
rect 5790 10116 5878 10173
rect 5790 10070 5803 10116
rect 5849 10070 5878 10116
rect 5790 10013 5878 10070
rect 5790 9967 5803 10013
rect 5849 9967 5878 10013
rect 5790 9954 5878 9967
rect 5998 11757 6102 11770
rect 5998 10997 6027 11757
rect 6073 10997 6102 11757
rect 5998 10940 6102 10997
rect 5998 10894 6027 10940
rect 6073 10894 6102 10940
rect 5998 10837 6102 10894
rect 5998 10791 6027 10837
rect 6073 10791 6102 10837
rect 5998 10734 6102 10791
rect 5998 10688 6027 10734
rect 6073 10688 6102 10734
rect 5998 10631 6102 10688
rect 5998 10585 6027 10631
rect 6073 10585 6102 10631
rect 5998 10528 6102 10585
rect 5998 10482 6027 10528
rect 6073 10482 6102 10528
rect 5998 10425 6102 10482
rect 5998 10379 6027 10425
rect 6073 10379 6102 10425
rect 5998 10322 6102 10379
rect 5998 10276 6027 10322
rect 6073 10276 6102 10322
rect 5998 10219 6102 10276
rect 5998 10173 6027 10219
rect 6073 10173 6102 10219
rect 5998 10116 6102 10173
rect 5998 10070 6027 10116
rect 6073 10070 6102 10116
rect 5998 10013 6102 10070
rect 5998 9967 6027 10013
rect 6073 9967 6102 10013
rect 5998 9954 6102 9967
rect 6222 11757 6326 11770
rect 6222 10997 6251 11757
rect 6297 10997 6326 11757
rect 6222 10940 6326 10997
rect 6222 10894 6251 10940
rect 6297 10894 6326 10940
rect 6222 10837 6326 10894
rect 6222 10791 6251 10837
rect 6297 10791 6326 10837
rect 6222 10734 6326 10791
rect 6222 10688 6251 10734
rect 6297 10688 6326 10734
rect 6222 10631 6326 10688
rect 6222 10585 6251 10631
rect 6297 10585 6326 10631
rect 6222 10528 6326 10585
rect 6222 10482 6251 10528
rect 6297 10482 6326 10528
rect 6222 10425 6326 10482
rect 6222 10379 6251 10425
rect 6297 10379 6326 10425
rect 6222 10322 6326 10379
rect 6222 10276 6251 10322
rect 6297 10276 6326 10322
rect 6222 10219 6326 10276
rect 6222 10173 6251 10219
rect 6297 10173 6326 10219
rect 6222 10116 6326 10173
rect 6222 10070 6251 10116
rect 6297 10070 6326 10116
rect 6222 10013 6326 10070
rect 6222 9967 6251 10013
rect 6297 9967 6326 10013
rect 6222 9954 6326 9967
rect 6446 11757 6550 11770
rect 6446 10997 6475 11757
rect 6521 10997 6550 11757
rect 6446 10940 6550 10997
rect 6446 10894 6475 10940
rect 6521 10894 6550 10940
rect 6446 10837 6550 10894
rect 6446 10791 6475 10837
rect 6521 10791 6550 10837
rect 6446 10734 6550 10791
rect 6446 10688 6475 10734
rect 6521 10688 6550 10734
rect 6446 10631 6550 10688
rect 6446 10585 6475 10631
rect 6521 10585 6550 10631
rect 6446 10528 6550 10585
rect 6446 10482 6475 10528
rect 6521 10482 6550 10528
rect 6446 10425 6550 10482
rect 6446 10379 6475 10425
rect 6521 10379 6550 10425
rect 6446 10322 6550 10379
rect 6446 10276 6475 10322
rect 6521 10276 6550 10322
rect 6446 10219 6550 10276
rect 6446 10173 6475 10219
rect 6521 10173 6550 10219
rect 6446 10116 6550 10173
rect 6446 10070 6475 10116
rect 6521 10070 6550 10116
rect 6446 10013 6550 10070
rect 6446 9967 6475 10013
rect 6521 9967 6550 10013
rect 6446 9954 6550 9967
rect 6670 11757 6758 11770
rect 6670 10997 6699 11757
rect 6745 10997 6758 11757
rect 6670 10940 6758 10997
rect 6670 10894 6699 10940
rect 6745 10894 6758 10940
rect 6670 10837 6758 10894
rect 6670 10791 6699 10837
rect 6745 10791 6758 10837
rect 6670 10734 6758 10791
rect 6670 10688 6699 10734
rect 6745 10688 6758 10734
rect 6670 10631 6758 10688
rect 6670 10585 6699 10631
rect 6745 10585 6758 10631
rect 6670 10528 6758 10585
rect 6670 10482 6699 10528
rect 6745 10482 6758 10528
rect 6670 10425 6758 10482
rect 6670 10379 6699 10425
rect 6745 10379 6758 10425
rect 6670 10322 6758 10379
rect 6670 10276 6699 10322
rect 6745 10276 6758 10322
rect 6670 10219 6758 10276
rect 6670 10173 6699 10219
rect 6745 10173 6758 10219
rect 6670 10116 6758 10173
rect 6670 10070 6699 10116
rect 6745 10070 6758 10116
rect 6670 10013 6758 10070
rect 6670 9967 6699 10013
rect 6745 9967 6758 10013
rect 6670 9954 6758 9967
rect 6910 11757 6998 11770
rect 6910 10997 6923 11757
rect 6969 10997 6998 11757
rect 6910 10940 6998 10997
rect 6910 10894 6923 10940
rect 6969 10894 6998 10940
rect 6910 10837 6998 10894
rect 6910 10791 6923 10837
rect 6969 10791 6998 10837
rect 6910 10734 6998 10791
rect 6910 10688 6923 10734
rect 6969 10688 6998 10734
rect 6910 10631 6998 10688
rect 6910 10585 6923 10631
rect 6969 10585 6998 10631
rect 6910 10528 6998 10585
rect 6910 10482 6923 10528
rect 6969 10482 6998 10528
rect 6910 10425 6998 10482
rect 6910 10379 6923 10425
rect 6969 10379 6998 10425
rect 6910 10322 6998 10379
rect 6910 10276 6923 10322
rect 6969 10276 6998 10322
rect 6910 10219 6998 10276
rect 6910 10173 6923 10219
rect 6969 10173 6998 10219
rect 6910 10116 6998 10173
rect 6910 10070 6923 10116
rect 6969 10070 6998 10116
rect 6910 10013 6998 10070
rect 6910 9967 6923 10013
rect 6969 9967 6998 10013
rect 6910 9954 6998 9967
rect 7118 11757 7222 11770
rect 7118 10997 7147 11757
rect 7193 10997 7222 11757
rect 7118 10940 7222 10997
rect 7118 10894 7147 10940
rect 7193 10894 7222 10940
rect 7118 10837 7222 10894
rect 7118 10791 7147 10837
rect 7193 10791 7222 10837
rect 7118 10734 7222 10791
rect 7118 10688 7147 10734
rect 7193 10688 7222 10734
rect 7118 10631 7222 10688
rect 7118 10585 7147 10631
rect 7193 10585 7222 10631
rect 7118 10528 7222 10585
rect 7118 10482 7147 10528
rect 7193 10482 7222 10528
rect 7118 10425 7222 10482
rect 7118 10379 7147 10425
rect 7193 10379 7222 10425
rect 7118 10322 7222 10379
rect 7118 10276 7147 10322
rect 7193 10276 7222 10322
rect 7118 10219 7222 10276
rect 7118 10173 7147 10219
rect 7193 10173 7222 10219
rect 7118 10116 7222 10173
rect 7118 10070 7147 10116
rect 7193 10070 7222 10116
rect 7118 10013 7222 10070
rect 7118 9967 7147 10013
rect 7193 9967 7222 10013
rect 7118 9954 7222 9967
rect 7342 11757 7446 11770
rect 7342 10997 7371 11757
rect 7417 10997 7446 11757
rect 7342 10940 7446 10997
rect 7342 10894 7371 10940
rect 7417 10894 7446 10940
rect 7342 10837 7446 10894
rect 7342 10791 7371 10837
rect 7417 10791 7446 10837
rect 7342 10734 7446 10791
rect 7342 10688 7371 10734
rect 7417 10688 7446 10734
rect 7342 10631 7446 10688
rect 7342 10585 7371 10631
rect 7417 10585 7446 10631
rect 7342 10528 7446 10585
rect 7342 10482 7371 10528
rect 7417 10482 7446 10528
rect 7342 10425 7446 10482
rect 7342 10379 7371 10425
rect 7417 10379 7446 10425
rect 7342 10322 7446 10379
rect 7342 10276 7371 10322
rect 7417 10276 7446 10322
rect 7342 10219 7446 10276
rect 7342 10173 7371 10219
rect 7417 10173 7446 10219
rect 7342 10116 7446 10173
rect 7342 10070 7371 10116
rect 7417 10070 7446 10116
rect 7342 10013 7446 10070
rect 7342 9967 7371 10013
rect 7417 9967 7446 10013
rect 7342 9954 7446 9967
rect 7566 11757 7670 11770
rect 7566 10997 7595 11757
rect 7641 10997 7670 11757
rect 7566 10940 7670 10997
rect 7566 10894 7595 10940
rect 7641 10894 7670 10940
rect 7566 10837 7670 10894
rect 7566 10791 7595 10837
rect 7641 10791 7670 10837
rect 7566 10734 7670 10791
rect 7566 10688 7595 10734
rect 7641 10688 7670 10734
rect 7566 10631 7670 10688
rect 7566 10585 7595 10631
rect 7641 10585 7670 10631
rect 7566 10528 7670 10585
rect 7566 10482 7595 10528
rect 7641 10482 7670 10528
rect 7566 10425 7670 10482
rect 7566 10379 7595 10425
rect 7641 10379 7670 10425
rect 7566 10322 7670 10379
rect 7566 10276 7595 10322
rect 7641 10276 7670 10322
rect 7566 10219 7670 10276
rect 7566 10173 7595 10219
rect 7641 10173 7670 10219
rect 7566 10116 7670 10173
rect 7566 10070 7595 10116
rect 7641 10070 7670 10116
rect 7566 10013 7670 10070
rect 7566 9967 7595 10013
rect 7641 9967 7670 10013
rect 7566 9954 7670 9967
rect 7790 11757 7878 11770
rect 7790 10997 7819 11757
rect 7865 10997 7878 11757
rect 7790 10940 7878 10997
rect 7790 10894 7819 10940
rect 7865 10894 7878 10940
rect 7790 10837 7878 10894
rect 7790 10791 7819 10837
rect 7865 10791 7878 10837
rect 7790 10734 7878 10791
rect 7790 10688 7819 10734
rect 7865 10688 7878 10734
rect 7790 10631 7878 10688
rect 7790 10585 7819 10631
rect 7865 10585 7878 10631
rect 7790 10528 7878 10585
rect 7790 10482 7819 10528
rect 7865 10482 7878 10528
rect 7790 10425 7878 10482
rect 7790 10379 7819 10425
rect 7865 10379 7878 10425
rect 7790 10322 7878 10379
rect 7790 10276 7819 10322
rect 7865 10276 7878 10322
rect 7790 10219 7878 10276
rect 7790 10173 7819 10219
rect 7865 10173 7878 10219
rect 7790 10116 7878 10173
rect 7790 10070 7819 10116
rect 7865 10070 7878 10116
rect 7790 10013 7878 10070
rect 7790 9967 7819 10013
rect 7865 9967 7878 10013
rect 7790 9954 7878 9967
rect 8030 11757 8118 11770
rect 8030 10997 8043 11757
rect 8089 10997 8118 11757
rect 8030 10940 8118 10997
rect 8030 10894 8043 10940
rect 8089 10894 8118 10940
rect 8030 10837 8118 10894
rect 8030 10791 8043 10837
rect 8089 10791 8118 10837
rect 8030 10734 8118 10791
rect 8030 10688 8043 10734
rect 8089 10688 8118 10734
rect 8030 10631 8118 10688
rect 8030 10585 8043 10631
rect 8089 10585 8118 10631
rect 8030 10528 8118 10585
rect 8030 10482 8043 10528
rect 8089 10482 8118 10528
rect 8030 10425 8118 10482
rect 8030 10379 8043 10425
rect 8089 10379 8118 10425
rect 8030 10322 8118 10379
rect 8030 10276 8043 10322
rect 8089 10276 8118 10322
rect 8030 10219 8118 10276
rect 8030 10173 8043 10219
rect 8089 10173 8118 10219
rect 8030 10116 8118 10173
rect 8030 10070 8043 10116
rect 8089 10070 8118 10116
rect 8030 10013 8118 10070
rect 8030 9967 8043 10013
rect 8089 9967 8118 10013
rect 8030 9954 8118 9967
rect 8238 11757 8342 11770
rect 8238 10997 8267 11757
rect 8313 10997 8342 11757
rect 8238 10940 8342 10997
rect 8238 10894 8267 10940
rect 8313 10894 8342 10940
rect 8238 10837 8342 10894
rect 8238 10791 8267 10837
rect 8313 10791 8342 10837
rect 8238 10734 8342 10791
rect 8238 10688 8267 10734
rect 8313 10688 8342 10734
rect 8238 10631 8342 10688
rect 8238 10585 8267 10631
rect 8313 10585 8342 10631
rect 8238 10528 8342 10585
rect 8238 10482 8267 10528
rect 8313 10482 8342 10528
rect 8238 10425 8342 10482
rect 8238 10379 8267 10425
rect 8313 10379 8342 10425
rect 8238 10322 8342 10379
rect 8238 10276 8267 10322
rect 8313 10276 8342 10322
rect 8238 10219 8342 10276
rect 8238 10173 8267 10219
rect 8313 10173 8342 10219
rect 8238 10116 8342 10173
rect 8238 10070 8267 10116
rect 8313 10070 8342 10116
rect 8238 10013 8342 10070
rect 8238 9967 8267 10013
rect 8313 9967 8342 10013
rect 8238 9954 8342 9967
rect 8462 11757 8566 11770
rect 8462 10997 8491 11757
rect 8537 10997 8566 11757
rect 8462 10940 8566 10997
rect 8462 10894 8491 10940
rect 8537 10894 8566 10940
rect 8462 10837 8566 10894
rect 8462 10791 8491 10837
rect 8537 10791 8566 10837
rect 8462 10734 8566 10791
rect 8462 10688 8491 10734
rect 8537 10688 8566 10734
rect 8462 10631 8566 10688
rect 8462 10585 8491 10631
rect 8537 10585 8566 10631
rect 8462 10528 8566 10585
rect 8462 10482 8491 10528
rect 8537 10482 8566 10528
rect 8462 10425 8566 10482
rect 8462 10379 8491 10425
rect 8537 10379 8566 10425
rect 8462 10322 8566 10379
rect 8462 10276 8491 10322
rect 8537 10276 8566 10322
rect 8462 10219 8566 10276
rect 8462 10173 8491 10219
rect 8537 10173 8566 10219
rect 8462 10116 8566 10173
rect 8462 10070 8491 10116
rect 8537 10070 8566 10116
rect 8462 10013 8566 10070
rect 8462 9967 8491 10013
rect 8537 9967 8566 10013
rect 8462 9954 8566 9967
rect 8686 11757 8790 11770
rect 8686 10997 8715 11757
rect 8761 10997 8790 11757
rect 8686 10940 8790 10997
rect 8686 10894 8715 10940
rect 8761 10894 8790 10940
rect 8686 10837 8790 10894
rect 8686 10791 8715 10837
rect 8761 10791 8790 10837
rect 8686 10734 8790 10791
rect 8686 10688 8715 10734
rect 8761 10688 8790 10734
rect 8686 10631 8790 10688
rect 8686 10585 8715 10631
rect 8761 10585 8790 10631
rect 8686 10528 8790 10585
rect 8686 10482 8715 10528
rect 8761 10482 8790 10528
rect 8686 10425 8790 10482
rect 8686 10379 8715 10425
rect 8761 10379 8790 10425
rect 8686 10322 8790 10379
rect 8686 10276 8715 10322
rect 8761 10276 8790 10322
rect 8686 10219 8790 10276
rect 8686 10173 8715 10219
rect 8761 10173 8790 10219
rect 8686 10116 8790 10173
rect 8686 10070 8715 10116
rect 8761 10070 8790 10116
rect 8686 10013 8790 10070
rect 8686 9967 8715 10013
rect 8761 9967 8790 10013
rect 8686 9954 8790 9967
rect 8910 11757 8998 11770
rect 8910 10997 8939 11757
rect 8985 10997 8998 11757
rect 8910 10940 8998 10997
rect 8910 10894 8939 10940
rect 8985 10894 8998 10940
rect 8910 10837 8998 10894
rect 8910 10791 8939 10837
rect 8985 10791 8998 10837
rect 8910 10734 8998 10791
rect 8910 10688 8939 10734
rect 8985 10688 8998 10734
rect 8910 10631 8998 10688
rect 8910 10585 8939 10631
rect 8985 10585 8998 10631
rect 8910 10528 8998 10585
rect 8910 10482 8939 10528
rect 8985 10482 8998 10528
rect 8910 10425 8998 10482
rect 8910 10379 8939 10425
rect 8985 10379 8998 10425
rect 8910 10322 8998 10379
rect 8910 10276 8939 10322
rect 8985 10276 8998 10322
rect 8910 10219 8998 10276
rect 8910 10173 8939 10219
rect 8985 10173 8998 10219
rect 8910 10116 8998 10173
rect 8910 10070 8939 10116
rect 8985 10070 8998 10116
rect 8910 10013 8998 10070
rect 8910 9967 8939 10013
rect 8985 9967 8998 10013
rect 8910 9954 8998 9967
rect 9150 11757 9238 11770
rect 9150 10997 9163 11757
rect 9209 10997 9238 11757
rect 9150 10940 9238 10997
rect 9150 10894 9163 10940
rect 9209 10894 9238 10940
rect 9150 10837 9238 10894
rect 9150 10791 9163 10837
rect 9209 10791 9238 10837
rect 9150 10734 9238 10791
rect 9150 10688 9163 10734
rect 9209 10688 9238 10734
rect 9150 10631 9238 10688
rect 9150 10585 9163 10631
rect 9209 10585 9238 10631
rect 9150 10528 9238 10585
rect 9150 10482 9163 10528
rect 9209 10482 9238 10528
rect 9150 10425 9238 10482
rect 9150 10379 9163 10425
rect 9209 10379 9238 10425
rect 9150 10322 9238 10379
rect 9150 10276 9163 10322
rect 9209 10276 9238 10322
rect 9150 10219 9238 10276
rect 9150 10173 9163 10219
rect 9209 10173 9238 10219
rect 9150 10116 9238 10173
rect 9150 10070 9163 10116
rect 9209 10070 9238 10116
rect 9150 10013 9238 10070
rect 9150 9967 9163 10013
rect 9209 9967 9238 10013
rect 9150 9954 9238 9967
rect 9358 11757 9462 11770
rect 9358 10997 9387 11757
rect 9433 10997 9462 11757
rect 9358 10940 9462 10997
rect 9358 10894 9387 10940
rect 9433 10894 9462 10940
rect 9358 10837 9462 10894
rect 9358 10791 9387 10837
rect 9433 10791 9462 10837
rect 9358 10734 9462 10791
rect 9358 10688 9387 10734
rect 9433 10688 9462 10734
rect 9358 10631 9462 10688
rect 9358 10585 9387 10631
rect 9433 10585 9462 10631
rect 9358 10528 9462 10585
rect 9358 10482 9387 10528
rect 9433 10482 9462 10528
rect 9358 10425 9462 10482
rect 9358 10379 9387 10425
rect 9433 10379 9462 10425
rect 9358 10322 9462 10379
rect 9358 10276 9387 10322
rect 9433 10276 9462 10322
rect 9358 10219 9462 10276
rect 9358 10173 9387 10219
rect 9433 10173 9462 10219
rect 9358 10116 9462 10173
rect 9358 10070 9387 10116
rect 9433 10070 9462 10116
rect 9358 10013 9462 10070
rect 9358 9967 9387 10013
rect 9433 9967 9462 10013
rect 9358 9954 9462 9967
rect 9582 11757 9686 11770
rect 9582 10997 9611 11757
rect 9657 10997 9686 11757
rect 9582 10940 9686 10997
rect 9582 10894 9611 10940
rect 9657 10894 9686 10940
rect 9582 10837 9686 10894
rect 9582 10791 9611 10837
rect 9657 10791 9686 10837
rect 9582 10734 9686 10791
rect 9582 10688 9611 10734
rect 9657 10688 9686 10734
rect 9582 10631 9686 10688
rect 9582 10585 9611 10631
rect 9657 10585 9686 10631
rect 9582 10528 9686 10585
rect 9582 10482 9611 10528
rect 9657 10482 9686 10528
rect 9582 10425 9686 10482
rect 9582 10379 9611 10425
rect 9657 10379 9686 10425
rect 9582 10322 9686 10379
rect 9582 10276 9611 10322
rect 9657 10276 9686 10322
rect 9582 10219 9686 10276
rect 9582 10173 9611 10219
rect 9657 10173 9686 10219
rect 9582 10116 9686 10173
rect 9582 10070 9611 10116
rect 9657 10070 9686 10116
rect 9582 10013 9686 10070
rect 9582 9967 9611 10013
rect 9657 9967 9686 10013
rect 9582 9954 9686 9967
rect 9806 11757 9910 11770
rect 9806 10997 9835 11757
rect 9881 10997 9910 11757
rect 9806 10940 9910 10997
rect 9806 10894 9835 10940
rect 9881 10894 9910 10940
rect 9806 10837 9910 10894
rect 9806 10791 9835 10837
rect 9881 10791 9910 10837
rect 9806 10734 9910 10791
rect 9806 10688 9835 10734
rect 9881 10688 9910 10734
rect 9806 10631 9910 10688
rect 9806 10585 9835 10631
rect 9881 10585 9910 10631
rect 9806 10528 9910 10585
rect 9806 10482 9835 10528
rect 9881 10482 9910 10528
rect 9806 10425 9910 10482
rect 9806 10379 9835 10425
rect 9881 10379 9910 10425
rect 9806 10322 9910 10379
rect 9806 10276 9835 10322
rect 9881 10276 9910 10322
rect 9806 10219 9910 10276
rect 9806 10173 9835 10219
rect 9881 10173 9910 10219
rect 9806 10116 9910 10173
rect 9806 10070 9835 10116
rect 9881 10070 9910 10116
rect 9806 10013 9910 10070
rect 9806 9967 9835 10013
rect 9881 9967 9910 10013
rect 9806 9954 9910 9967
rect 10030 11757 10118 11770
rect 10030 10997 10059 11757
rect 10105 10997 10118 11757
rect 10030 10940 10118 10997
rect 10030 10894 10059 10940
rect 10105 10894 10118 10940
rect 10030 10837 10118 10894
rect 10030 10791 10059 10837
rect 10105 10791 10118 10837
rect 10030 10734 10118 10791
rect 10030 10688 10059 10734
rect 10105 10688 10118 10734
rect 10030 10631 10118 10688
rect 10030 10585 10059 10631
rect 10105 10585 10118 10631
rect 10030 10528 10118 10585
rect 10030 10482 10059 10528
rect 10105 10482 10118 10528
rect 10030 10425 10118 10482
rect 10030 10379 10059 10425
rect 10105 10379 10118 10425
rect 10030 10322 10118 10379
rect 10030 10276 10059 10322
rect 10105 10276 10118 10322
rect 10030 10219 10118 10276
rect 10030 10173 10059 10219
rect 10105 10173 10118 10219
rect 10030 10116 10118 10173
rect 10030 10070 10059 10116
rect 10105 10070 10118 10116
rect 10030 10013 10118 10070
rect 10030 9967 10059 10013
rect 10105 9967 10118 10013
rect 10030 9954 10118 9967
rect 10270 11757 10358 11770
rect 10270 10997 10283 11757
rect 10329 10997 10358 11757
rect 10270 10940 10358 10997
rect 10270 10894 10283 10940
rect 10329 10894 10358 10940
rect 10270 10837 10358 10894
rect 10270 10791 10283 10837
rect 10329 10791 10358 10837
rect 10270 10734 10358 10791
rect 10270 10688 10283 10734
rect 10329 10688 10358 10734
rect 10270 10631 10358 10688
rect 10270 10585 10283 10631
rect 10329 10585 10358 10631
rect 10270 10528 10358 10585
rect 10270 10482 10283 10528
rect 10329 10482 10358 10528
rect 10270 10425 10358 10482
rect 10270 10379 10283 10425
rect 10329 10379 10358 10425
rect 10270 10322 10358 10379
rect 10270 10276 10283 10322
rect 10329 10276 10358 10322
rect 10270 10219 10358 10276
rect 10270 10173 10283 10219
rect 10329 10173 10358 10219
rect 10270 10116 10358 10173
rect 10270 10070 10283 10116
rect 10329 10070 10358 10116
rect 10270 10013 10358 10070
rect 10270 9967 10283 10013
rect 10329 9967 10358 10013
rect 10270 9954 10358 9967
rect 10478 11757 10582 11770
rect 10478 10997 10507 11757
rect 10553 10997 10582 11757
rect 10478 10940 10582 10997
rect 10478 10894 10507 10940
rect 10553 10894 10582 10940
rect 10478 10837 10582 10894
rect 10478 10791 10507 10837
rect 10553 10791 10582 10837
rect 10478 10734 10582 10791
rect 10478 10688 10507 10734
rect 10553 10688 10582 10734
rect 10478 10631 10582 10688
rect 10478 10585 10507 10631
rect 10553 10585 10582 10631
rect 10478 10528 10582 10585
rect 10478 10482 10507 10528
rect 10553 10482 10582 10528
rect 10478 10425 10582 10482
rect 10478 10379 10507 10425
rect 10553 10379 10582 10425
rect 10478 10322 10582 10379
rect 10478 10276 10507 10322
rect 10553 10276 10582 10322
rect 10478 10219 10582 10276
rect 10478 10173 10507 10219
rect 10553 10173 10582 10219
rect 10478 10116 10582 10173
rect 10478 10070 10507 10116
rect 10553 10070 10582 10116
rect 10478 10013 10582 10070
rect 10478 9967 10507 10013
rect 10553 9967 10582 10013
rect 10478 9954 10582 9967
rect 10702 11757 10806 11770
rect 10702 10997 10731 11757
rect 10777 10997 10806 11757
rect 10702 10940 10806 10997
rect 10702 10894 10731 10940
rect 10777 10894 10806 10940
rect 10702 10837 10806 10894
rect 10702 10791 10731 10837
rect 10777 10791 10806 10837
rect 10702 10734 10806 10791
rect 10702 10688 10731 10734
rect 10777 10688 10806 10734
rect 10702 10631 10806 10688
rect 10702 10585 10731 10631
rect 10777 10585 10806 10631
rect 10702 10528 10806 10585
rect 10702 10482 10731 10528
rect 10777 10482 10806 10528
rect 10702 10425 10806 10482
rect 10702 10379 10731 10425
rect 10777 10379 10806 10425
rect 10702 10322 10806 10379
rect 10702 10276 10731 10322
rect 10777 10276 10806 10322
rect 10702 10219 10806 10276
rect 10702 10173 10731 10219
rect 10777 10173 10806 10219
rect 10702 10116 10806 10173
rect 10702 10070 10731 10116
rect 10777 10070 10806 10116
rect 10702 10013 10806 10070
rect 10702 9967 10731 10013
rect 10777 9967 10806 10013
rect 10702 9954 10806 9967
rect 10926 11757 11030 11770
rect 10926 10997 10955 11757
rect 11001 10997 11030 11757
rect 10926 10940 11030 10997
rect 10926 10894 10955 10940
rect 11001 10894 11030 10940
rect 10926 10837 11030 10894
rect 10926 10791 10955 10837
rect 11001 10791 11030 10837
rect 10926 10734 11030 10791
rect 10926 10688 10955 10734
rect 11001 10688 11030 10734
rect 10926 10631 11030 10688
rect 10926 10585 10955 10631
rect 11001 10585 11030 10631
rect 10926 10528 11030 10585
rect 10926 10482 10955 10528
rect 11001 10482 11030 10528
rect 10926 10425 11030 10482
rect 10926 10379 10955 10425
rect 11001 10379 11030 10425
rect 10926 10322 11030 10379
rect 10926 10276 10955 10322
rect 11001 10276 11030 10322
rect 10926 10219 11030 10276
rect 10926 10173 10955 10219
rect 11001 10173 11030 10219
rect 10926 10116 11030 10173
rect 10926 10070 10955 10116
rect 11001 10070 11030 10116
rect 10926 10013 11030 10070
rect 10926 9967 10955 10013
rect 11001 9967 11030 10013
rect 10926 9954 11030 9967
rect 11150 11757 11238 11770
rect 11150 10997 11179 11757
rect 11225 10997 11238 11757
rect 11150 10940 11238 10997
rect 11150 10894 11179 10940
rect 11225 10894 11238 10940
rect 11150 10837 11238 10894
rect 11150 10791 11179 10837
rect 11225 10791 11238 10837
rect 11150 10734 11238 10791
rect 11150 10688 11179 10734
rect 11225 10688 11238 10734
rect 11150 10631 11238 10688
rect 11150 10585 11179 10631
rect 11225 10585 11238 10631
rect 11150 10528 11238 10585
rect 11150 10482 11179 10528
rect 11225 10482 11238 10528
rect 11150 10425 11238 10482
rect 11150 10379 11179 10425
rect 11225 10379 11238 10425
rect 11150 10322 11238 10379
rect 11150 10276 11179 10322
rect 11225 10276 11238 10322
rect 11150 10219 11238 10276
rect 11150 10173 11179 10219
rect 11225 10173 11238 10219
rect 11150 10116 11238 10173
rect 11150 10070 11179 10116
rect 11225 10070 11238 10116
rect 11150 10013 11238 10070
rect 11150 9967 11179 10013
rect 11225 9967 11238 10013
rect 11150 9954 11238 9967
rect 11390 11757 11478 11770
rect 11390 10997 11403 11757
rect 11449 10997 11478 11757
rect 11390 10940 11478 10997
rect 11390 10894 11403 10940
rect 11449 10894 11478 10940
rect 11390 10837 11478 10894
rect 11390 10791 11403 10837
rect 11449 10791 11478 10837
rect 11390 10734 11478 10791
rect 11390 10688 11403 10734
rect 11449 10688 11478 10734
rect 11390 10631 11478 10688
rect 11390 10585 11403 10631
rect 11449 10585 11478 10631
rect 11390 10528 11478 10585
rect 11390 10482 11403 10528
rect 11449 10482 11478 10528
rect 11390 10425 11478 10482
rect 11390 10379 11403 10425
rect 11449 10379 11478 10425
rect 11390 10322 11478 10379
rect 11390 10276 11403 10322
rect 11449 10276 11478 10322
rect 11390 10219 11478 10276
rect 11390 10173 11403 10219
rect 11449 10173 11478 10219
rect 11390 10116 11478 10173
rect 11390 10070 11403 10116
rect 11449 10070 11478 10116
rect 11390 10013 11478 10070
rect 11390 9967 11403 10013
rect 11449 9967 11478 10013
rect 11390 9954 11478 9967
rect 11598 11757 11702 11770
rect 11598 10997 11627 11757
rect 11673 10997 11702 11757
rect 11598 10940 11702 10997
rect 11598 10894 11627 10940
rect 11673 10894 11702 10940
rect 11598 10837 11702 10894
rect 11598 10791 11627 10837
rect 11673 10791 11702 10837
rect 11598 10734 11702 10791
rect 11598 10688 11627 10734
rect 11673 10688 11702 10734
rect 11598 10631 11702 10688
rect 11598 10585 11627 10631
rect 11673 10585 11702 10631
rect 11598 10528 11702 10585
rect 11598 10482 11627 10528
rect 11673 10482 11702 10528
rect 11598 10425 11702 10482
rect 11598 10379 11627 10425
rect 11673 10379 11702 10425
rect 11598 10322 11702 10379
rect 11598 10276 11627 10322
rect 11673 10276 11702 10322
rect 11598 10219 11702 10276
rect 11598 10173 11627 10219
rect 11673 10173 11702 10219
rect 11598 10116 11702 10173
rect 11598 10070 11627 10116
rect 11673 10070 11702 10116
rect 11598 10013 11702 10070
rect 11598 9967 11627 10013
rect 11673 9967 11702 10013
rect 11598 9954 11702 9967
rect 11822 11757 11926 11770
rect 11822 10997 11851 11757
rect 11897 10997 11926 11757
rect 11822 10940 11926 10997
rect 11822 10894 11851 10940
rect 11897 10894 11926 10940
rect 11822 10837 11926 10894
rect 11822 10791 11851 10837
rect 11897 10791 11926 10837
rect 11822 10734 11926 10791
rect 11822 10688 11851 10734
rect 11897 10688 11926 10734
rect 11822 10631 11926 10688
rect 11822 10585 11851 10631
rect 11897 10585 11926 10631
rect 11822 10528 11926 10585
rect 11822 10482 11851 10528
rect 11897 10482 11926 10528
rect 11822 10425 11926 10482
rect 11822 10379 11851 10425
rect 11897 10379 11926 10425
rect 11822 10322 11926 10379
rect 11822 10276 11851 10322
rect 11897 10276 11926 10322
rect 11822 10219 11926 10276
rect 11822 10173 11851 10219
rect 11897 10173 11926 10219
rect 11822 10116 11926 10173
rect 11822 10070 11851 10116
rect 11897 10070 11926 10116
rect 11822 10013 11926 10070
rect 11822 9967 11851 10013
rect 11897 9967 11926 10013
rect 11822 9954 11926 9967
rect 12046 11757 12150 11770
rect 12046 10997 12075 11757
rect 12121 10997 12150 11757
rect 12046 10940 12150 10997
rect 12046 10894 12075 10940
rect 12121 10894 12150 10940
rect 12046 10837 12150 10894
rect 12046 10791 12075 10837
rect 12121 10791 12150 10837
rect 12046 10734 12150 10791
rect 12046 10688 12075 10734
rect 12121 10688 12150 10734
rect 12046 10631 12150 10688
rect 12046 10585 12075 10631
rect 12121 10585 12150 10631
rect 12046 10528 12150 10585
rect 12046 10482 12075 10528
rect 12121 10482 12150 10528
rect 12046 10425 12150 10482
rect 12046 10379 12075 10425
rect 12121 10379 12150 10425
rect 12046 10322 12150 10379
rect 12046 10276 12075 10322
rect 12121 10276 12150 10322
rect 12046 10219 12150 10276
rect 12046 10173 12075 10219
rect 12121 10173 12150 10219
rect 12046 10116 12150 10173
rect 12046 10070 12075 10116
rect 12121 10070 12150 10116
rect 12046 10013 12150 10070
rect 12046 9967 12075 10013
rect 12121 9967 12150 10013
rect 12046 9954 12150 9967
rect 12270 11757 12358 11770
rect 12270 10997 12299 11757
rect 12345 10997 12358 11757
rect 12270 10940 12358 10997
rect 12270 10894 12299 10940
rect 12345 10894 12358 10940
rect 12270 10837 12358 10894
rect 12270 10791 12299 10837
rect 12345 10791 12358 10837
rect 12270 10734 12358 10791
rect 12270 10688 12299 10734
rect 12345 10688 12358 10734
rect 12270 10631 12358 10688
rect 12270 10585 12299 10631
rect 12345 10585 12358 10631
rect 12270 10528 12358 10585
rect 12270 10482 12299 10528
rect 12345 10482 12358 10528
rect 12270 10425 12358 10482
rect 12270 10379 12299 10425
rect 12345 10379 12358 10425
rect 12270 10322 12358 10379
rect 12270 10276 12299 10322
rect 12345 10276 12358 10322
rect 12270 10219 12358 10276
rect 12270 10173 12299 10219
rect 12345 10173 12358 10219
rect 12270 10116 12358 10173
rect 12270 10070 12299 10116
rect 12345 10070 12358 10116
rect 12270 10013 12358 10070
rect 12270 9967 12299 10013
rect 12345 9967 12358 10013
rect 12270 9954 12358 9967
rect 12510 11757 12598 11770
rect 12510 10997 12523 11757
rect 12569 10997 12598 11757
rect 12510 10940 12598 10997
rect 12510 10894 12523 10940
rect 12569 10894 12598 10940
rect 12510 10837 12598 10894
rect 12510 10791 12523 10837
rect 12569 10791 12598 10837
rect 12510 10734 12598 10791
rect 12510 10688 12523 10734
rect 12569 10688 12598 10734
rect 12510 10631 12598 10688
rect 12510 10585 12523 10631
rect 12569 10585 12598 10631
rect 12510 10528 12598 10585
rect 12510 10482 12523 10528
rect 12569 10482 12598 10528
rect 12510 10425 12598 10482
rect 12510 10379 12523 10425
rect 12569 10379 12598 10425
rect 12510 10322 12598 10379
rect 12510 10276 12523 10322
rect 12569 10276 12598 10322
rect 12510 10219 12598 10276
rect 12510 10173 12523 10219
rect 12569 10173 12598 10219
rect 12510 10116 12598 10173
rect 12510 10070 12523 10116
rect 12569 10070 12598 10116
rect 12510 10013 12598 10070
rect 12510 9967 12523 10013
rect 12569 9967 12598 10013
rect 12510 9954 12598 9967
rect 12718 11757 12822 11770
rect 12718 10997 12747 11757
rect 12793 10997 12822 11757
rect 12718 10940 12822 10997
rect 12718 10894 12747 10940
rect 12793 10894 12822 10940
rect 12718 10837 12822 10894
rect 12718 10791 12747 10837
rect 12793 10791 12822 10837
rect 12718 10734 12822 10791
rect 12718 10688 12747 10734
rect 12793 10688 12822 10734
rect 12718 10631 12822 10688
rect 12718 10585 12747 10631
rect 12793 10585 12822 10631
rect 12718 10528 12822 10585
rect 12718 10482 12747 10528
rect 12793 10482 12822 10528
rect 12718 10425 12822 10482
rect 12718 10379 12747 10425
rect 12793 10379 12822 10425
rect 12718 10322 12822 10379
rect 12718 10276 12747 10322
rect 12793 10276 12822 10322
rect 12718 10219 12822 10276
rect 12718 10173 12747 10219
rect 12793 10173 12822 10219
rect 12718 10116 12822 10173
rect 12718 10070 12747 10116
rect 12793 10070 12822 10116
rect 12718 10013 12822 10070
rect 12718 9967 12747 10013
rect 12793 9967 12822 10013
rect 12718 9954 12822 9967
rect 12942 11757 13046 11770
rect 12942 10997 12971 11757
rect 13017 10997 13046 11757
rect 12942 10940 13046 10997
rect 12942 10894 12971 10940
rect 13017 10894 13046 10940
rect 12942 10837 13046 10894
rect 12942 10791 12971 10837
rect 13017 10791 13046 10837
rect 12942 10734 13046 10791
rect 12942 10688 12971 10734
rect 13017 10688 13046 10734
rect 12942 10631 13046 10688
rect 12942 10585 12971 10631
rect 13017 10585 13046 10631
rect 12942 10528 13046 10585
rect 12942 10482 12971 10528
rect 13017 10482 13046 10528
rect 12942 10425 13046 10482
rect 12942 10379 12971 10425
rect 13017 10379 13046 10425
rect 12942 10322 13046 10379
rect 12942 10276 12971 10322
rect 13017 10276 13046 10322
rect 12942 10219 13046 10276
rect 12942 10173 12971 10219
rect 13017 10173 13046 10219
rect 12942 10116 13046 10173
rect 12942 10070 12971 10116
rect 13017 10070 13046 10116
rect 12942 10013 13046 10070
rect 12942 9967 12971 10013
rect 13017 9967 13046 10013
rect 12942 9954 13046 9967
rect 13166 11757 13270 11770
rect 13166 10997 13195 11757
rect 13241 10997 13270 11757
rect 13166 10940 13270 10997
rect 13166 10894 13195 10940
rect 13241 10894 13270 10940
rect 13166 10837 13270 10894
rect 13166 10791 13195 10837
rect 13241 10791 13270 10837
rect 13166 10734 13270 10791
rect 13166 10688 13195 10734
rect 13241 10688 13270 10734
rect 13166 10631 13270 10688
rect 13166 10585 13195 10631
rect 13241 10585 13270 10631
rect 13166 10528 13270 10585
rect 13166 10482 13195 10528
rect 13241 10482 13270 10528
rect 13166 10425 13270 10482
rect 13166 10379 13195 10425
rect 13241 10379 13270 10425
rect 13166 10322 13270 10379
rect 13166 10276 13195 10322
rect 13241 10276 13270 10322
rect 13166 10219 13270 10276
rect 13166 10173 13195 10219
rect 13241 10173 13270 10219
rect 13166 10116 13270 10173
rect 13166 10070 13195 10116
rect 13241 10070 13270 10116
rect 13166 10013 13270 10070
rect 13166 9967 13195 10013
rect 13241 9967 13270 10013
rect 13166 9954 13270 9967
rect 13390 11757 13478 11770
rect 13390 10997 13419 11757
rect 13465 10997 13478 11757
rect 13390 10940 13478 10997
rect 13390 10894 13419 10940
rect 13465 10894 13478 10940
rect 13390 10837 13478 10894
rect 13390 10791 13419 10837
rect 13465 10791 13478 10837
rect 13390 10734 13478 10791
rect 13390 10688 13419 10734
rect 13465 10688 13478 10734
rect 13390 10631 13478 10688
rect 13390 10585 13419 10631
rect 13465 10585 13478 10631
rect 13390 10528 13478 10585
rect 13390 10482 13419 10528
rect 13465 10482 13478 10528
rect 13390 10425 13478 10482
rect 13390 10379 13419 10425
rect 13465 10379 13478 10425
rect 13390 10322 13478 10379
rect 13390 10276 13419 10322
rect 13465 10276 13478 10322
rect 13390 10219 13478 10276
rect 13390 10173 13419 10219
rect 13465 10173 13478 10219
rect 13390 10116 13478 10173
rect 13390 10070 13419 10116
rect 13465 10070 13478 10116
rect 13390 10013 13478 10070
rect 13390 9967 13419 10013
rect 13465 9967 13478 10013
rect 13390 9954 13478 9967
rect 13630 11757 13718 11770
rect 13630 10997 13643 11757
rect 13689 10997 13718 11757
rect 13630 10940 13718 10997
rect 13630 10894 13643 10940
rect 13689 10894 13718 10940
rect 13630 10837 13718 10894
rect 13630 10791 13643 10837
rect 13689 10791 13718 10837
rect 13630 10734 13718 10791
rect 13630 10688 13643 10734
rect 13689 10688 13718 10734
rect 13630 10631 13718 10688
rect 13630 10585 13643 10631
rect 13689 10585 13718 10631
rect 13630 10528 13718 10585
rect 13630 10482 13643 10528
rect 13689 10482 13718 10528
rect 13630 10425 13718 10482
rect 13630 10379 13643 10425
rect 13689 10379 13718 10425
rect 13630 10322 13718 10379
rect 13630 10276 13643 10322
rect 13689 10276 13718 10322
rect 13630 10219 13718 10276
rect 13630 10173 13643 10219
rect 13689 10173 13718 10219
rect 13630 10116 13718 10173
rect 13630 10070 13643 10116
rect 13689 10070 13718 10116
rect 13630 10013 13718 10070
rect 13630 9967 13643 10013
rect 13689 9967 13718 10013
rect 13630 9954 13718 9967
rect 13838 11757 13942 11770
rect 13838 10997 13867 11757
rect 13913 10997 13942 11757
rect 13838 10940 13942 10997
rect 13838 10894 13867 10940
rect 13913 10894 13942 10940
rect 13838 10837 13942 10894
rect 13838 10791 13867 10837
rect 13913 10791 13942 10837
rect 13838 10734 13942 10791
rect 13838 10688 13867 10734
rect 13913 10688 13942 10734
rect 13838 10631 13942 10688
rect 13838 10585 13867 10631
rect 13913 10585 13942 10631
rect 13838 10528 13942 10585
rect 13838 10482 13867 10528
rect 13913 10482 13942 10528
rect 13838 10425 13942 10482
rect 13838 10379 13867 10425
rect 13913 10379 13942 10425
rect 13838 10322 13942 10379
rect 13838 10276 13867 10322
rect 13913 10276 13942 10322
rect 13838 10219 13942 10276
rect 13838 10173 13867 10219
rect 13913 10173 13942 10219
rect 13838 10116 13942 10173
rect 13838 10070 13867 10116
rect 13913 10070 13942 10116
rect 13838 10013 13942 10070
rect 13838 9967 13867 10013
rect 13913 9967 13942 10013
rect 13838 9954 13942 9967
rect 14062 11757 14166 11770
rect 14062 10997 14091 11757
rect 14137 10997 14166 11757
rect 14062 10940 14166 10997
rect 14062 10894 14091 10940
rect 14137 10894 14166 10940
rect 14062 10837 14166 10894
rect 14062 10791 14091 10837
rect 14137 10791 14166 10837
rect 14062 10734 14166 10791
rect 14062 10688 14091 10734
rect 14137 10688 14166 10734
rect 14062 10631 14166 10688
rect 14062 10585 14091 10631
rect 14137 10585 14166 10631
rect 14062 10528 14166 10585
rect 14062 10482 14091 10528
rect 14137 10482 14166 10528
rect 14062 10425 14166 10482
rect 14062 10379 14091 10425
rect 14137 10379 14166 10425
rect 14062 10322 14166 10379
rect 14062 10276 14091 10322
rect 14137 10276 14166 10322
rect 14062 10219 14166 10276
rect 14062 10173 14091 10219
rect 14137 10173 14166 10219
rect 14062 10116 14166 10173
rect 14062 10070 14091 10116
rect 14137 10070 14166 10116
rect 14062 10013 14166 10070
rect 14062 9967 14091 10013
rect 14137 9967 14166 10013
rect 14062 9954 14166 9967
rect 14286 11757 14390 11770
rect 14286 10997 14315 11757
rect 14361 10997 14390 11757
rect 14286 10940 14390 10997
rect 14286 10894 14315 10940
rect 14361 10894 14390 10940
rect 14286 10837 14390 10894
rect 14286 10791 14315 10837
rect 14361 10791 14390 10837
rect 14286 10734 14390 10791
rect 14286 10688 14315 10734
rect 14361 10688 14390 10734
rect 14286 10631 14390 10688
rect 14286 10585 14315 10631
rect 14361 10585 14390 10631
rect 14286 10528 14390 10585
rect 14286 10482 14315 10528
rect 14361 10482 14390 10528
rect 14286 10425 14390 10482
rect 14286 10379 14315 10425
rect 14361 10379 14390 10425
rect 14286 10322 14390 10379
rect 14286 10276 14315 10322
rect 14361 10276 14390 10322
rect 14286 10219 14390 10276
rect 14286 10173 14315 10219
rect 14361 10173 14390 10219
rect 14286 10116 14390 10173
rect 14286 10070 14315 10116
rect 14361 10070 14390 10116
rect 14286 10013 14390 10070
rect 14286 9967 14315 10013
rect 14361 9967 14390 10013
rect 14286 9954 14390 9967
rect 14510 11757 14598 11770
rect 14510 10997 14539 11757
rect 14585 10997 14598 11757
rect 14510 10940 14598 10997
rect 14510 10894 14539 10940
rect 14585 10894 14598 10940
rect 14510 10837 14598 10894
rect 14510 10791 14539 10837
rect 14585 10791 14598 10837
rect 14510 10734 14598 10791
rect 14510 10688 14539 10734
rect 14585 10688 14598 10734
rect 14510 10631 14598 10688
rect 14510 10585 14539 10631
rect 14585 10585 14598 10631
rect 14510 10528 14598 10585
rect 14510 10482 14539 10528
rect 14585 10482 14598 10528
rect 14510 10425 14598 10482
rect 14510 10379 14539 10425
rect 14585 10379 14598 10425
rect 14510 10322 14598 10379
rect 14510 10276 14539 10322
rect 14585 10276 14598 10322
rect 14510 10219 14598 10276
rect 14510 10173 14539 10219
rect 14585 10173 14598 10219
rect 14510 10116 14598 10173
rect 14510 10070 14539 10116
rect 14585 10070 14598 10116
rect 14510 10013 14598 10070
rect 14510 9967 14539 10013
rect 14585 9967 14598 10013
rect 14510 9954 14598 9967
rect 14750 11757 14838 11770
rect 14750 10997 14763 11757
rect 14809 10997 14838 11757
rect 14750 10940 14838 10997
rect 14750 10894 14763 10940
rect 14809 10894 14838 10940
rect 14750 10837 14838 10894
rect 14750 10791 14763 10837
rect 14809 10791 14838 10837
rect 14750 10734 14838 10791
rect 14750 10688 14763 10734
rect 14809 10688 14838 10734
rect 14750 10631 14838 10688
rect 14750 10585 14763 10631
rect 14809 10585 14838 10631
rect 14750 10528 14838 10585
rect 14750 10482 14763 10528
rect 14809 10482 14838 10528
rect 14750 10425 14838 10482
rect 14750 10379 14763 10425
rect 14809 10379 14838 10425
rect 14750 10322 14838 10379
rect 14750 10276 14763 10322
rect 14809 10276 14838 10322
rect 14750 10219 14838 10276
rect 14750 10173 14763 10219
rect 14809 10173 14838 10219
rect 14750 10116 14838 10173
rect 14750 10070 14763 10116
rect 14809 10070 14838 10116
rect 14750 10013 14838 10070
rect 14750 9967 14763 10013
rect 14809 9967 14838 10013
rect 14750 9954 14838 9967
rect 14958 11757 15062 11770
rect 14958 10997 14987 11757
rect 15033 10997 15062 11757
rect 14958 10940 15062 10997
rect 14958 10894 14987 10940
rect 15033 10894 15062 10940
rect 14958 10837 15062 10894
rect 14958 10791 14987 10837
rect 15033 10791 15062 10837
rect 14958 10734 15062 10791
rect 14958 10688 14987 10734
rect 15033 10688 15062 10734
rect 14958 10631 15062 10688
rect 14958 10585 14987 10631
rect 15033 10585 15062 10631
rect 14958 10528 15062 10585
rect 14958 10482 14987 10528
rect 15033 10482 15062 10528
rect 14958 10425 15062 10482
rect 14958 10379 14987 10425
rect 15033 10379 15062 10425
rect 14958 10322 15062 10379
rect 14958 10276 14987 10322
rect 15033 10276 15062 10322
rect 14958 10219 15062 10276
rect 14958 10173 14987 10219
rect 15033 10173 15062 10219
rect 14958 10116 15062 10173
rect 14958 10070 14987 10116
rect 15033 10070 15062 10116
rect 14958 10013 15062 10070
rect 14958 9967 14987 10013
rect 15033 9967 15062 10013
rect 14958 9954 15062 9967
rect 15182 11757 15286 11770
rect 15182 10997 15211 11757
rect 15257 10997 15286 11757
rect 15182 10940 15286 10997
rect 15182 10894 15211 10940
rect 15257 10894 15286 10940
rect 15182 10837 15286 10894
rect 15182 10791 15211 10837
rect 15257 10791 15286 10837
rect 15182 10734 15286 10791
rect 15182 10688 15211 10734
rect 15257 10688 15286 10734
rect 15182 10631 15286 10688
rect 15182 10585 15211 10631
rect 15257 10585 15286 10631
rect 15182 10528 15286 10585
rect 15182 10482 15211 10528
rect 15257 10482 15286 10528
rect 15182 10425 15286 10482
rect 15182 10379 15211 10425
rect 15257 10379 15286 10425
rect 15182 10322 15286 10379
rect 15182 10276 15211 10322
rect 15257 10276 15286 10322
rect 15182 10219 15286 10276
rect 15182 10173 15211 10219
rect 15257 10173 15286 10219
rect 15182 10116 15286 10173
rect 15182 10070 15211 10116
rect 15257 10070 15286 10116
rect 15182 10013 15286 10070
rect 15182 9967 15211 10013
rect 15257 9967 15286 10013
rect 15182 9954 15286 9967
rect 15406 11757 15510 11770
rect 15406 10997 15435 11757
rect 15481 10997 15510 11757
rect 15406 10940 15510 10997
rect 15406 10894 15435 10940
rect 15481 10894 15510 10940
rect 15406 10837 15510 10894
rect 15406 10791 15435 10837
rect 15481 10791 15510 10837
rect 15406 10734 15510 10791
rect 15406 10688 15435 10734
rect 15481 10688 15510 10734
rect 15406 10631 15510 10688
rect 15406 10585 15435 10631
rect 15481 10585 15510 10631
rect 15406 10528 15510 10585
rect 15406 10482 15435 10528
rect 15481 10482 15510 10528
rect 15406 10425 15510 10482
rect 15406 10379 15435 10425
rect 15481 10379 15510 10425
rect 15406 10322 15510 10379
rect 15406 10276 15435 10322
rect 15481 10276 15510 10322
rect 15406 10219 15510 10276
rect 15406 10173 15435 10219
rect 15481 10173 15510 10219
rect 15406 10116 15510 10173
rect 15406 10070 15435 10116
rect 15481 10070 15510 10116
rect 15406 10013 15510 10070
rect 15406 9967 15435 10013
rect 15481 9967 15510 10013
rect 15406 9954 15510 9967
rect 15630 11757 15718 11770
rect 15630 10997 15659 11757
rect 15705 10997 15718 11757
rect 15630 10940 15718 10997
rect 15630 10894 15659 10940
rect 15705 10894 15718 10940
rect 15630 10837 15718 10894
rect 15630 10791 15659 10837
rect 15705 10791 15718 10837
rect 15630 10734 15718 10791
rect 15630 10688 15659 10734
rect 15705 10688 15718 10734
rect 15630 10631 15718 10688
rect 15630 10585 15659 10631
rect 15705 10585 15718 10631
rect 15630 10528 15718 10585
rect 15630 10482 15659 10528
rect 15705 10482 15718 10528
rect 15630 10425 15718 10482
rect 15630 10379 15659 10425
rect 15705 10379 15718 10425
rect 15630 10322 15718 10379
rect 15630 10276 15659 10322
rect 15705 10276 15718 10322
rect 15630 10219 15718 10276
rect 15630 10173 15659 10219
rect 15705 10173 15718 10219
rect 15630 10116 15718 10173
rect 15630 10070 15659 10116
rect 15705 10070 15718 10116
rect 15630 10013 15718 10070
rect 15630 9967 15659 10013
rect 15705 9967 15718 10013
rect 15630 9954 15718 9967
rect 15870 11757 15958 11770
rect 15870 10997 15883 11757
rect 15929 10997 15958 11757
rect 15870 10940 15958 10997
rect 15870 10894 15883 10940
rect 15929 10894 15958 10940
rect 15870 10837 15958 10894
rect 15870 10791 15883 10837
rect 15929 10791 15958 10837
rect 15870 10734 15958 10791
rect 15870 10688 15883 10734
rect 15929 10688 15958 10734
rect 15870 10631 15958 10688
rect 15870 10585 15883 10631
rect 15929 10585 15958 10631
rect 15870 10528 15958 10585
rect 15870 10482 15883 10528
rect 15929 10482 15958 10528
rect 15870 10425 15958 10482
rect 15870 10379 15883 10425
rect 15929 10379 15958 10425
rect 15870 10322 15958 10379
rect 15870 10276 15883 10322
rect 15929 10276 15958 10322
rect 15870 10219 15958 10276
rect 15870 10173 15883 10219
rect 15929 10173 15958 10219
rect 15870 10116 15958 10173
rect 15870 10070 15883 10116
rect 15929 10070 15958 10116
rect 15870 10013 15958 10070
rect 15870 9967 15883 10013
rect 15929 9967 15958 10013
rect 15870 9954 15958 9967
rect 16078 11757 16182 11770
rect 16078 10997 16107 11757
rect 16153 10997 16182 11757
rect 16078 10940 16182 10997
rect 16078 10894 16107 10940
rect 16153 10894 16182 10940
rect 16078 10837 16182 10894
rect 16078 10791 16107 10837
rect 16153 10791 16182 10837
rect 16078 10734 16182 10791
rect 16078 10688 16107 10734
rect 16153 10688 16182 10734
rect 16078 10631 16182 10688
rect 16078 10585 16107 10631
rect 16153 10585 16182 10631
rect 16078 10528 16182 10585
rect 16078 10482 16107 10528
rect 16153 10482 16182 10528
rect 16078 10425 16182 10482
rect 16078 10379 16107 10425
rect 16153 10379 16182 10425
rect 16078 10322 16182 10379
rect 16078 10276 16107 10322
rect 16153 10276 16182 10322
rect 16078 10219 16182 10276
rect 16078 10173 16107 10219
rect 16153 10173 16182 10219
rect 16078 10116 16182 10173
rect 16078 10070 16107 10116
rect 16153 10070 16182 10116
rect 16078 10013 16182 10070
rect 16078 9967 16107 10013
rect 16153 9967 16182 10013
rect 16078 9954 16182 9967
rect 16302 11757 16406 11770
rect 16302 10997 16331 11757
rect 16377 10997 16406 11757
rect 16302 10940 16406 10997
rect 16302 10894 16331 10940
rect 16377 10894 16406 10940
rect 16302 10837 16406 10894
rect 16302 10791 16331 10837
rect 16377 10791 16406 10837
rect 16302 10734 16406 10791
rect 16302 10688 16331 10734
rect 16377 10688 16406 10734
rect 16302 10631 16406 10688
rect 16302 10585 16331 10631
rect 16377 10585 16406 10631
rect 16302 10528 16406 10585
rect 16302 10482 16331 10528
rect 16377 10482 16406 10528
rect 16302 10425 16406 10482
rect 16302 10379 16331 10425
rect 16377 10379 16406 10425
rect 16302 10322 16406 10379
rect 16302 10276 16331 10322
rect 16377 10276 16406 10322
rect 16302 10219 16406 10276
rect 16302 10173 16331 10219
rect 16377 10173 16406 10219
rect 16302 10116 16406 10173
rect 16302 10070 16331 10116
rect 16377 10070 16406 10116
rect 16302 10013 16406 10070
rect 16302 9967 16331 10013
rect 16377 9967 16406 10013
rect 16302 9954 16406 9967
rect 16526 11757 16630 11770
rect 16526 10997 16555 11757
rect 16601 10997 16630 11757
rect 16526 10940 16630 10997
rect 16526 10894 16555 10940
rect 16601 10894 16630 10940
rect 16526 10837 16630 10894
rect 16526 10791 16555 10837
rect 16601 10791 16630 10837
rect 16526 10734 16630 10791
rect 16526 10688 16555 10734
rect 16601 10688 16630 10734
rect 16526 10631 16630 10688
rect 16526 10585 16555 10631
rect 16601 10585 16630 10631
rect 16526 10528 16630 10585
rect 16526 10482 16555 10528
rect 16601 10482 16630 10528
rect 16526 10425 16630 10482
rect 16526 10379 16555 10425
rect 16601 10379 16630 10425
rect 16526 10322 16630 10379
rect 16526 10276 16555 10322
rect 16601 10276 16630 10322
rect 16526 10219 16630 10276
rect 16526 10173 16555 10219
rect 16601 10173 16630 10219
rect 16526 10116 16630 10173
rect 16526 10070 16555 10116
rect 16601 10070 16630 10116
rect 16526 10013 16630 10070
rect 16526 9967 16555 10013
rect 16601 9967 16630 10013
rect 16526 9954 16630 9967
rect 16750 11757 16838 11770
rect 16750 10997 16779 11757
rect 16825 10997 16838 11757
rect 16750 10940 16838 10997
rect 16750 10894 16779 10940
rect 16825 10894 16838 10940
rect 16750 10837 16838 10894
rect 16750 10791 16779 10837
rect 16825 10791 16838 10837
rect 16750 10734 16838 10791
rect 16750 10688 16779 10734
rect 16825 10688 16838 10734
rect 16750 10631 16838 10688
rect 16750 10585 16779 10631
rect 16825 10585 16838 10631
rect 16750 10528 16838 10585
rect 16750 10482 16779 10528
rect 16825 10482 16838 10528
rect 16750 10425 16838 10482
rect 16750 10379 16779 10425
rect 16825 10379 16838 10425
rect 16750 10322 16838 10379
rect 16750 10276 16779 10322
rect 16825 10276 16838 10322
rect 16750 10219 16838 10276
rect 16750 10173 16779 10219
rect 16825 10173 16838 10219
rect 16750 10116 16838 10173
rect 16750 10070 16779 10116
rect 16825 10070 16838 10116
rect 16750 10013 16838 10070
rect 16750 9967 16779 10013
rect 16825 9967 16838 10013
rect 16750 9954 16838 9967
rect 16990 11757 17078 11770
rect 16990 10997 17003 11757
rect 17049 10997 17078 11757
rect 16990 10940 17078 10997
rect 16990 10894 17003 10940
rect 17049 10894 17078 10940
rect 16990 10837 17078 10894
rect 16990 10791 17003 10837
rect 17049 10791 17078 10837
rect 16990 10734 17078 10791
rect 16990 10688 17003 10734
rect 17049 10688 17078 10734
rect 16990 10631 17078 10688
rect 16990 10585 17003 10631
rect 17049 10585 17078 10631
rect 16990 10528 17078 10585
rect 16990 10482 17003 10528
rect 17049 10482 17078 10528
rect 16990 10425 17078 10482
rect 16990 10379 17003 10425
rect 17049 10379 17078 10425
rect 16990 10322 17078 10379
rect 16990 10276 17003 10322
rect 17049 10276 17078 10322
rect 16990 10219 17078 10276
rect 16990 10173 17003 10219
rect 17049 10173 17078 10219
rect 16990 10116 17078 10173
rect 16990 10070 17003 10116
rect 17049 10070 17078 10116
rect 16990 10013 17078 10070
rect 16990 9967 17003 10013
rect 17049 9967 17078 10013
rect 16990 9954 17078 9967
rect 17198 11757 17302 11770
rect 17198 10997 17227 11757
rect 17273 10997 17302 11757
rect 17198 10940 17302 10997
rect 17198 10894 17227 10940
rect 17273 10894 17302 10940
rect 17198 10837 17302 10894
rect 17198 10791 17227 10837
rect 17273 10791 17302 10837
rect 17198 10734 17302 10791
rect 17198 10688 17227 10734
rect 17273 10688 17302 10734
rect 17198 10631 17302 10688
rect 17198 10585 17227 10631
rect 17273 10585 17302 10631
rect 17198 10528 17302 10585
rect 17198 10482 17227 10528
rect 17273 10482 17302 10528
rect 17198 10425 17302 10482
rect 17198 10379 17227 10425
rect 17273 10379 17302 10425
rect 17198 10322 17302 10379
rect 17198 10276 17227 10322
rect 17273 10276 17302 10322
rect 17198 10219 17302 10276
rect 17198 10173 17227 10219
rect 17273 10173 17302 10219
rect 17198 10116 17302 10173
rect 17198 10070 17227 10116
rect 17273 10070 17302 10116
rect 17198 10013 17302 10070
rect 17198 9967 17227 10013
rect 17273 9967 17302 10013
rect 17198 9954 17302 9967
rect 17422 11757 17526 11770
rect 17422 10997 17451 11757
rect 17497 10997 17526 11757
rect 17422 10940 17526 10997
rect 17422 10894 17451 10940
rect 17497 10894 17526 10940
rect 17422 10837 17526 10894
rect 17422 10791 17451 10837
rect 17497 10791 17526 10837
rect 17422 10734 17526 10791
rect 17422 10688 17451 10734
rect 17497 10688 17526 10734
rect 17422 10631 17526 10688
rect 17422 10585 17451 10631
rect 17497 10585 17526 10631
rect 17422 10528 17526 10585
rect 17422 10482 17451 10528
rect 17497 10482 17526 10528
rect 17422 10425 17526 10482
rect 17422 10379 17451 10425
rect 17497 10379 17526 10425
rect 17422 10322 17526 10379
rect 17422 10276 17451 10322
rect 17497 10276 17526 10322
rect 17422 10219 17526 10276
rect 17422 10173 17451 10219
rect 17497 10173 17526 10219
rect 17422 10116 17526 10173
rect 17422 10070 17451 10116
rect 17497 10070 17526 10116
rect 17422 10013 17526 10070
rect 17422 9967 17451 10013
rect 17497 9967 17526 10013
rect 17422 9954 17526 9967
rect 17646 11757 17750 11770
rect 17646 10997 17675 11757
rect 17721 10997 17750 11757
rect 17646 10940 17750 10997
rect 17646 10894 17675 10940
rect 17721 10894 17750 10940
rect 17646 10837 17750 10894
rect 17646 10791 17675 10837
rect 17721 10791 17750 10837
rect 17646 10734 17750 10791
rect 17646 10688 17675 10734
rect 17721 10688 17750 10734
rect 17646 10631 17750 10688
rect 17646 10585 17675 10631
rect 17721 10585 17750 10631
rect 17646 10528 17750 10585
rect 17646 10482 17675 10528
rect 17721 10482 17750 10528
rect 17646 10425 17750 10482
rect 17646 10379 17675 10425
rect 17721 10379 17750 10425
rect 17646 10322 17750 10379
rect 17646 10276 17675 10322
rect 17721 10276 17750 10322
rect 17646 10219 17750 10276
rect 17646 10173 17675 10219
rect 17721 10173 17750 10219
rect 17646 10116 17750 10173
rect 17646 10070 17675 10116
rect 17721 10070 17750 10116
rect 17646 10013 17750 10070
rect 17646 9967 17675 10013
rect 17721 9967 17750 10013
rect 17646 9954 17750 9967
rect 17870 11757 17958 11770
rect 17870 10997 17899 11757
rect 17945 10997 17958 11757
rect 17870 10940 17958 10997
rect 17870 10894 17899 10940
rect 17945 10894 17958 10940
rect 17870 10837 17958 10894
rect 17870 10791 17899 10837
rect 17945 10791 17958 10837
rect 17870 10734 17958 10791
rect 17870 10688 17899 10734
rect 17945 10688 17958 10734
rect 17870 10631 17958 10688
rect 17870 10585 17899 10631
rect 17945 10585 17958 10631
rect 17870 10528 17958 10585
rect 17870 10482 17899 10528
rect 17945 10482 17958 10528
rect 17870 10425 17958 10482
rect 17870 10379 17899 10425
rect 17945 10379 17958 10425
rect 17870 10322 17958 10379
rect 17870 10276 17899 10322
rect 17945 10276 17958 10322
rect 17870 10219 17958 10276
rect 17870 10173 17899 10219
rect 17945 10173 17958 10219
rect 17870 10116 17958 10173
rect 17870 10070 17899 10116
rect 17945 10070 17958 10116
rect 17870 10013 17958 10070
rect 17870 9967 17899 10013
rect 17945 9967 17958 10013
rect 17870 9954 17958 9967
rect 18110 11757 18198 11770
rect 18110 10997 18123 11757
rect 18169 10997 18198 11757
rect 18110 10940 18198 10997
rect 18110 10894 18123 10940
rect 18169 10894 18198 10940
rect 18110 10837 18198 10894
rect 18110 10791 18123 10837
rect 18169 10791 18198 10837
rect 18110 10734 18198 10791
rect 18110 10688 18123 10734
rect 18169 10688 18198 10734
rect 18110 10631 18198 10688
rect 18110 10585 18123 10631
rect 18169 10585 18198 10631
rect 18110 10528 18198 10585
rect 18110 10482 18123 10528
rect 18169 10482 18198 10528
rect 18110 10425 18198 10482
rect 18110 10379 18123 10425
rect 18169 10379 18198 10425
rect 18110 10322 18198 10379
rect 18110 10276 18123 10322
rect 18169 10276 18198 10322
rect 18110 10219 18198 10276
rect 18110 10173 18123 10219
rect 18169 10173 18198 10219
rect 18110 10116 18198 10173
rect 18110 10070 18123 10116
rect 18169 10070 18198 10116
rect 18110 10013 18198 10070
rect 18110 9967 18123 10013
rect 18169 9967 18198 10013
rect 18110 9954 18198 9967
rect 18318 11757 18422 11770
rect 18318 10997 18347 11757
rect 18393 10997 18422 11757
rect 18318 10940 18422 10997
rect 18318 10894 18347 10940
rect 18393 10894 18422 10940
rect 18318 10837 18422 10894
rect 18318 10791 18347 10837
rect 18393 10791 18422 10837
rect 18318 10734 18422 10791
rect 18318 10688 18347 10734
rect 18393 10688 18422 10734
rect 18318 10631 18422 10688
rect 18318 10585 18347 10631
rect 18393 10585 18422 10631
rect 18318 10528 18422 10585
rect 18318 10482 18347 10528
rect 18393 10482 18422 10528
rect 18318 10425 18422 10482
rect 18318 10379 18347 10425
rect 18393 10379 18422 10425
rect 18318 10322 18422 10379
rect 18318 10276 18347 10322
rect 18393 10276 18422 10322
rect 18318 10219 18422 10276
rect 18318 10173 18347 10219
rect 18393 10173 18422 10219
rect 18318 10116 18422 10173
rect 18318 10070 18347 10116
rect 18393 10070 18422 10116
rect 18318 10013 18422 10070
rect 18318 9967 18347 10013
rect 18393 9967 18422 10013
rect 18318 9954 18422 9967
rect 18542 11757 18646 11770
rect 18542 10997 18571 11757
rect 18617 10997 18646 11757
rect 18542 10940 18646 10997
rect 18542 10894 18571 10940
rect 18617 10894 18646 10940
rect 18542 10837 18646 10894
rect 18542 10791 18571 10837
rect 18617 10791 18646 10837
rect 18542 10734 18646 10791
rect 18542 10688 18571 10734
rect 18617 10688 18646 10734
rect 18542 10631 18646 10688
rect 18542 10585 18571 10631
rect 18617 10585 18646 10631
rect 18542 10528 18646 10585
rect 18542 10482 18571 10528
rect 18617 10482 18646 10528
rect 18542 10425 18646 10482
rect 18542 10379 18571 10425
rect 18617 10379 18646 10425
rect 18542 10322 18646 10379
rect 18542 10276 18571 10322
rect 18617 10276 18646 10322
rect 18542 10219 18646 10276
rect 18542 10173 18571 10219
rect 18617 10173 18646 10219
rect 18542 10116 18646 10173
rect 18542 10070 18571 10116
rect 18617 10070 18646 10116
rect 18542 10013 18646 10070
rect 18542 9967 18571 10013
rect 18617 9967 18646 10013
rect 18542 9954 18646 9967
rect 18766 11757 18870 11770
rect 18766 10997 18795 11757
rect 18841 10997 18870 11757
rect 18766 10940 18870 10997
rect 18766 10894 18795 10940
rect 18841 10894 18870 10940
rect 18766 10837 18870 10894
rect 18766 10791 18795 10837
rect 18841 10791 18870 10837
rect 18766 10734 18870 10791
rect 18766 10688 18795 10734
rect 18841 10688 18870 10734
rect 18766 10631 18870 10688
rect 18766 10585 18795 10631
rect 18841 10585 18870 10631
rect 18766 10528 18870 10585
rect 18766 10482 18795 10528
rect 18841 10482 18870 10528
rect 18766 10425 18870 10482
rect 18766 10379 18795 10425
rect 18841 10379 18870 10425
rect 18766 10322 18870 10379
rect 18766 10276 18795 10322
rect 18841 10276 18870 10322
rect 18766 10219 18870 10276
rect 18766 10173 18795 10219
rect 18841 10173 18870 10219
rect 18766 10116 18870 10173
rect 18766 10070 18795 10116
rect 18841 10070 18870 10116
rect 18766 10013 18870 10070
rect 18766 9967 18795 10013
rect 18841 9967 18870 10013
rect 18766 9954 18870 9967
rect 18990 11757 19078 11770
rect 18990 10997 19019 11757
rect 19065 10997 19078 11757
rect 18990 10940 19078 10997
rect 18990 10894 19019 10940
rect 19065 10894 19078 10940
rect 18990 10837 19078 10894
rect 18990 10791 19019 10837
rect 19065 10791 19078 10837
rect 18990 10734 19078 10791
rect 18990 10688 19019 10734
rect 19065 10688 19078 10734
rect 18990 10631 19078 10688
rect 18990 10585 19019 10631
rect 19065 10585 19078 10631
rect 18990 10528 19078 10585
rect 18990 10482 19019 10528
rect 19065 10482 19078 10528
rect 18990 10425 19078 10482
rect 18990 10379 19019 10425
rect 19065 10379 19078 10425
rect 18990 10322 19078 10379
rect 18990 10276 19019 10322
rect 19065 10276 19078 10322
rect 18990 10219 19078 10276
rect 18990 10173 19019 10219
rect 19065 10173 19078 10219
rect 18990 10116 19078 10173
rect 18990 10070 19019 10116
rect 19065 10070 19078 10116
rect 18990 10013 19078 10070
rect 18990 9967 19019 10013
rect 19065 9967 19078 10013
rect 18990 9954 19078 9967
rect 19230 11757 19318 11770
rect 19230 10997 19243 11757
rect 19289 10997 19318 11757
rect 19230 10940 19318 10997
rect 19230 10894 19243 10940
rect 19289 10894 19318 10940
rect 19230 10837 19318 10894
rect 19230 10791 19243 10837
rect 19289 10791 19318 10837
rect 19230 10734 19318 10791
rect 19230 10688 19243 10734
rect 19289 10688 19318 10734
rect 19230 10631 19318 10688
rect 19230 10585 19243 10631
rect 19289 10585 19318 10631
rect 19230 10528 19318 10585
rect 19230 10482 19243 10528
rect 19289 10482 19318 10528
rect 19230 10425 19318 10482
rect 19230 10379 19243 10425
rect 19289 10379 19318 10425
rect 19230 10322 19318 10379
rect 19230 10276 19243 10322
rect 19289 10276 19318 10322
rect 19230 10219 19318 10276
rect 19230 10173 19243 10219
rect 19289 10173 19318 10219
rect 19230 10116 19318 10173
rect 19230 10070 19243 10116
rect 19289 10070 19318 10116
rect 19230 10013 19318 10070
rect 19230 9967 19243 10013
rect 19289 9967 19318 10013
rect 19230 9954 19318 9967
rect 19438 11757 19542 11770
rect 19438 10997 19467 11757
rect 19513 10997 19542 11757
rect 19438 10940 19542 10997
rect 19438 10894 19467 10940
rect 19513 10894 19542 10940
rect 19438 10837 19542 10894
rect 19438 10791 19467 10837
rect 19513 10791 19542 10837
rect 19438 10734 19542 10791
rect 19438 10688 19467 10734
rect 19513 10688 19542 10734
rect 19438 10631 19542 10688
rect 19438 10585 19467 10631
rect 19513 10585 19542 10631
rect 19438 10528 19542 10585
rect 19438 10482 19467 10528
rect 19513 10482 19542 10528
rect 19438 10425 19542 10482
rect 19438 10379 19467 10425
rect 19513 10379 19542 10425
rect 19438 10322 19542 10379
rect 19438 10276 19467 10322
rect 19513 10276 19542 10322
rect 19438 10219 19542 10276
rect 19438 10173 19467 10219
rect 19513 10173 19542 10219
rect 19438 10116 19542 10173
rect 19438 10070 19467 10116
rect 19513 10070 19542 10116
rect 19438 10013 19542 10070
rect 19438 9967 19467 10013
rect 19513 9967 19542 10013
rect 19438 9954 19542 9967
rect 19662 11757 19766 11770
rect 19662 10997 19691 11757
rect 19737 10997 19766 11757
rect 19662 10940 19766 10997
rect 19662 10894 19691 10940
rect 19737 10894 19766 10940
rect 19662 10837 19766 10894
rect 19662 10791 19691 10837
rect 19737 10791 19766 10837
rect 19662 10734 19766 10791
rect 19662 10688 19691 10734
rect 19737 10688 19766 10734
rect 19662 10631 19766 10688
rect 19662 10585 19691 10631
rect 19737 10585 19766 10631
rect 19662 10528 19766 10585
rect 19662 10482 19691 10528
rect 19737 10482 19766 10528
rect 19662 10425 19766 10482
rect 19662 10379 19691 10425
rect 19737 10379 19766 10425
rect 19662 10322 19766 10379
rect 19662 10276 19691 10322
rect 19737 10276 19766 10322
rect 19662 10219 19766 10276
rect 19662 10173 19691 10219
rect 19737 10173 19766 10219
rect 19662 10116 19766 10173
rect 19662 10070 19691 10116
rect 19737 10070 19766 10116
rect 19662 10013 19766 10070
rect 19662 9967 19691 10013
rect 19737 9967 19766 10013
rect 19662 9954 19766 9967
rect 19886 11757 19974 11770
rect 19886 10997 19915 11757
rect 19961 10997 19974 11757
rect 19886 10940 19974 10997
rect 19886 10894 19915 10940
rect 19961 10894 19974 10940
rect 19886 10837 19974 10894
rect 19886 10791 19915 10837
rect 19961 10791 19974 10837
rect 19886 10734 19974 10791
rect 19886 10688 19915 10734
rect 19961 10688 19974 10734
rect 19886 10631 19974 10688
rect 19886 10585 19915 10631
rect 19961 10585 19974 10631
rect 19886 10528 19974 10585
rect 19886 10482 19915 10528
rect 19961 10482 19974 10528
rect 19886 10425 19974 10482
rect 19886 10379 19915 10425
rect 19961 10379 19974 10425
rect 19886 10322 19974 10379
rect 19886 10276 19915 10322
rect 19961 10276 19974 10322
rect 19886 10219 19974 10276
rect 19886 10173 19915 10219
rect 19961 10173 19974 10219
rect 19886 10116 19974 10173
rect 19886 10070 19915 10116
rect 19961 10070 19974 10116
rect 19886 10013 19974 10070
rect 19886 9967 19915 10013
rect 19961 9967 19974 10013
rect 19886 9954 19974 9967
rect 2608 9152 2696 9165
rect 2608 9106 2621 9152
rect 2667 9106 2696 9152
rect 2608 9048 2696 9106
rect 2608 9002 2621 9048
rect 2667 9002 2696 9048
rect 2608 8944 2696 9002
rect 2608 8898 2621 8944
rect 2667 8898 2696 8944
rect 2608 8840 2696 8898
rect 2608 8794 2621 8840
rect 2667 8794 2696 8840
rect 2608 8736 2696 8794
rect 2608 8690 2621 8736
rect 2667 8690 2696 8736
rect 2608 8631 2696 8690
rect 2608 8585 2621 8631
rect 2667 8585 2696 8631
rect 2608 8526 2696 8585
rect 2608 8480 2621 8526
rect 2667 8480 2696 8526
rect 2608 8421 2696 8480
rect 2608 8375 2621 8421
rect 2667 8375 2696 8421
rect 2608 8316 2696 8375
rect 2608 8270 2621 8316
rect 2667 8270 2696 8316
rect 2608 8257 2696 8270
rect 2816 9152 2904 9165
rect 2816 9106 2845 9152
rect 2891 9106 2904 9152
rect 2816 9048 2904 9106
rect 2816 9002 2845 9048
rect 2891 9002 2904 9048
rect 2816 8944 2904 9002
rect 2816 8898 2845 8944
rect 2891 8898 2904 8944
rect 2816 8840 2904 8898
rect 2816 8794 2845 8840
rect 2891 8794 2904 8840
rect 2816 8736 2904 8794
rect 2816 8690 2845 8736
rect 2891 8690 2904 8736
rect 2816 8631 2904 8690
rect 2816 8585 2845 8631
rect 2891 8585 2904 8631
rect 2816 8526 2904 8585
rect 2816 8480 2845 8526
rect 2891 8480 2904 8526
rect 2816 8421 2904 8480
rect 2816 8375 2845 8421
rect 2891 8375 2904 8421
rect 2816 8316 2904 8375
rect 2816 8270 2845 8316
rect 2891 8270 2904 8316
rect 2816 8257 2904 8270
rect 3122 9152 3210 9165
rect 3122 9106 3135 9152
rect 3181 9106 3210 9152
rect 3122 9048 3210 9106
rect 3122 9002 3135 9048
rect 3181 9002 3210 9048
rect 3122 8944 3210 9002
rect 3122 8898 3135 8944
rect 3181 8898 3210 8944
rect 3122 8840 3210 8898
rect 3122 8794 3135 8840
rect 3181 8794 3210 8840
rect 3122 8736 3210 8794
rect 3122 8690 3135 8736
rect 3181 8690 3210 8736
rect 3122 8631 3210 8690
rect 3122 8585 3135 8631
rect 3181 8585 3210 8631
rect 3122 8526 3210 8585
rect 3122 8480 3135 8526
rect 3181 8480 3210 8526
rect 3122 8421 3210 8480
rect 3122 8375 3135 8421
rect 3181 8375 3210 8421
rect 3122 8316 3210 8375
rect 3122 8270 3135 8316
rect 3181 8270 3210 8316
rect 3122 8257 3210 8270
rect 3330 9152 3418 9165
rect 3330 9106 3359 9152
rect 3405 9106 3418 9152
rect 3330 9048 3418 9106
rect 3330 9002 3359 9048
rect 3405 9002 3418 9048
rect 3330 8944 3418 9002
rect 3330 8898 3359 8944
rect 3405 8898 3418 8944
rect 3330 8840 3418 8898
rect 3330 8794 3359 8840
rect 3405 8794 3418 8840
rect 3330 8736 3418 8794
rect 3330 8690 3359 8736
rect 3405 8690 3418 8736
rect 3330 8631 3418 8690
rect 3330 8585 3359 8631
rect 3405 8585 3418 8631
rect 3330 8526 3418 8585
rect 3330 8480 3359 8526
rect 3405 8480 3418 8526
rect 4299 9152 4387 9165
rect 4299 9106 4312 9152
rect 4358 9106 4387 9152
rect 4299 9048 4387 9106
rect 4299 9002 4312 9048
rect 4358 9002 4387 9048
rect 4299 8944 4387 9002
rect 4299 8898 4312 8944
rect 4358 8898 4387 8944
rect 4299 8840 4387 8898
rect 4299 8794 4312 8840
rect 4358 8794 4387 8840
rect 4299 8736 4387 8794
rect 4299 8690 4312 8736
rect 4358 8690 4387 8736
rect 4299 8631 4387 8690
rect 4299 8585 4312 8631
rect 4358 8585 4387 8631
rect 4299 8526 4387 8585
rect 3330 8421 3418 8480
rect 3330 8375 3359 8421
rect 3405 8375 3418 8421
rect 3330 8316 3418 8375
rect 3330 8270 3359 8316
rect 3405 8270 3418 8316
rect 3330 8257 3418 8270
rect 4299 8480 4312 8526
rect 4358 8480 4387 8526
rect 4299 8421 4387 8480
rect 4299 8375 4312 8421
rect 4358 8375 4387 8421
rect 4299 8316 4387 8375
rect 4299 8270 4312 8316
rect 4358 8270 4387 8316
rect 4299 8257 4387 8270
rect 4507 9152 4595 9165
rect 4507 9106 4536 9152
rect 4582 9106 4595 9152
rect 4507 9048 4595 9106
rect 4507 9002 4536 9048
rect 4582 9002 4595 9048
rect 4507 8944 4595 9002
rect 4507 8898 4536 8944
rect 4582 8898 4595 8944
rect 4507 8840 4595 8898
rect 4507 8794 4536 8840
rect 4582 8794 4595 8840
rect 4507 8736 4595 8794
rect 4507 8690 4536 8736
rect 4582 8690 4595 8736
rect 4507 8631 4595 8690
rect 4507 8585 4536 8631
rect 4582 8585 4595 8631
rect 4507 8526 4595 8585
rect 4507 8480 4536 8526
rect 4582 8480 4595 8526
rect 4507 8421 4595 8480
rect 4507 8375 4536 8421
rect 4582 8375 4595 8421
rect 4507 8316 4595 8375
rect 4507 8270 4536 8316
rect 4582 8270 4595 8316
rect 4507 8257 4595 8270
rect 4813 9152 4901 9165
rect 4813 9106 4826 9152
rect 4872 9106 4901 9152
rect 4813 9048 4901 9106
rect 4813 9002 4826 9048
rect 4872 9002 4901 9048
rect 4813 8944 4901 9002
rect 4813 8898 4826 8944
rect 4872 8898 4901 8944
rect 4813 8840 4901 8898
rect 4813 8794 4826 8840
rect 4872 8794 4901 8840
rect 4813 8736 4901 8794
rect 4813 8690 4826 8736
rect 4872 8690 4901 8736
rect 4813 8631 4901 8690
rect 4813 8585 4826 8631
rect 4872 8585 4901 8631
rect 4813 8526 4901 8585
rect 4813 8480 4826 8526
rect 4872 8480 4901 8526
rect 4813 8421 4901 8480
rect 4813 8375 4826 8421
rect 4872 8375 4901 8421
rect 4813 8316 4901 8375
rect 4813 8270 4826 8316
rect 4872 8270 4901 8316
rect 4813 8257 4901 8270
rect 5021 9152 5109 9165
rect 5021 9106 5050 9152
rect 5096 9106 5109 9152
rect 5021 9048 5109 9106
rect 5021 9002 5050 9048
rect 5096 9002 5109 9048
rect 5021 8944 5109 9002
rect 5021 8898 5050 8944
rect 5096 8898 5109 8944
rect 5021 8840 5109 8898
rect 5021 8794 5050 8840
rect 5096 8794 5109 8840
rect 5021 8736 5109 8794
rect 5021 8690 5050 8736
rect 5096 8690 5109 8736
rect 5021 8631 5109 8690
rect 5021 8585 5050 8631
rect 5096 8585 5109 8631
rect 5021 8526 5109 8585
rect 5021 8480 5050 8526
rect 5096 8480 5109 8526
rect 5990 9152 6078 9165
rect 5990 9106 6003 9152
rect 6049 9106 6078 9152
rect 5990 9048 6078 9106
rect 5990 9002 6003 9048
rect 6049 9002 6078 9048
rect 5990 8944 6078 9002
rect 5990 8898 6003 8944
rect 6049 8898 6078 8944
rect 5990 8840 6078 8898
rect 5990 8794 6003 8840
rect 6049 8794 6078 8840
rect 5990 8736 6078 8794
rect 5990 8690 6003 8736
rect 6049 8690 6078 8736
rect 5990 8631 6078 8690
rect 5990 8585 6003 8631
rect 6049 8585 6078 8631
rect 5990 8526 6078 8585
rect 5021 8421 5109 8480
rect 5021 8375 5050 8421
rect 5096 8375 5109 8421
rect 5021 8316 5109 8375
rect 5021 8270 5050 8316
rect 5096 8270 5109 8316
rect 5021 8257 5109 8270
rect 5990 8480 6003 8526
rect 6049 8480 6078 8526
rect 5990 8421 6078 8480
rect 5990 8375 6003 8421
rect 6049 8375 6078 8421
rect 5990 8316 6078 8375
rect 5990 8270 6003 8316
rect 6049 8270 6078 8316
rect 5990 8257 6078 8270
rect 6198 9152 6286 9165
rect 6198 9106 6227 9152
rect 6273 9106 6286 9152
rect 6198 9048 6286 9106
rect 6198 9002 6227 9048
rect 6273 9002 6286 9048
rect 6198 8944 6286 9002
rect 6198 8898 6227 8944
rect 6273 8898 6286 8944
rect 6198 8840 6286 8898
rect 6198 8794 6227 8840
rect 6273 8794 6286 8840
rect 6198 8736 6286 8794
rect 6198 8690 6227 8736
rect 6273 8690 6286 8736
rect 6198 8631 6286 8690
rect 6198 8585 6227 8631
rect 6273 8585 6286 8631
rect 6198 8526 6286 8585
rect 6198 8480 6227 8526
rect 6273 8480 6286 8526
rect 6198 8421 6286 8480
rect 6198 8375 6227 8421
rect 6273 8375 6286 8421
rect 6198 8316 6286 8375
rect 6198 8270 6227 8316
rect 6273 8270 6286 8316
rect 6198 8257 6286 8270
rect 6504 9152 6592 9165
rect 6504 9106 6517 9152
rect 6563 9106 6592 9152
rect 6504 9048 6592 9106
rect 6504 9002 6517 9048
rect 6563 9002 6592 9048
rect 6504 8944 6592 9002
rect 6504 8898 6517 8944
rect 6563 8898 6592 8944
rect 6504 8840 6592 8898
rect 6504 8794 6517 8840
rect 6563 8794 6592 8840
rect 6504 8736 6592 8794
rect 6504 8690 6517 8736
rect 6563 8690 6592 8736
rect 6504 8631 6592 8690
rect 6504 8585 6517 8631
rect 6563 8585 6592 8631
rect 6504 8526 6592 8585
rect 6504 8480 6517 8526
rect 6563 8480 6592 8526
rect 6504 8421 6592 8480
rect 6504 8375 6517 8421
rect 6563 8375 6592 8421
rect 6504 8316 6592 8375
rect 6504 8270 6517 8316
rect 6563 8270 6592 8316
rect 6504 8257 6592 8270
rect 6712 9152 6800 9165
rect 6712 9106 6741 9152
rect 6787 9106 6800 9152
rect 6712 9048 6800 9106
rect 6712 9002 6741 9048
rect 6787 9002 6800 9048
rect 6712 8944 6800 9002
rect 6712 8898 6741 8944
rect 6787 8898 6800 8944
rect 6712 8840 6800 8898
rect 6712 8794 6741 8840
rect 6787 8794 6800 8840
rect 6712 8736 6800 8794
rect 6712 8690 6741 8736
rect 6787 8690 6800 8736
rect 6712 8631 6800 8690
rect 6712 8585 6741 8631
rect 6787 8585 6800 8631
rect 6712 8526 6800 8585
rect 7437 9008 7525 9021
rect 7437 8962 7450 9008
rect 7496 8962 7525 9008
rect 7437 8880 7525 8962
rect 7437 8834 7450 8880
rect 7496 8834 7525 8880
rect 7437 8753 7525 8834
rect 7437 8707 7450 8753
rect 7496 8707 7525 8753
rect 7437 8626 7525 8707
rect 7437 8580 7450 8626
rect 7496 8580 7525 8626
rect 7437 8567 7525 8580
rect 7645 9008 7749 9021
rect 7645 8962 7674 9008
rect 7720 8962 7749 9008
rect 7645 8880 7749 8962
rect 7645 8834 7674 8880
rect 7720 8834 7749 8880
rect 7645 8753 7749 8834
rect 7645 8707 7674 8753
rect 7720 8707 7749 8753
rect 7645 8626 7749 8707
rect 7645 8580 7674 8626
rect 7720 8580 7749 8626
rect 7645 8567 7749 8580
rect 7869 9008 7973 9021
rect 7869 8962 7898 9008
rect 7944 8962 7973 9008
rect 7869 8880 7973 8962
rect 7869 8834 7898 8880
rect 7944 8834 7973 8880
rect 7869 8753 7973 8834
rect 7869 8707 7898 8753
rect 7944 8707 7973 8753
rect 7869 8626 7973 8707
rect 7869 8580 7898 8626
rect 7944 8580 7973 8626
rect 7869 8567 7973 8580
rect 8093 9008 8197 9021
rect 8093 8962 8122 9008
rect 8168 8962 8197 9008
rect 8093 8880 8197 8962
rect 8093 8834 8122 8880
rect 8168 8834 8197 8880
rect 8093 8753 8197 8834
rect 8093 8707 8122 8753
rect 8168 8707 8197 8753
rect 8093 8626 8197 8707
rect 8093 8580 8122 8626
rect 8168 8580 8197 8626
rect 8093 8567 8197 8580
rect 8317 9008 8421 9021
rect 8317 8962 8346 9008
rect 8392 8962 8421 9008
rect 8317 8880 8421 8962
rect 8317 8834 8346 8880
rect 8392 8834 8421 8880
rect 8317 8753 8421 8834
rect 8317 8707 8346 8753
rect 8392 8707 8421 8753
rect 8317 8626 8421 8707
rect 8317 8580 8346 8626
rect 8392 8580 8421 8626
rect 8317 8567 8421 8580
rect 8541 9008 8645 9021
rect 8541 8962 8570 9008
rect 8616 8962 8645 9008
rect 8541 8880 8645 8962
rect 8541 8834 8570 8880
rect 8616 8834 8645 8880
rect 8541 8753 8645 8834
rect 8541 8707 8570 8753
rect 8616 8707 8645 8753
rect 8541 8626 8645 8707
rect 8541 8580 8570 8626
rect 8616 8580 8645 8626
rect 8541 8567 8645 8580
rect 8765 9008 8853 9021
rect 8765 8962 8794 9008
rect 8840 8962 8853 9008
rect 8765 8880 8853 8962
rect 8765 8834 8794 8880
rect 8840 8834 8853 8880
rect 8765 8753 8853 8834
rect 8765 8707 8794 8753
rect 8840 8707 8853 8753
rect 8765 8626 8853 8707
rect 8765 8580 8794 8626
rect 8840 8580 8853 8626
rect 8765 8567 8853 8580
rect 9070 9008 9158 9021
rect 9070 8962 9083 9008
rect 9129 8962 9158 9008
rect 9070 8880 9158 8962
rect 9070 8834 9083 8880
rect 9129 8834 9158 8880
rect 9070 8753 9158 8834
rect 9070 8707 9083 8753
rect 9129 8707 9158 8753
rect 9070 8626 9158 8707
rect 9070 8580 9083 8626
rect 9129 8580 9158 8626
rect 9070 8567 9158 8580
rect 9278 9008 9382 9021
rect 9278 8962 9307 9008
rect 9353 8962 9382 9008
rect 9278 8880 9382 8962
rect 9278 8834 9307 8880
rect 9353 8834 9382 8880
rect 9278 8753 9382 8834
rect 9278 8707 9307 8753
rect 9353 8707 9382 8753
rect 9278 8626 9382 8707
rect 9278 8580 9307 8626
rect 9353 8580 9382 8626
rect 9278 8567 9382 8580
rect 9502 9008 9606 9021
rect 9502 8962 9531 9008
rect 9577 8962 9606 9008
rect 9502 8880 9606 8962
rect 9502 8834 9531 8880
rect 9577 8834 9606 8880
rect 9502 8753 9606 8834
rect 9502 8707 9531 8753
rect 9577 8707 9606 8753
rect 9502 8626 9606 8707
rect 9502 8580 9531 8626
rect 9577 8580 9606 8626
rect 9502 8567 9606 8580
rect 9726 9008 9830 9021
rect 9726 8962 9755 9008
rect 9801 8962 9830 9008
rect 9726 8880 9830 8962
rect 9726 8834 9755 8880
rect 9801 8834 9830 8880
rect 9726 8753 9830 8834
rect 9726 8707 9755 8753
rect 9801 8707 9830 8753
rect 9726 8626 9830 8707
rect 9726 8580 9755 8626
rect 9801 8580 9830 8626
rect 9726 8567 9830 8580
rect 9950 9008 10054 9021
rect 9950 8962 9979 9008
rect 10025 8962 10054 9008
rect 9950 8880 10054 8962
rect 9950 8834 9979 8880
rect 10025 8834 10054 8880
rect 9950 8753 10054 8834
rect 9950 8707 9979 8753
rect 10025 8707 10054 8753
rect 9950 8626 10054 8707
rect 9950 8580 9979 8626
rect 10025 8580 10054 8626
rect 9950 8567 10054 8580
rect 10174 9008 10278 9021
rect 10174 8962 10203 9008
rect 10249 8962 10278 9008
rect 10174 8880 10278 8962
rect 10174 8834 10203 8880
rect 10249 8834 10278 8880
rect 10174 8753 10278 8834
rect 10174 8707 10203 8753
rect 10249 8707 10278 8753
rect 10174 8626 10278 8707
rect 10174 8580 10203 8626
rect 10249 8580 10278 8626
rect 10174 8567 10278 8580
rect 10398 9008 10486 9021
rect 10398 8962 10427 9008
rect 10473 8962 10486 9008
rect 10398 8880 10486 8962
rect 10398 8834 10427 8880
rect 10473 8834 10486 8880
rect 10398 8753 10486 8834
rect 10398 8707 10427 8753
rect 10473 8707 10486 8753
rect 10398 8626 10486 8707
rect 10398 8580 10427 8626
rect 10473 8580 10486 8626
rect 10398 8567 10486 8580
rect 10704 9008 10792 9021
rect 10704 8962 10717 9008
rect 10763 8962 10792 9008
rect 10704 8880 10792 8962
rect 10704 8834 10717 8880
rect 10763 8834 10792 8880
rect 10704 8753 10792 8834
rect 10704 8707 10717 8753
rect 10763 8707 10792 8753
rect 10704 8626 10792 8707
rect 10704 8580 10717 8626
rect 10763 8580 10792 8626
rect 10704 8567 10792 8580
rect 10912 9008 11016 9021
rect 10912 8962 10941 9008
rect 10987 8962 11016 9008
rect 10912 8880 11016 8962
rect 10912 8834 10941 8880
rect 10987 8834 11016 8880
rect 10912 8753 11016 8834
rect 10912 8707 10941 8753
rect 10987 8707 11016 8753
rect 10912 8626 11016 8707
rect 10912 8580 10941 8626
rect 10987 8580 11016 8626
rect 10912 8567 11016 8580
rect 11136 9008 11240 9021
rect 11136 8962 11165 9008
rect 11211 8962 11240 9008
rect 11136 8880 11240 8962
rect 11136 8834 11165 8880
rect 11211 8834 11240 8880
rect 11136 8753 11240 8834
rect 11136 8707 11165 8753
rect 11211 8707 11240 8753
rect 11136 8626 11240 8707
rect 11136 8580 11165 8626
rect 11211 8580 11240 8626
rect 11136 8567 11240 8580
rect 11360 9008 11464 9021
rect 11360 8962 11389 9008
rect 11435 8962 11464 9008
rect 11360 8880 11464 8962
rect 11360 8834 11389 8880
rect 11435 8834 11464 8880
rect 11360 8753 11464 8834
rect 11360 8707 11389 8753
rect 11435 8707 11464 8753
rect 11360 8626 11464 8707
rect 11360 8580 11389 8626
rect 11435 8580 11464 8626
rect 11360 8567 11464 8580
rect 11584 9008 11688 9021
rect 11584 8962 11613 9008
rect 11659 8962 11688 9008
rect 11584 8880 11688 8962
rect 11584 8834 11613 8880
rect 11659 8834 11688 8880
rect 11584 8753 11688 8834
rect 11584 8707 11613 8753
rect 11659 8707 11688 8753
rect 11584 8626 11688 8707
rect 11584 8580 11613 8626
rect 11659 8580 11688 8626
rect 11584 8567 11688 8580
rect 11808 9008 11912 9021
rect 11808 8962 11837 9008
rect 11883 8962 11912 9008
rect 11808 8880 11912 8962
rect 11808 8834 11837 8880
rect 11883 8834 11912 8880
rect 11808 8753 11912 8834
rect 11808 8707 11837 8753
rect 11883 8707 11912 8753
rect 11808 8626 11912 8707
rect 11808 8580 11837 8626
rect 11883 8580 11912 8626
rect 11808 8567 11912 8580
rect 12032 9008 12120 9021
rect 12032 8962 12061 9008
rect 12107 8962 12120 9008
rect 12032 8880 12120 8962
rect 12032 8834 12061 8880
rect 12107 8834 12120 8880
rect 12032 8753 12120 8834
rect 12032 8707 12061 8753
rect 12107 8707 12120 8753
rect 12032 8626 12120 8707
rect 12032 8580 12061 8626
rect 12107 8580 12120 8626
rect 12032 8567 12120 8580
rect 12338 9008 12426 9021
rect 12338 8962 12351 9008
rect 12397 8962 12426 9008
rect 12338 8880 12426 8962
rect 12338 8834 12351 8880
rect 12397 8834 12426 8880
rect 12338 8753 12426 8834
rect 12338 8707 12351 8753
rect 12397 8707 12426 8753
rect 12338 8626 12426 8707
rect 12338 8580 12351 8626
rect 12397 8580 12426 8626
rect 12338 8567 12426 8580
rect 12546 9008 12650 9021
rect 12546 8962 12575 9008
rect 12621 8962 12650 9008
rect 12546 8880 12650 8962
rect 12546 8834 12575 8880
rect 12621 8834 12650 8880
rect 12546 8753 12650 8834
rect 12546 8707 12575 8753
rect 12621 8707 12650 8753
rect 12546 8626 12650 8707
rect 12546 8580 12575 8626
rect 12621 8580 12650 8626
rect 12546 8567 12650 8580
rect 12770 9008 12874 9021
rect 12770 8962 12799 9008
rect 12845 8962 12874 9008
rect 12770 8880 12874 8962
rect 12770 8834 12799 8880
rect 12845 8834 12874 8880
rect 12770 8753 12874 8834
rect 12770 8707 12799 8753
rect 12845 8707 12874 8753
rect 12770 8626 12874 8707
rect 12770 8580 12799 8626
rect 12845 8580 12874 8626
rect 12770 8567 12874 8580
rect 12994 9008 13098 9021
rect 12994 8962 13023 9008
rect 13069 8962 13098 9008
rect 12994 8880 13098 8962
rect 12994 8834 13023 8880
rect 13069 8834 13098 8880
rect 12994 8753 13098 8834
rect 12994 8707 13023 8753
rect 13069 8707 13098 8753
rect 12994 8626 13098 8707
rect 12994 8580 13023 8626
rect 13069 8580 13098 8626
rect 12994 8567 13098 8580
rect 13218 9008 13322 9021
rect 13218 8962 13247 9008
rect 13293 8962 13322 9008
rect 13218 8880 13322 8962
rect 13218 8834 13247 8880
rect 13293 8834 13322 8880
rect 13218 8753 13322 8834
rect 13218 8707 13247 8753
rect 13293 8707 13322 8753
rect 13218 8626 13322 8707
rect 13218 8580 13247 8626
rect 13293 8580 13322 8626
rect 13218 8567 13322 8580
rect 13442 9008 13546 9021
rect 13442 8962 13471 9008
rect 13517 8962 13546 9008
rect 13442 8880 13546 8962
rect 13442 8834 13471 8880
rect 13517 8834 13546 8880
rect 13442 8753 13546 8834
rect 13442 8707 13471 8753
rect 13517 8707 13546 8753
rect 13442 8626 13546 8707
rect 13442 8580 13471 8626
rect 13517 8580 13546 8626
rect 13442 8567 13546 8580
rect 13666 9008 13754 9021
rect 13666 8962 13695 9008
rect 13741 8962 13754 9008
rect 13666 8880 13754 8962
rect 13666 8834 13695 8880
rect 13741 8834 13754 8880
rect 13666 8753 13754 8834
rect 13666 8707 13695 8753
rect 13741 8707 13754 8753
rect 13666 8626 13754 8707
rect 13666 8580 13695 8626
rect 13741 8580 13754 8626
rect 13666 8567 13754 8580
rect 6712 8480 6741 8526
rect 6787 8480 6800 8526
rect 6712 8421 6800 8480
rect 6712 8375 6741 8421
rect 6787 8375 6800 8421
rect 6712 8316 6800 8375
rect 6712 8270 6741 8316
rect 6787 8270 6800 8316
rect 6712 8257 6800 8270
rect 7407 3866 7526 3912
rect 7407 3820 7450 3866
rect 7496 3820 7526 3866
rect 7407 3698 7526 3820
rect 7407 3652 7450 3698
rect 7496 3652 7526 3698
rect 7407 3530 7526 3652
rect 7407 3484 7450 3530
rect 7496 3484 7526 3530
rect 7407 3363 7526 3484
rect 7407 3317 7450 3363
rect 7496 3317 7526 3363
rect 7407 3195 7526 3317
rect 7407 3149 7450 3195
rect 7496 3149 7526 3195
rect 7407 3027 7526 3149
rect 7407 2981 7450 3027
rect 7496 2981 7526 3027
rect 7407 2859 7526 2981
rect 7407 2813 7450 2859
rect 7496 2813 7526 2859
rect 7407 2692 7526 2813
rect 7407 2646 7450 2692
rect 7496 2646 7526 2692
rect 7407 2550 7526 2646
rect 7646 2550 7748 3912
rect 7868 2550 7972 3912
rect 8092 3866 8198 3912
rect 8092 3820 8122 3866
rect 8168 3820 8198 3866
rect 8092 3698 8198 3820
rect 8092 3652 8122 3698
rect 8168 3652 8198 3698
rect 8092 3530 8198 3652
rect 8092 3484 8122 3530
rect 8168 3484 8198 3530
rect 8092 3363 8198 3484
rect 8092 3317 8122 3363
rect 8168 3317 8198 3363
rect 8092 3195 8198 3317
rect 8092 3149 8122 3195
rect 8168 3149 8198 3195
rect 8092 3027 8198 3149
rect 8092 2981 8122 3027
rect 8168 2981 8198 3027
rect 8092 2859 8198 2981
rect 8092 2813 8122 2859
rect 8168 2813 8198 2859
rect 8092 2692 8198 2813
rect 8092 2646 8122 2692
rect 8168 2646 8198 2692
rect 8092 2550 8198 2646
rect 8318 2550 8422 3912
rect 8542 2550 8644 3912
rect 8764 3866 8883 3912
rect 8764 3820 8794 3866
rect 8840 3820 8883 3866
rect 8764 3698 8883 3820
rect 8764 3652 8794 3698
rect 8840 3652 8883 3698
rect 8764 3530 8883 3652
rect 8764 3484 8794 3530
rect 8840 3484 8883 3530
rect 8764 3363 8883 3484
rect 8764 3317 8794 3363
rect 8840 3317 8883 3363
rect 8764 3195 8883 3317
rect 8764 3149 8794 3195
rect 8840 3149 8883 3195
rect 8764 3027 8883 3149
rect 8764 2981 8794 3027
rect 8840 2981 8883 3027
rect 8764 2859 8883 2981
rect 8764 2813 8794 2859
rect 8840 2813 8883 2859
rect 8764 2692 8883 2813
rect 8764 2646 8794 2692
rect 8840 2646 8883 2692
rect 8764 2550 8883 2646
rect 9040 3866 9159 3912
rect 9040 3820 9083 3866
rect 9129 3820 9159 3866
rect 9040 3698 9159 3820
rect 9040 3652 9083 3698
rect 9129 3652 9159 3698
rect 9040 3530 9159 3652
rect 9040 3484 9083 3530
rect 9129 3484 9159 3530
rect 9040 3363 9159 3484
rect 9040 3317 9083 3363
rect 9129 3317 9159 3363
rect 9040 3195 9159 3317
rect 9040 3149 9083 3195
rect 9129 3149 9159 3195
rect 9040 3027 9159 3149
rect 9040 2981 9083 3027
rect 9129 2981 9159 3027
rect 9040 2859 9159 2981
rect 9040 2813 9083 2859
rect 9129 2813 9159 2859
rect 9040 2692 9159 2813
rect 9040 2646 9083 2692
rect 9129 2646 9159 2692
rect 9040 2550 9159 2646
rect 9279 2550 9381 3912
rect 9501 2550 9605 3912
rect 9725 3866 9831 3912
rect 9725 3820 9755 3866
rect 9801 3820 9831 3866
rect 9725 3698 9831 3820
rect 9725 3652 9755 3698
rect 9801 3652 9831 3698
rect 9725 3530 9831 3652
rect 9725 3484 9755 3530
rect 9801 3484 9831 3530
rect 9725 3363 9831 3484
rect 9725 3317 9755 3363
rect 9801 3317 9831 3363
rect 9725 3195 9831 3317
rect 9725 3149 9755 3195
rect 9801 3149 9831 3195
rect 9725 3027 9831 3149
rect 9725 2981 9755 3027
rect 9801 2981 9831 3027
rect 9725 2859 9831 2981
rect 9725 2813 9755 2859
rect 9801 2813 9831 2859
rect 9725 2692 9831 2813
rect 9725 2646 9755 2692
rect 9801 2646 9831 2692
rect 9725 2550 9831 2646
rect 9951 2550 10055 3912
rect 10175 2550 10277 3912
rect 10397 3866 10516 3912
rect 10397 3820 10427 3866
rect 10473 3820 10516 3866
rect 10397 3698 10516 3820
rect 10397 3652 10427 3698
rect 10473 3652 10516 3698
rect 10397 3530 10516 3652
rect 10397 3484 10427 3530
rect 10473 3484 10516 3530
rect 10397 3363 10516 3484
rect 10397 3317 10427 3363
rect 10473 3317 10516 3363
rect 10397 3195 10516 3317
rect 10397 3149 10427 3195
rect 10473 3149 10516 3195
rect 10397 3027 10516 3149
rect 10397 2981 10427 3027
rect 10473 2981 10516 3027
rect 10397 2859 10516 2981
rect 10397 2813 10427 2859
rect 10473 2813 10516 2859
rect 10397 2692 10516 2813
rect 10397 2646 10427 2692
rect 10473 2646 10516 2692
rect 10397 2550 10516 2646
rect 10674 3866 10793 3912
rect 10674 3820 10717 3866
rect 10763 3820 10793 3866
rect 10674 3698 10793 3820
rect 10674 3652 10717 3698
rect 10763 3652 10793 3698
rect 10674 3530 10793 3652
rect 10674 3484 10717 3530
rect 10763 3484 10793 3530
rect 10674 3363 10793 3484
rect 10674 3317 10717 3363
rect 10763 3317 10793 3363
rect 10674 3195 10793 3317
rect 10674 3149 10717 3195
rect 10763 3149 10793 3195
rect 10674 3027 10793 3149
rect 10674 2981 10717 3027
rect 10763 2981 10793 3027
rect 10674 2859 10793 2981
rect 10674 2813 10717 2859
rect 10763 2813 10793 2859
rect 10674 2692 10793 2813
rect 10674 2646 10717 2692
rect 10763 2646 10793 2692
rect 10674 2550 10793 2646
rect 10913 2550 11015 3912
rect 11135 2550 11239 3912
rect 11359 3866 11465 3912
rect 11359 3820 11389 3866
rect 11435 3820 11465 3866
rect 11359 3698 11465 3820
rect 11359 3652 11389 3698
rect 11435 3652 11465 3698
rect 11359 3530 11465 3652
rect 11359 3484 11389 3530
rect 11435 3484 11465 3530
rect 11359 3363 11465 3484
rect 11359 3317 11389 3363
rect 11435 3317 11465 3363
rect 11359 3195 11465 3317
rect 11359 3149 11389 3195
rect 11435 3149 11465 3195
rect 11359 3027 11465 3149
rect 11359 2981 11389 3027
rect 11435 2981 11465 3027
rect 11359 2859 11465 2981
rect 11359 2813 11389 2859
rect 11435 2813 11465 2859
rect 11359 2692 11465 2813
rect 11359 2646 11389 2692
rect 11435 2646 11465 2692
rect 11359 2550 11465 2646
rect 11585 2550 11689 3912
rect 11809 2550 11911 3912
rect 12031 3866 12150 3912
rect 12031 3820 12061 3866
rect 12107 3820 12150 3866
rect 12031 3698 12150 3820
rect 12031 3652 12061 3698
rect 12107 3652 12150 3698
rect 12031 3530 12150 3652
rect 12031 3484 12061 3530
rect 12107 3484 12150 3530
rect 12031 3363 12150 3484
rect 12031 3317 12061 3363
rect 12107 3317 12150 3363
rect 12031 3195 12150 3317
rect 12031 3149 12061 3195
rect 12107 3149 12150 3195
rect 12031 3027 12150 3149
rect 12031 2981 12061 3027
rect 12107 2981 12150 3027
rect 12031 2859 12150 2981
rect 12031 2813 12061 2859
rect 12107 2813 12150 2859
rect 12031 2692 12150 2813
rect 12031 2646 12061 2692
rect 12107 2646 12150 2692
rect 12031 2550 12150 2646
rect 12308 3866 12427 3912
rect 12308 3820 12351 3866
rect 12397 3820 12427 3866
rect 12308 3698 12427 3820
rect 12308 3652 12351 3698
rect 12397 3652 12427 3698
rect 12308 3530 12427 3652
rect 12308 3484 12351 3530
rect 12397 3484 12427 3530
rect 12308 3363 12427 3484
rect 12308 3317 12351 3363
rect 12397 3317 12427 3363
rect 12308 3195 12427 3317
rect 12308 3149 12351 3195
rect 12397 3149 12427 3195
rect 12308 3027 12427 3149
rect 12308 2981 12351 3027
rect 12397 2981 12427 3027
rect 12308 2859 12427 2981
rect 12308 2813 12351 2859
rect 12397 2813 12427 2859
rect 12308 2692 12427 2813
rect 12308 2646 12351 2692
rect 12397 2646 12427 2692
rect 12308 2550 12427 2646
rect 12547 2550 12649 3912
rect 12769 2550 12873 3912
rect 12993 3866 13099 3912
rect 12993 3820 13023 3866
rect 13069 3820 13099 3866
rect 12993 3698 13099 3820
rect 12993 3652 13023 3698
rect 13069 3652 13099 3698
rect 12993 3530 13099 3652
rect 12993 3484 13023 3530
rect 13069 3484 13099 3530
rect 12993 3363 13099 3484
rect 12993 3317 13023 3363
rect 13069 3317 13099 3363
rect 12993 3195 13099 3317
rect 12993 3149 13023 3195
rect 13069 3149 13099 3195
rect 12993 3027 13099 3149
rect 12993 2981 13023 3027
rect 13069 2981 13099 3027
rect 12993 2859 13099 2981
rect 12993 2813 13023 2859
rect 13069 2813 13099 2859
rect 12993 2692 13099 2813
rect 12993 2646 13023 2692
rect 13069 2646 13099 2692
rect 12993 2550 13099 2646
rect 13219 2550 13323 3912
rect 13443 2550 13545 3912
rect 13665 3866 13784 3912
rect 13665 3820 13695 3866
rect 13741 3820 13784 3866
rect 13665 3698 13784 3820
rect 13665 3652 13695 3698
rect 13741 3652 13784 3698
rect 13665 3530 13784 3652
rect 13665 3484 13695 3530
rect 13741 3484 13784 3530
rect 13665 3363 13784 3484
rect 13665 3317 13695 3363
rect 13741 3317 13784 3363
rect 13665 3195 13784 3317
rect 13665 3149 13695 3195
rect 13741 3149 13784 3195
rect 13665 3027 13784 3149
rect 13665 2981 13695 3027
rect 13741 2981 13784 3027
rect 13665 2859 13784 2981
rect 13665 2813 13695 2859
rect 13741 2813 13784 2859
rect 13665 2692 13784 2813
rect 13665 2646 13695 2692
rect 13741 2646 13784 2692
rect 13665 2550 13784 2646
rect 9195 1931 9283 1944
rect 9195 1885 9208 1931
rect 9254 1885 9283 1931
rect 7825 1816 7913 1829
rect 7825 1570 7838 1816
rect 7884 1570 7913 1816
rect 7825 1557 7913 1570
rect 8033 1816 8121 1829
rect 8033 1570 8062 1816
rect 8108 1570 8121 1816
rect 9195 1828 9283 1885
rect 8033 1557 8121 1570
rect 9195 1782 9208 1828
rect 9254 1782 9283 1828
rect 9195 1725 9283 1782
rect 9195 1679 9208 1725
rect 9254 1679 9283 1725
rect 9195 1621 9283 1679
rect 9195 1575 9208 1621
rect 9254 1575 9283 1621
rect 9195 1562 9283 1575
rect 9403 1931 9507 1944
rect 9403 1885 9432 1931
rect 9478 1885 9507 1931
rect 9403 1828 9507 1885
rect 9403 1782 9432 1828
rect 9478 1782 9507 1828
rect 9403 1725 9507 1782
rect 9403 1679 9432 1725
rect 9478 1679 9507 1725
rect 9403 1621 9507 1679
rect 9403 1575 9432 1621
rect 9478 1575 9507 1621
rect 9403 1562 9507 1575
rect 9627 1931 9715 1944
rect 9627 1885 9656 1931
rect 9702 1885 9715 1931
rect 9627 1828 9715 1885
rect 9627 1782 9656 1828
rect 9702 1782 9715 1828
rect 9627 1725 9715 1782
rect 9627 1679 9656 1725
rect 9702 1679 9715 1725
rect 9627 1621 9715 1679
rect 9627 1575 9656 1621
rect 9702 1575 9715 1621
rect 9627 1562 9715 1575
<< mvpdiff >>
rect 1646 27452 1734 27465
rect 1646 27406 1659 27452
rect 1705 27406 1734 27452
rect 1646 27347 1734 27406
rect 1646 27301 1659 27347
rect 1705 27301 1734 27347
rect 1646 27242 1734 27301
rect 1646 27196 1659 27242
rect 1705 27196 1734 27242
rect 1646 27137 1734 27196
rect 1646 27091 1659 27137
rect 1705 27091 1734 27137
rect 1646 27032 1734 27091
rect 1646 26986 1659 27032
rect 1705 26986 1734 27032
rect 1646 26927 1734 26986
rect 1646 26881 1659 26927
rect 1705 26881 1734 26927
rect 1646 26822 1734 26881
rect 1646 26776 1659 26822
rect 1705 26776 1734 26822
rect 1646 26717 1734 26776
rect 1646 26671 1659 26717
rect 1705 26671 1734 26717
rect 1646 26612 1734 26671
rect 1646 26566 1659 26612
rect 1705 26566 1734 26612
rect 1646 26507 1734 26566
rect 1646 26461 1659 26507
rect 1705 26461 1734 26507
rect 1646 26402 1734 26461
rect 1646 26356 1659 26402
rect 1705 26356 1734 26402
rect 1646 26297 1734 26356
rect 1646 26251 1659 26297
rect 1705 26251 1734 26297
rect 1646 26192 1734 26251
rect 1646 26146 1659 26192
rect 1705 26146 1734 26192
rect 1646 26088 1734 26146
rect 1646 26042 1659 26088
rect 1705 26042 1734 26088
rect 1646 25984 1734 26042
rect 1646 25938 1659 25984
rect 1705 25938 1734 25984
rect 1646 25880 1734 25938
rect 1646 25834 1659 25880
rect 1705 25834 1734 25880
rect 1646 25776 1734 25834
rect 1646 25730 1659 25776
rect 1705 25730 1734 25776
rect 1646 25672 1734 25730
rect 1646 25626 1659 25672
rect 1705 25626 1734 25672
rect 1646 25568 1734 25626
rect 1646 25522 1659 25568
rect 1705 25522 1734 25568
rect 1646 25464 1734 25522
rect 1646 25418 1659 25464
rect 1705 25418 1734 25464
rect 1646 25360 1734 25418
rect 1646 25314 1659 25360
rect 1705 25314 1734 25360
rect 1646 25256 1734 25314
rect 1646 25210 1659 25256
rect 1705 25210 1734 25256
rect 1646 25197 1734 25210
rect 1854 27452 1958 27465
rect 1854 27406 1883 27452
rect 1929 27406 1958 27452
rect 1854 27347 1958 27406
rect 1854 27301 1883 27347
rect 1929 27301 1958 27347
rect 1854 27242 1958 27301
rect 1854 27196 1883 27242
rect 1929 27196 1958 27242
rect 1854 27137 1958 27196
rect 1854 27091 1883 27137
rect 1929 27091 1958 27137
rect 1854 27032 1958 27091
rect 1854 26986 1883 27032
rect 1929 26986 1958 27032
rect 1854 26927 1958 26986
rect 1854 26881 1883 26927
rect 1929 26881 1958 26927
rect 1854 26822 1958 26881
rect 1854 26776 1883 26822
rect 1929 26776 1958 26822
rect 1854 26717 1958 26776
rect 1854 26671 1883 26717
rect 1929 26671 1958 26717
rect 1854 26612 1958 26671
rect 1854 26566 1883 26612
rect 1929 26566 1958 26612
rect 1854 26507 1958 26566
rect 1854 26461 1883 26507
rect 1929 26461 1958 26507
rect 1854 26402 1958 26461
rect 1854 26356 1883 26402
rect 1929 26356 1958 26402
rect 1854 26297 1958 26356
rect 1854 26251 1883 26297
rect 1929 26251 1958 26297
rect 1854 26192 1958 26251
rect 1854 26146 1883 26192
rect 1929 26146 1958 26192
rect 1854 26088 1958 26146
rect 1854 26042 1883 26088
rect 1929 26042 1958 26088
rect 1854 25984 1958 26042
rect 1854 25938 1883 25984
rect 1929 25938 1958 25984
rect 1854 25880 1958 25938
rect 1854 25834 1883 25880
rect 1929 25834 1958 25880
rect 1854 25776 1958 25834
rect 1854 25730 1883 25776
rect 1929 25730 1958 25776
rect 1854 25672 1958 25730
rect 1854 25626 1883 25672
rect 1929 25626 1958 25672
rect 1854 25568 1958 25626
rect 1854 25522 1883 25568
rect 1929 25522 1958 25568
rect 1854 25464 1958 25522
rect 1854 25418 1883 25464
rect 1929 25418 1958 25464
rect 1854 25360 1958 25418
rect 1854 25314 1883 25360
rect 1929 25314 1958 25360
rect 1854 25256 1958 25314
rect 1854 25210 1883 25256
rect 1929 25210 1958 25256
rect 1854 25197 1958 25210
rect 2078 27452 2182 27465
rect 2078 27406 2107 27452
rect 2153 27406 2182 27452
rect 2078 27347 2182 27406
rect 2078 27301 2107 27347
rect 2153 27301 2182 27347
rect 2078 27242 2182 27301
rect 2078 27196 2107 27242
rect 2153 27196 2182 27242
rect 2078 27137 2182 27196
rect 2078 27091 2107 27137
rect 2153 27091 2182 27137
rect 2078 27032 2182 27091
rect 2078 26986 2107 27032
rect 2153 26986 2182 27032
rect 2078 26927 2182 26986
rect 2078 26881 2107 26927
rect 2153 26881 2182 26927
rect 2078 26822 2182 26881
rect 2078 26776 2107 26822
rect 2153 26776 2182 26822
rect 2078 26717 2182 26776
rect 2078 26671 2107 26717
rect 2153 26671 2182 26717
rect 2078 26612 2182 26671
rect 2078 26566 2107 26612
rect 2153 26566 2182 26612
rect 2078 26507 2182 26566
rect 2078 26461 2107 26507
rect 2153 26461 2182 26507
rect 2078 26402 2182 26461
rect 2078 26356 2107 26402
rect 2153 26356 2182 26402
rect 2078 26297 2182 26356
rect 2078 26251 2107 26297
rect 2153 26251 2182 26297
rect 2078 26192 2182 26251
rect 2078 26146 2107 26192
rect 2153 26146 2182 26192
rect 2078 26088 2182 26146
rect 2078 26042 2107 26088
rect 2153 26042 2182 26088
rect 2078 25984 2182 26042
rect 2078 25938 2107 25984
rect 2153 25938 2182 25984
rect 2078 25880 2182 25938
rect 2078 25834 2107 25880
rect 2153 25834 2182 25880
rect 2078 25776 2182 25834
rect 2078 25730 2107 25776
rect 2153 25730 2182 25776
rect 2078 25672 2182 25730
rect 2078 25626 2107 25672
rect 2153 25626 2182 25672
rect 2078 25568 2182 25626
rect 2078 25522 2107 25568
rect 2153 25522 2182 25568
rect 2078 25464 2182 25522
rect 2078 25418 2107 25464
rect 2153 25418 2182 25464
rect 2078 25360 2182 25418
rect 2078 25314 2107 25360
rect 2153 25314 2182 25360
rect 2078 25256 2182 25314
rect 2078 25210 2107 25256
rect 2153 25210 2182 25256
rect 2078 25197 2182 25210
rect 2302 27452 2406 27465
rect 2302 27406 2331 27452
rect 2377 27406 2406 27452
rect 2302 27347 2406 27406
rect 2302 27301 2331 27347
rect 2377 27301 2406 27347
rect 2302 27242 2406 27301
rect 2302 27196 2331 27242
rect 2377 27196 2406 27242
rect 2302 27137 2406 27196
rect 2302 27091 2331 27137
rect 2377 27091 2406 27137
rect 2302 27032 2406 27091
rect 2302 26986 2331 27032
rect 2377 26986 2406 27032
rect 2302 26927 2406 26986
rect 2302 26881 2331 26927
rect 2377 26881 2406 26927
rect 2302 26822 2406 26881
rect 2302 26776 2331 26822
rect 2377 26776 2406 26822
rect 2302 26717 2406 26776
rect 2302 26671 2331 26717
rect 2377 26671 2406 26717
rect 2302 26612 2406 26671
rect 2302 26566 2331 26612
rect 2377 26566 2406 26612
rect 2302 26507 2406 26566
rect 2302 26461 2331 26507
rect 2377 26461 2406 26507
rect 2302 26402 2406 26461
rect 2302 26356 2331 26402
rect 2377 26356 2406 26402
rect 2302 26297 2406 26356
rect 2302 26251 2331 26297
rect 2377 26251 2406 26297
rect 2302 26192 2406 26251
rect 2302 26146 2331 26192
rect 2377 26146 2406 26192
rect 2302 26088 2406 26146
rect 2302 26042 2331 26088
rect 2377 26042 2406 26088
rect 2302 25984 2406 26042
rect 2302 25938 2331 25984
rect 2377 25938 2406 25984
rect 2302 25880 2406 25938
rect 2302 25834 2331 25880
rect 2377 25834 2406 25880
rect 2302 25776 2406 25834
rect 2302 25730 2331 25776
rect 2377 25730 2406 25776
rect 2302 25672 2406 25730
rect 2302 25626 2331 25672
rect 2377 25626 2406 25672
rect 2302 25568 2406 25626
rect 2302 25522 2331 25568
rect 2377 25522 2406 25568
rect 2302 25464 2406 25522
rect 2302 25418 2331 25464
rect 2377 25418 2406 25464
rect 2302 25360 2406 25418
rect 2302 25314 2331 25360
rect 2377 25314 2406 25360
rect 2302 25256 2406 25314
rect 2302 25210 2331 25256
rect 2377 25210 2406 25256
rect 2302 25197 2406 25210
rect 2526 27452 2630 27465
rect 2526 27406 2555 27452
rect 2601 27406 2630 27452
rect 2526 27347 2630 27406
rect 2526 27301 2555 27347
rect 2601 27301 2630 27347
rect 2526 27242 2630 27301
rect 2526 27196 2555 27242
rect 2601 27196 2630 27242
rect 2526 27137 2630 27196
rect 2526 27091 2555 27137
rect 2601 27091 2630 27137
rect 2526 27032 2630 27091
rect 2526 26986 2555 27032
rect 2601 26986 2630 27032
rect 2526 26927 2630 26986
rect 2526 26881 2555 26927
rect 2601 26881 2630 26927
rect 2526 26822 2630 26881
rect 2526 26776 2555 26822
rect 2601 26776 2630 26822
rect 2526 26717 2630 26776
rect 2526 26671 2555 26717
rect 2601 26671 2630 26717
rect 2526 26612 2630 26671
rect 2526 26566 2555 26612
rect 2601 26566 2630 26612
rect 2526 26507 2630 26566
rect 2526 26461 2555 26507
rect 2601 26461 2630 26507
rect 2526 26402 2630 26461
rect 2526 26356 2555 26402
rect 2601 26356 2630 26402
rect 2526 26297 2630 26356
rect 2526 26251 2555 26297
rect 2601 26251 2630 26297
rect 2526 26192 2630 26251
rect 2526 26146 2555 26192
rect 2601 26146 2630 26192
rect 2526 26088 2630 26146
rect 2526 26042 2555 26088
rect 2601 26042 2630 26088
rect 2526 25984 2630 26042
rect 2526 25938 2555 25984
rect 2601 25938 2630 25984
rect 2526 25880 2630 25938
rect 2526 25834 2555 25880
rect 2601 25834 2630 25880
rect 2526 25776 2630 25834
rect 2526 25730 2555 25776
rect 2601 25730 2630 25776
rect 2526 25672 2630 25730
rect 2526 25626 2555 25672
rect 2601 25626 2630 25672
rect 2526 25568 2630 25626
rect 2526 25522 2555 25568
rect 2601 25522 2630 25568
rect 2526 25464 2630 25522
rect 2526 25418 2555 25464
rect 2601 25418 2630 25464
rect 2526 25360 2630 25418
rect 2526 25314 2555 25360
rect 2601 25314 2630 25360
rect 2526 25256 2630 25314
rect 2526 25210 2555 25256
rect 2601 25210 2630 25256
rect 2526 25197 2630 25210
rect 2750 27452 2854 27465
rect 2750 27406 2779 27452
rect 2825 27406 2854 27452
rect 2750 27347 2854 27406
rect 2750 27301 2779 27347
rect 2825 27301 2854 27347
rect 2750 27242 2854 27301
rect 2750 27196 2779 27242
rect 2825 27196 2854 27242
rect 2750 27137 2854 27196
rect 2750 27091 2779 27137
rect 2825 27091 2854 27137
rect 2750 27032 2854 27091
rect 2750 26986 2779 27032
rect 2825 26986 2854 27032
rect 2750 26927 2854 26986
rect 2750 26881 2779 26927
rect 2825 26881 2854 26927
rect 2750 26822 2854 26881
rect 2750 26776 2779 26822
rect 2825 26776 2854 26822
rect 2750 26717 2854 26776
rect 2750 26671 2779 26717
rect 2825 26671 2854 26717
rect 2750 26612 2854 26671
rect 2750 26566 2779 26612
rect 2825 26566 2854 26612
rect 2750 26507 2854 26566
rect 2750 26461 2779 26507
rect 2825 26461 2854 26507
rect 2750 26402 2854 26461
rect 2750 26356 2779 26402
rect 2825 26356 2854 26402
rect 2750 26297 2854 26356
rect 2750 26251 2779 26297
rect 2825 26251 2854 26297
rect 2750 26192 2854 26251
rect 2750 26146 2779 26192
rect 2825 26146 2854 26192
rect 2750 26088 2854 26146
rect 2750 26042 2779 26088
rect 2825 26042 2854 26088
rect 2750 25984 2854 26042
rect 2750 25938 2779 25984
rect 2825 25938 2854 25984
rect 2750 25880 2854 25938
rect 2750 25834 2779 25880
rect 2825 25834 2854 25880
rect 2750 25776 2854 25834
rect 2750 25730 2779 25776
rect 2825 25730 2854 25776
rect 2750 25672 2854 25730
rect 2750 25626 2779 25672
rect 2825 25626 2854 25672
rect 2750 25568 2854 25626
rect 2750 25522 2779 25568
rect 2825 25522 2854 25568
rect 2750 25464 2854 25522
rect 2750 25418 2779 25464
rect 2825 25418 2854 25464
rect 2750 25360 2854 25418
rect 2750 25314 2779 25360
rect 2825 25314 2854 25360
rect 2750 25256 2854 25314
rect 2750 25210 2779 25256
rect 2825 25210 2854 25256
rect 2750 25197 2854 25210
rect 2974 27452 3078 27465
rect 2974 27406 3003 27452
rect 3049 27406 3078 27452
rect 2974 27347 3078 27406
rect 2974 27301 3003 27347
rect 3049 27301 3078 27347
rect 2974 27242 3078 27301
rect 2974 27196 3003 27242
rect 3049 27196 3078 27242
rect 2974 27137 3078 27196
rect 2974 27091 3003 27137
rect 3049 27091 3078 27137
rect 2974 27032 3078 27091
rect 2974 26986 3003 27032
rect 3049 26986 3078 27032
rect 2974 26927 3078 26986
rect 2974 26881 3003 26927
rect 3049 26881 3078 26927
rect 2974 26822 3078 26881
rect 2974 26776 3003 26822
rect 3049 26776 3078 26822
rect 2974 26717 3078 26776
rect 2974 26671 3003 26717
rect 3049 26671 3078 26717
rect 2974 26612 3078 26671
rect 2974 26566 3003 26612
rect 3049 26566 3078 26612
rect 2974 26507 3078 26566
rect 2974 26461 3003 26507
rect 3049 26461 3078 26507
rect 2974 26402 3078 26461
rect 2974 26356 3003 26402
rect 3049 26356 3078 26402
rect 2974 26297 3078 26356
rect 2974 26251 3003 26297
rect 3049 26251 3078 26297
rect 2974 26192 3078 26251
rect 2974 26146 3003 26192
rect 3049 26146 3078 26192
rect 2974 26088 3078 26146
rect 2974 26042 3003 26088
rect 3049 26042 3078 26088
rect 2974 25984 3078 26042
rect 2974 25938 3003 25984
rect 3049 25938 3078 25984
rect 2974 25880 3078 25938
rect 2974 25834 3003 25880
rect 3049 25834 3078 25880
rect 2974 25776 3078 25834
rect 2974 25730 3003 25776
rect 3049 25730 3078 25776
rect 2974 25672 3078 25730
rect 2974 25626 3003 25672
rect 3049 25626 3078 25672
rect 2974 25568 3078 25626
rect 2974 25522 3003 25568
rect 3049 25522 3078 25568
rect 2974 25464 3078 25522
rect 2974 25418 3003 25464
rect 3049 25418 3078 25464
rect 2974 25360 3078 25418
rect 2974 25314 3003 25360
rect 3049 25314 3078 25360
rect 2974 25256 3078 25314
rect 2974 25210 3003 25256
rect 3049 25210 3078 25256
rect 2974 25197 3078 25210
rect 3198 27452 3302 27465
rect 3198 27406 3227 27452
rect 3273 27406 3302 27452
rect 3198 27347 3302 27406
rect 3198 27301 3227 27347
rect 3273 27301 3302 27347
rect 3198 27242 3302 27301
rect 3198 27196 3227 27242
rect 3273 27196 3302 27242
rect 3198 27137 3302 27196
rect 3198 27091 3227 27137
rect 3273 27091 3302 27137
rect 3198 27032 3302 27091
rect 3198 26986 3227 27032
rect 3273 26986 3302 27032
rect 3198 26927 3302 26986
rect 3198 26881 3227 26927
rect 3273 26881 3302 26927
rect 3198 26822 3302 26881
rect 3198 26776 3227 26822
rect 3273 26776 3302 26822
rect 3198 26717 3302 26776
rect 3198 26671 3227 26717
rect 3273 26671 3302 26717
rect 3198 26612 3302 26671
rect 3198 26566 3227 26612
rect 3273 26566 3302 26612
rect 3198 26507 3302 26566
rect 3198 26461 3227 26507
rect 3273 26461 3302 26507
rect 3198 26402 3302 26461
rect 3198 26356 3227 26402
rect 3273 26356 3302 26402
rect 3198 26297 3302 26356
rect 3198 26251 3227 26297
rect 3273 26251 3302 26297
rect 3198 26192 3302 26251
rect 3198 26146 3227 26192
rect 3273 26146 3302 26192
rect 3198 26088 3302 26146
rect 3198 26042 3227 26088
rect 3273 26042 3302 26088
rect 3198 25984 3302 26042
rect 3198 25938 3227 25984
rect 3273 25938 3302 25984
rect 3198 25880 3302 25938
rect 3198 25834 3227 25880
rect 3273 25834 3302 25880
rect 3198 25776 3302 25834
rect 3198 25730 3227 25776
rect 3273 25730 3302 25776
rect 3198 25672 3302 25730
rect 3198 25626 3227 25672
rect 3273 25626 3302 25672
rect 3198 25568 3302 25626
rect 3198 25522 3227 25568
rect 3273 25522 3302 25568
rect 3198 25464 3302 25522
rect 3198 25418 3227 25464
rect 3273 25418 3302 25464
rect 3198 25360 3302 25418
rect 3198 25314 3227 25360
rect 3273 25314 3302 25360
rect 3198 25256 3302 25314
rect 3198 25210 3227 25256
rect 3273 25210 3302 25256
rect 3198 25197 3302 25210
rect 3422 27452 3526 27465
rect 3422 27406 3451 27452
rect 3497 27406 3526 27452
rect 3422 27347 3526 27406
rect 3422 27301 3451 27347
rect 3497 27301 3526 27347
rect 3422 27242 3526 27301
rect 3422 27196 3451 27242
rect 3497 27196 3526 27242
rect 3422 27137 3526 27196
rect 3422 27091 3451 27137
rect 3497 27091 3526 27137
rect 3422 27032 3526 27091
rect 3422 26986 3451 27032
rect 3497 26986 3526 27032
rect 3422 26927 3526 26986
rect 3422 26881 3451 26927
rect 3497 26881 3526 26927
rect 3422 26822 3526 26881
rect 3422 26776 3451 26822
rect 3497 26776 3526 26822
rect 3422 26717 3526 26776
rect 3422 26671 3451 26717
rect 3497 26671 3526 26717
rect 3422 26612 3526 26671
rect 3422 26566 3451 26612
rect 3497 26566 3526 26612
rect 3422 26507 3526 26566
rect 3422 26461 3451 26507
rect 3497 26461 3526 26507
rect 3422 26402 3526 26461
rect 3422 26356 3451 26402
rect 3497 26356 3526 26402
rect 3422 26297 3526 26356
rect 3422 26251 3451 26297
rect 3497 26251 3526 26297
rect 3422 26192 3526 26251
rect 3422 26146 3451 26192
rect 3497 26146 3526 26192
rect 3422 26088 3526 26146
rect 3422 26042 3451 26088
rect 3497 26042 3526 26088
rect 3422 25984 3526 26042
rect 3422 25938 3451 25984
rect 3497 25938 3526 25984
rect 3422 25880 3526 25938
rect 3422 25834 3451 25880
rect 3497 25834 3526 25880
rect 3422 25776 3526 25834
rect 3422 25730 3451 25776
rect 3497 25730 3526 25776
rect 3422 25672 3526 25730
rect 3422 25626 3451 25672
rect 3497 25626 3526 25672
rect 3422 25568 3526 25626
rect 3422 25522 3451 25568
rect 3497 25522 3526 25568
rect 3422 25464 3526 25522
rect 3422 25418 3451 25464
rect 3497 25418 3526 25464
rect 3422 25360 3526 25418
rect 3422 25314 3451 25360
rect 3497 25314 3526 25360
rect 3422 25256 3526 25314
rect 3422 25210 3451 25256
rect 3497 25210 3526 25256
rect 3422 25197 3526 25210
rect 3646 27452 3750 27465
rect 3646 27406 3675 27452
rect 3721 27406 3750 27452
rect 3646 27347 3750 27406
rect 3646 27301 3675 27347
rect 3721 27301 3750 27347
rect 3646 27242 3750 27301
rect 3646 27196 3675 27242
rect 3721 27196 3750 27242
rect 3646 27137 3750 27196
rect 3646 27091 3675 27137
rect 3721 27091 3750 27137
rect 3646 27032 3750 27091
rect 3646 26986 3675 27032
rect 3721 26986 3750 27032
rect 3646 26927 3750 26986
rect 3646 26881 3675 26927
rect 3721 26881 3750 26927
rect 3646 26822 3750 26881
rect 3646 26776 3675 26822
rect 3721 26776 3750 26822
rect 3646 26717 3750 26776
rect 3646 26671 3675 26717
rect 3721 26671 3750 26717
rect 3646 26612 3750 26671
rect 3646 26566 3675 26612
rect 3721 26566 3750 26612
rect 3646 26507 3750 26566
rect 3646 26461 3675 26507
rect 3721 26461 3750 26507
rect 3646 26402 3750 26461
rect 3646 26356 3675 26402
rect 3721 26356 3750 26402
rect 3646 26297 3750 26356
rect 3646 26251 3675 26297
rect 3721 26251 3750 26297
rect 3646 26192 3750 26251
rect 3646 26146 3675 26192
rect 3721 26146 3750 26192
rect 3646 26088 3750 26146
rect 3646 26042 3675 26088
rect 3721 26042 3750 26088
rect 3646 25984 3750 26042
rect 3646 25938 3675 25984
rect 3721 25938 3750 25984
rect 3646 25880 3750 25938
rect 3646 25834 3675 25880
rect 3721 25834 3750 25880
rect 3646 25776 3750 25834
rect 3646 25730 3675 25776
rect 3721 25730 3750 25776
rect 3646 25672 3750 25730
rect 3646 25626 3675 25672
rect 3721 25626 3750 25672
rect 3646 25568 3750 25626
rect 3646 25522 3675 25568
rect 3721 25522 3750 25568
rect 3646 25464 3750 25522
rect 3646 25418 3675 25464
rect 3721 25418 3750 25464
rect 3646 25360 3750 25418
rect 3646 25314 3675 25360
rect 3721 25314 3750 25360
rect 3646 25256 3750 25314
rect 3646 25210 3675 25256
rect 3721 25210 3750 25256
rect 3646 25197 3750 25210
rect 3870 27452 3974 27465
rect 3870 27406 3899 27452
rect 3945 27406 3974 27452
rect 3870 27347 3974 27406
rect 3870 27301 3899 27347
rect 3945 27301 3974 27347
rect 3870 27242 3974 27301
rect 3870 27196 3899 27242
rect 3945 27196 3974 27242
rect 3870 27137 3974 27196
rect 3870 27091 3899 27137
rect 3945 27091 3974 27137
rect 3870 27032 3974 27091
rect 3870 26986 3899 27032
rect 3945 26986 3974 27032
rect 3870 26927 3974 26986
rect 3870 26881 3899 26927
rect 3945 26881 3974 26927
rect 3870 26822 3974 26881
rect 3870 26776 3899 26822
rect 3945 26776 3974 26822
rect 3870 26717 3974 26776
rect 3870 26671 3899 26717
rect 3945 26671 3974 26717
rect 3870 26612 3974 26671
rect 3870 26566 3899 26612
rect 3945 26566 3974 26612
rect 3870 26507 3974 26566
rect 3870 26461 3899 26507
rect 3945 26461 3974 26507
rect 3870 26402 3974 26461
rect 3870 26356 3899 26402
rect 3945 26356 3974 26402
rect 3870 26297 3974 26356
rect 3870 26251 3899 26297
rect 3945 26251 3974 26297
rect 3870 26192 3974 26251
rect 3870 26146 3899 26192
rect 3945 26146 3974 26192
rect 3870 26088 3974 26146
rect 3870 26042 3899 26088
rect 3945 26042 3974 26088
rect 3870 25984 3974 26042
rect 3870 25938 3899 25984
rect 3945 25938 3974 25984
rect 3870 25880 3974 25938
rect 3870 25834 3899 25880
rect 3945 25834 3974 25880
rect 3870 25776 3974 25834
rect 3870 25730 3899 25776
rect 3945 25730 3974 25776
rect 3870 25672 3974 25730
rect 3870 25626 3899 25672
rect 3945 25626 3974 25672
rect 3870 25568 3974 25626
rect 3870 25522 3899 25568
rect 3945 25522 3974 25568
rect 3870 25464 3974 25522
rect 3870 25418 3899 25464
rect 3945 25418 3974 25464
rect 3870 25360 3974 25418
rect 3870 25314 3899 25360
rect 3945 25314 3974 25360
rect 3870 25256 3974 25314
rect 3870 25210 3899 25256
rect 3945 25210 3974 25256
rect 3870 25197 3974 25210
rect 4094 27452 4198 27465
rect 4094 27406 4123 27452
rect 4169 27406 4198 27452
rect 4094 27347 4198 27406
rect 4094 27301 4123 27347
rect 4169 27301 4198 27347
rect 4094 27242 4198 27301
rect 4094 27196 4123 27242
rect 4169 27196 4198 27242
rect 4094 27137 4198 27196
rect 4094 27091 4123 27137
rect 4169 27091 4198 27137
rect 4094 27032 4198 27091
rect 4094 26986 4123 27032
rect 4169 26986 4198 27032
rect 4094 26927 4198 26986
rect 4094 26881 4123 26927
rect 4169 26881 4198 26927
rect 4094 26822 4198 26881
rect 4094 26776 4123 26822
rect 4169 26776 4198 26822
rect 4094 26717 4198 26776
rect 4094 26671 4123 26717
rect 4169 26671 4198 26717
rect 4094 26612 4198 26671
rect 4094 26566 4123 26612
rect 4169 26566 4198 26612
rect 4094 26507 4198 26566
rect 4094 26461 4123 26507
rect 4169 26461 4198 26507
rect 4094 26402 4198 26461
rect 4094 26356 4123 26402
rect 4169 26356 4198 26402
rect 4094 26297 4198 26356
rect 4094 26251 4123 26297
rect 4169 26251 4198 26297
rect 4094 26192 4198 26251
rect 4094 26146 4123 26192
rect 4169 26146 4198 26192
rect 4094 26088 4198 26146
rect 4094 26042 4123 26088
rect 4169 26042 4198 26088
rect 4094 25984 4198 26042
rect 4094 25938 4123 25984
rect 4169 25938 4198 25984
rect 4094 25880 4198 25938
rect 4094 25834 4123 25880
rect 4169 25834 4198 25880
rect 4094 25776 4198 25834
rect 4094 25730 4123 25776
rect 4169 25730 4198 25776
rect 4094 25672 4198 25730
rect 4094 25626 4123 25672
rect 4169 25626 4198 25672
rect 4094 25568 4198 25626
rect 4094 25522 4123 25568
rect 4169 25522 4198 25568
rect 4094 25464 4198 25522
rect 4094 25418 4123 25464
rect 4169 25418 4198 25464
rect 4094 25360 4198 25418
rect 4094 25314 4123 25360
rect 4169 25314 4198 25360
rect 4094 25256 4198 25314
rect 4094 25210 4123 25256
rect 4169 25210 4198 25256
rect 4094 25197 4198 25210
rect 4318 27452 4422 27465
rect 4318 27406 4347 27452
rect 4393 27406 4422 27452
rect 4318 27347 4422 27406
rect 4318 27301 4347 27347
rect 4393 27301 4422 27347
rect 4318 27242 4422 27301
rect 4318 27196 4347 27242
rect 4393 27196 4422 27242
rect 4318 27137 4422 27196
rect 4318 27091 4347 27137
rect 4393 27091 4422 27137
rect 4318 27032 4422 27091
rect 4318 26986 4347 27032
rect 4393 26986 4422 27032
rect 4318 26927 4422 26986
rect 4318 26881 4347 26927
rect 4393 26881 4422 26927
rect 4318 26822 4422 26881
rect 4318 26776 4347 26822
rect 4393 26776 4422 26822
rect 4318 26717 4422 26776
rect 4318 26671 4347 26717
rect 4393 26671 4422 26717
rect 4318 26612 4422 26671
rect 4318 26566 4347 26612
rect 4393 26566 4422 26612
rect 4318 26507 4422 26566
rect 4318 26461 4347 26507
rect 4393 26461 4422 26507
rect 4318 26402 4422 26461
rect 4318 26356 4347 26402
rect 4393 26356 4422 26402
rect 4318 26297 4422 26356
rect 4318 26251 4347 26297
rect 4393 26251 4422 26297
rect 4318 26192 4422 26251
rect 4318 26146 4347 26192
rect 4393 26146 4422 26192
rect 4318 26088 4422 26146
rect 4318 26042 4347 26088
rect 4393 26042 4422 26088
rect 4318 25984 4422 26042
rect 4318 25938 4347 25984
rect 4393 25938 4422 25984
rect 4318 25880 4422 25938
rect 4318 25834 4347 25880
rect 4393 25834 4422 25880
rect 4318 25776 4422 25834
rect 4318 25730 4347 25776
rect 4393 25730 4422 25776
rect 4318 25672 4422 25730
rect 4318 25626 4347 25672
rect 4393 25626 4422 25672
rect 4318 25568 4422 25626
rect 4318 25522 4347 25568
rect 4393 25522 4422 25568
rect 4318 25464 4422 25522
rect 4318 25418 4347 25464
rect 4393 25418 4422 25464
rect 4318 25360 4422 25418
rect 4318 25314 4347 25360
rect 4393 25314 4422 25360
rect 4318 25256 4422 25314
rect 4318 25210 4347 25256
rect 4393 25210 4422 25256
rect 4318 25197 4422 25210
rect 4542 27452 4646 27465
rect 4542 27406 4571 27452
rect 4617 27406 4646 27452
rect 4542 27347 4646 27406
rect 4542 27301 4571 27347
rect 4617 27301 4646 27347
rect 4542 27242 4646 27301
rect 4542 27196 4571 27242
rect 4617 27196 4646 27242
rect 4542 27137 4646 27196
rect 4542 27091 4571 27137
rect 4617 27091 4646 27137
rect 4542 27032 4646 27091
rect 4542 26986 4571 27032
rect 4617 26986 4646 27032
rect 4542 26927 4646 26986
rect 4542 26881 4571 26927
rect 4617 26881 4646 26927
rect 4542 26822 4646 26881
rect 4542 26776 4571 26822
rect 4617 26776 4646 26822
rect 4542 26717 4646 26776
rect 4542 26671 4571 26717
rect 4617 26671 4646 26717
rect 4542 26612 4646 26671
rect 4542 26566 4571 26612
rect 4617 26566 4646 26612
rect 4542 26507 4646 26566
rect 4542 26461 4571 26507
rect 4617 26461 4646 26507
rect 4542 26402 4646 26461
rect 4542 26356 4571 26402
rect 4617 26356 4646 26402
rect 4542 26297 4646 26356
rect 4542 26251 4571 26297
rect 4617 26251 4646 26297
rect 4542 26192 4646 26251
rect 4542 26146 4571 26192
rect 4617 26146 4646 26192
rect 4542 26088 4646 26146
rect 4542 26042 4571 26088
rect 4617 26042 4646 26088
rect 4542 25984 4646 26042
rect 4542 25938 4571 25984
rect 4617 25938 4646 25984
rect 4542 25880 4646 25938
rect 4542 25834 4571 25880
rect 4617 25834 4646 25880
rect 4542 25776 4646 25834
rect 4542 25730 4571 25776
rect 4617 25730 4646 25776
rect 4542 25672 4646 25730
rect 4542 25626 4571 25672
rect 4617 25626 4646 25672
rect 4542 25568 4646 25626
rect 4542 25522 4571 25568
rect 4617 25522 4646 25568
rect 4542 25464 4646 25522
rect 4542 25418 4571 25464
rect 4617 25418 4646 25464
rect 4542 25360 4646 25418
rect 4542 25314 4571 25360
rect 4617 25314 4646 25360
rect 4542 25256 4646 25314
rect 4542 25210 4571 25256
rect 4617 25210 4646 25256
rect 4542 25197 4646 25210
rect 4766 27452 4870 27465
rect 4766 27406 4795 27452
rect 4841 27406 4870 27452
rect 4766 27347 4870 27406
rect 4766 27301 4795 27347
rect 4841 27301 4870 27347
rect 4766 27242 4870 27301
rect 4766 27196 4795 27242
rect 4841 27196 4870 27242
rect 4766 27137 4870 27196
rect 4766 27091 4795 27137
rect 4841 27091 4870 27137
rect 4766 27032 4870 27091
rect 4766 26986 4795 27032
rect 4841 26986 4870 27032
rect 4766 26927 4870 26986
rect 4766 26881 4795 26927
rect 4841 26881 4870 26927
rect 4766 26822 4870 26881
rect 4766 26776 4795 26822
rect 4841 26776 4870 26822
rect 4766 26717 4870 26776
rect 4766 26671 4795 26717
rect 4841 26671 4870 26717
rect 4766 26612 4870 26671
rect 4766 26566 4795 26612
rect 4841 26566 4870 26612
rect 4766 26507 4870 26566
rect 4766 26461 4795 26507
rect 4841 26461 4870 26507
rect 4766 26402 4870 26461
rect 4766 26356 4795 26402
rect 4841 26356 4870 26402
rect 4766 26297 4870 26356
rect 4766 26251 4795 26297
rect 4841 26251 4870 26297
rect 4766 26192 4870 26251
rect 4766 26146 4795 26192
rect 4841 26146 4870 26192
rect 4766 26088 4870 26146
rect 4766 26042 4795 26088
rect 4841 26042 4870 26088
rect 4766 25984 4870 26042
rect 4766 25938 4795 25984
rect 4841 25938 4870 25984
rect 4766 25880 4870 25938
rect 4766 25834 4795 25880
rect 4841 25834 4870 25880
rect 4766 25776 4870 25834
rect 4766 25730 4795 25776
rect 4841 25730 4870 25776
rect 4766 25672 4870 25730
rect 4766 25626 4795 25672
rect 4841 25626 4870 25672
rect 4766 25568 4870 25626
rect 4766 25522 4795 25568
rect 4841 25522 4870 25568
rect 4766 25464 4870 25522
rect 4766 25418 4795 25464
rect 4841 25418 4870 25464
rect 4766 25360 4870 25418
rect 4766 25314 4795 25360
rect 4841 25314 4870 25360
rect 4766 25256 4870 25314
rect 4766 25210 4795 25256
rect 4841 25210 4870 25256
rect 4766 25197 4870 25210
rect 4990 27452 5094 27465
rect 4990 27406 5019 27452
rect 5065 27406 5094 27452
rect 4990 27347 5094 27406
rect 4990 27301 5019 27347
rect 5065 27301 5094 27347
rect 4990 27242 5094 27301
rect 4990 27196 5019 27242
rect 5065 27196 5094 27242
rect 4990 27137 5094 27196
rect 4990 27091 5019 27137
rect 5065 27091 5094 27137
rect 4990 27032 5094 27091
rect 4990 26986 5019 27032
rect 5065 26986 5094 27032
rect 4990 26927 5094 26986
rect 4990 26881 5019 26927
rect 5065 26881 5094 26927
rect 4990 26822 5094 26881
rect 4990 26776 5019 26822
rect 5065 26776 5094 26822
rect 4990 26717 5094 26776
rect 4990 26671 5019 26717
rect 5065 26671 5094 26717
rect 4990 26612 5094 26671
rect 4990 26566 5019 26612
rect 5065 26566 5094 26612
rect 4990 26507 5094 26566
rect 4990 26461 5019 26507
rect 5065 26461 5094 26507
rect 4990 26402 5094 26461
rect 4990 26356 5019 26402
rect 5065 26356 5094 26402
rect 4990 26297 5094 26356
rect 4990 26251 5019 26297
rect 5065 26251 5094 26297
rect 4990 26192 5094 26251
rect 4990 26146 5019 26192
rect 5065 26146 5094 26192
rect 4990 26088 5094 26146
rect 4990 26042 5019 26088
rect 5065 26042 5094 26088
rect 4990 25984 5094 26042
rect 4990 25938 5019 25984
rect 5065 25938 5094 25984
rect 4990 25880 5094 25938
rect 4990 25834 5019 25880
rect 5065 25834 5094 25880
rect 4990 25776 5094 25834
rect 4990 25730 5019 25776
rect 5065 25730 5094 25776
rect 4990 25672 5094 25730
rect 4990 25626 5019 25672
rect 5065 25626 5094 25672
rect 4990 25568 5094 25626
rect 4990 25522 5019 25568
rect 5065 25522 5094 25568
rect 4990 25464 5094 25522
rect 4990 25418 5019 25464
rect 5065 25418 5094 25464
rect 4990 25360 5094 25418
rect 4990 25314 5019 25360
rect 5065 25314 5094 25360
rect 4990 25256 5094 25314
rect 4990 25210 5019 25256
rect 5065 25210 5094 25256
rect 4990 25197 5094 25210
rect 5214 27452 5302 27465
rect 5214 27406 5243 27452
rect 5289 27406 5302 27452
rect 5214 27347 5302 27406
rect 5214 27301 5243 27347
rect 5289 27301 5302 27347
rect 5214 27242 5302 27301
rect 5214 27196 5243 27242
rect 5289 27196 5302 27242
rect 5214 27137 5302 27196
rect 5214 27091 5243 27137
rect 5289 27091 5302 27137
rect 5889 27382 6008 27427
rect 5889 27336 5933 27382
rect 5979 27336 6008 27382
rect 5889 27178 6008 27336
rect 5889 27132 5933 27178
rect 5979 27132 6008 27178
rect 5214 27032 5302 27091
rect 5889 27086 6008 27132
rect 6128 27086 6231 27427
rect 6351 27382 6456 27427
rect 6351 27336 6381 27382
rect 6427 27336 6456 27382
rect 6351 27178 6456 27336
rect 6351 27132 6381 27178
rect 6427 27132 6456 27178
rect 6351 27086 6456 27132
rect 6576 27086 6679 27427
rect 6799 27382 6918 27427
rect 6799 27336 6829 27382
rect 6875 27336 6918 27382
rect 6799 27178 6918 27336
rect 9025 27452 9113 27465
rect 9025 27406 9038 27452
rect 9084 27406 9113 27452
rect 6799 27132 6829 27178
rect 6875 27132 6918 27178
rect 6799 27086 6918 27132
rect 7396 27315 7484 27328
rect 7396 27269 7409 27315
rect 7455 27269 7484 27315
rect 7396 27159 7484 27269
rect 7396 27113 7409 27159
rect 7455 27113 7484 27159
rect 7396 27100 7484 27113
rect 7604 27315 7708 27328
rect 7604 27269 7633 27315
rect 7679 27269 7708 27315
rect 7604 27159 7708 27269
rect 7604 27113 7633 27159
rect 7679 27113 7708 27159
rect 7604 27100 7708 27113
rect 7828 27315 7916 27328
rect 7828 27269 7857 27315
rect 7903 27269 7916 27315
rect 7828 27159 7916 27269
rect 7828 27113 7857 27159
rect 7903 27113 7916 27159
rect 9025 27347 9113 27406
rect 9025 27301 9038 27347
rect 9084 27301 9113 27347
rect 9025 27242 9113 27301
rect 9025 27196 9038 27242
rect 9084 27196 9113 27242
rect 9025 27137 9113 27196
rect 7828 27100 7916 27113
rect 5214 26986 5243 27032
rect 5289 26986 5302 27032
rect 5214 26927 5302 26986
rect 9025 27091 9038 27137
rect 9084 27091 9113 27137
rect 9025 27032 9113 27091
rect 9025 26986 9038 27032
rect 9084 26986 9113 27032
rect 5214 26881 5243 26927
rect 5289 26881 5302 26927
rect 5214 26822 5302 26881
rect 5214 26776 5243 26822
rect 5289 26776 5302 26822
rect 9025 26927 9113 26986
rect 9025 26881 9038 26927
rect 9084 26881 9113 26927
rect 9025 26822 9113 26881
rect 5214 26717 5302 26776
rect 9025 26776 9038 26822
rect 9084 26776 9113 26822
rect 5214 26671 5243 26717
rect 5289 26671 5302 26717
rect 5214 26612 5302 26671
rect 5214 26566 5243 26612
rect 5289 26566 5302 26612
rect 5214 26507 5302 26566
rect 5214 26461 5243 26507
rect 5289 26461 5302 26507
rect 5214 26402 5302 26461
rect 5214 26356 5243 26402
rect 5289 26356 5302 26402
rect 5214 26297 5302 26356
rect 5214 26251 5243 26297
rect 5289 26251 5302 26297
rect 5214 26192 5302 26251
rect 5214 26146 5243 26192
rect 5289 26146 5302 26192
rect 5214 26088 5302 26146
rect 5214 26042 5243 26088
rect 5289 26042 5302 26088
rect 5214 25984 5302 26042
rect 5214 25938 5243 25984
rect 5289 25938 5302 25984
rect 5214 25880 5302 25938
rect 5214 25834 5243 25880
rect 5289 25834 5302 25880
rect 5214 25776 5302 25834
rect 5214 25730 5243 25776
rect 5289 25730 5302 25776
rect 5214 25672 5302 25730
rect 5214 25626 5243 25672
rect 5289 25626 5302 25672
rect 5214 25568 5302 25626
rect 5214 25522 5243 25568
rect 5289 25522 5302 25568
rect 5214 25464 5302 25522
rect 5214 25418 5243 25464
rect 5289 25418 5302 25464
rect 5214 25360 5302 25418
rect 5214 25314 5243 25360
rect 5289 25314 5302 25360
rect 5214 25256 5302 25314
rect 9025 26717 9113 26776
rect 9025 26671 9038 26717
rect 9084 26671 9113 26717
rect 9025 26612 9113 26671
rect 9025 26566 9038 26612
rect 9084 26566 9113 26612
rect 9025 26507 9113 26566
rect 9025 26461 9038 26507
rect 9084 26461 9113 26507
rect 9025 26402 9113 26461
rect 9025 26356 9038 26402
rect 9084 26356 9113 26402
rect 9025 26297 9113 26356
rect 9025 26251 9038 26297
rect 9084 26251 9113 26297
rect 9025 26192 9113 26251
rect 9025 26146 9038 26192
rect 9084 26146 9113 26192
rect 9025 26088 9113 26146
rect 9025 26042 9038 26088
rect 9084 26042 9113 26088
rect 9025 25984 9113 26042
rect 9025 25938 9038 25984
rect 9084 25938 9113 25984
rect 9025 25880 9113 25938
rect 9025 25834 9038 25880
rect 9084 25834 9113 25880
rect 9025 25776 9113 25834
rect 9025 25730 9038 25776
rect 9084 25730 9113 25776
rect 9025 25672 9113 25730
rect 9025 25626 9038 25672
rect 9084 25626 9113 25672
rect 9025 25568 9113 25626
rect 9025 25522 9038 25568
rect 9084 25522 9113 25568
rect 9025 25464 9113 25522
rect 9025 25418 9038 25464
rect 9084 25418 9113 25464
rect 5214 25210 5243 25256
rect 5289 25210 5302 25256
rect 5214 25197 5302 25210
rect 9025 25360 9113 25418
rect 9025 25314 9038 25360
rect 9084 25314 9113 25360
rect 9025 25256 9113 25314
rect 9025 25210 9038 25256
rect 9084 25210 9113 25256
rect 9025 25197 9113 25210
rect 9233 27452 9337 27465
rect 9233 27406 9262 27452
rect 9308 27406 9337 27452
rect 9233 27347 9337 27406
rect 9233 27301 9262 27347
rect 9308 27301 9337 27347
rect 9233 27242 9337 27301
rect 9233 27196 9262 27242
rect 9308 27196 9337 27242
rect 9233 27137 9337 27196
rect 9233 27091 9262 27137
rect 9308 27091 9337 27137
rect 9233 27032 9337 27091
rect 9233 26986 9262 27032
rect 9308 26986 9337 27032
rect 9233 26927 9337 26986
rect 9233 26881 9262 26927
rect 9308 26881 9337 26927
rect 9233 26822 9337 26881
rect 9233 26776 9262 26822
rect 9308 26776 9337 26822
rect 9233 26717 9337 26776
rect 9233 26671 9262 26717
rect 9308 26671 9337 26717
rect 9233 26612 9337 26671
rect 9233 26566 9262 26612
rect 9308 26566 9337 26612
rect 9233 26507 9337 26566
rect 9233 26461 9262 26507
rect 9308 26461 9337 26507
rect 9233 26402 9337 26461
rect 9233 26356 9262 26402
rect 9308 26356 9337 26402
rect 9233 26297 9337 26356
rect 9233 26251 9262 26297
rect 9308 26251 9337 26297
rect 9233 26192 9337 26251
rect 9233 26146 9262 26192
rect 9308 26146 9337 26192
rect 9233 26088 9337 26146
rect 9233 26042 9262 26088
rect 9308 26042 9337 26088
rect 9233 25984 9337 26042
rect 9233 25938 9262 25984
rect 9308 25938 9337 25984
rect 9233 25880 9337 25938
rect 9233 25834 9262 25880
rect 9308 25834 9337 25880
rect 9233 25776 9337 25834
rect 9233 25730 9262 25776
rect 9308 25730 9337 25776
rect 9233 25672 9337 25730
rect 9233 25626 9262 25672
rect 9308 25626 9337 25672
rect 9233 25568 9337 25626
rect 9233 25522 9262 25568
rect 9308 25522 9337 25568
rect 9233 25464 9337 25522
rect 9233 25418 9262 25464
rect 9308 25418 9337 25464
rect 9233 25360 9337 25418
rect 9233 25314 9262 25360
rect 9308 25314 9337 25360
rect 9233 25256 9337 25314
rect 9233 25210 9262 25256
rect 9308 25210 9337 25256
rect 9233 25197 9337 25210
rect 9457 27452 9561 27465
rect 9457 27406 9486 27452
rect 9532 27406 9561 27452
rect 9457 27347 9561 27406
rect 9457 27301 9486 27347
rect 9532 27301 9561 27347
rect 9457 27242 9561 27301
rect 9457 27196 9486 27242
rect 9532 27196 9561 27242
rect 9457 27137 9561 27196
rect 9457 27091 9486 27137
rect 9532 27091 9561 27137
rect 9457 27032 9561 27091
rect 9457 26986 9486 27032
rect 9532 26986 9561 27032
rect 9457 26927 9561 26986
rect 9457 26881 9486 26927
rect 9532 26881 9561 26927
rect 9457 26822 9561 26881
rect 9457 26776 9486 26822
rect 9532 26776 9561 26822
rect 9457 26717 9561 26776
rect 9457 26671 9486 26717
rect 9532 26671 9561 26717
rect 9457 26612 9561 26671
rect 9457 26566 9486 26612
rect 9532 26566 9561 26612
rect 9457 26507 9561 26566
rect 9457 26461 9486 26507
rect 9532 26461 9561 26507
rect 9457 26402 9561 26461
rect 9457 26356 9486 26402
rect 9532 26356 9561 26402
rect 9457 26297 9561 26356
rect 9457 26251 9486 26297
rect 9532 26251 9561 26297
rect 9457 26192 9561 26251
rect 9457 26146 9486 26192
rect 9532 26146 9561 26192
rect 9457 26088 9561 26146
rect 9457 26042 9486 26088
rect 9532 26042 9561 26088
rect 9457 25984 9561 26042
rect 9457 25938 9486 25984
rect 9532 25938 9561 25984
rect 9457 25880 9561 25938
rect 9457 25834 9486 25880
rect 9532 25834 9561 25880
rect 9457 25776 9561 25834
rect 9457 25730 9486 25776
rect 9532 25730 9561 25776
rect 9457 25672 9561 25730
rect 9457 25626 9486 25672
rect 9532 25626 9561 25672
rect 9457 25568 9561 25626
rect 9457 25522 9486 25568
rect 9532 25522 9561 25568
rect 9457 25464 9561 25522
rect 9457 25418 9486 25464
rect 9532 25418 9561 25464
rect 9457 25360 9561 25418
rect 9457 25314 9486 25360
rect 9532 25314 9561 25360
rect 9457 25256 9561 25314
rect 9457 25210 9486 25256
rect 9532 25210 9561 25256
rect 9457 25197 9561 25210
rect 9681 27452 9785 27465
rect 9681 27406 9710 27452
rect 9756 27406 9785 27452
rect 9681 27347 9785 27406
rect 9681 27301 9710 27347
rect 9756 27301 9785 27347
rect 9681 27242 9785 27301
rect 9681 27196 9710 27242
rect 9756 27196 9785 27242
rect 9681 27137 9785 27196
rect 9681 27091 9710 27137
rect 9756 27091 9785 27137
rect 9681 27032 9785 27091
rect 9681 26986 9710 27032
rect 9756 26986 9785 27032
rect 9681 26927 9785 26986
rect 9681 26881 9710 26927
rect 9756 26881 9785 26927
rect 9681 26822 9785 26881
rect 9681 26776 9710 26822
rect 9756 26776 9785 26822
rect 9681 26717 9785 26776
rect 9681 26671 9710 26717
rect 9756 26671 9785 26717
rect 9681 26612 9785 26671
rect 9681 26566 9710 26612
rect 9756 26566 9785 26612
rect 9681 26507 9785 26566
rect 9681 26461 9710 26507
rect 9756 26461 9785 26507
rect 9681 26402 9785 26461
rect 9681 26356 9710 26402
rect 9756 26356 9785 26402
rect 9681 26297 9785 26356
rect 9681 26251 9710 26297
rect 9756 26251 9785 26297
rect 9681 26192 9785 26251
rect 9681 26146 9710 26192
rect 9756 26146 9785 26192
rect 9681 26088 9785 26146
rect 9681 26042 9710 26088
rect 9756 26042 9785 26088
rect 9681 25984 9785 26042
rect 9681 25938 9710 25984
rect 9756 25938 9785 25984
rect 9681 25880 9785 25938
rect 9681 25834 9710 25880
rect 9756 25834 9785 25880
rect 9681 25776 9785 25834
rect 9681 25730 9710 25776
rect 9756 25730 9785 25776
rect 9681 25672 9785 25730
rect 9681 25626 9710 25672
rect 9756 25626 9785 25672
rect 9681 25568 9785 25626
rect 9681 25522 9710 25568
rect 9756 25522 9785 25568
rect 9681 25464 9785 25522
rect 9681 25418 9710 25464
rect 9756 25418 9785 25464
rect 9681 25360 9785 25418
rect 9681 25314 9710 25360
rect 9756 25314 9785 25360
rect 9681 25256 9785 25314
rect 9681 25210 9710 25256
rect 9756 25210 9785 25256
rect 9681 25197 9785 25210
rect 9905 27452 10009 27465
rect 9905 27406 9934 27452
rect 9980 27406 10009 27452
rect 9905 27347 10009 27406
rect 9905 27301 9934 27347
rect 9980 27301 10009 27347
rect 9905 27242 10009 27301
rect 9905 27196 9934 27242
rect 9980 27196 10009 27242
rect 9905 27137 10009 27196
rect 9905 27091 9934 27137
rect 9980 27091 10009 27137
rect 9905 27032 10009 27091
rect 9905 26986 9934 27032
rect 9980 26986 10009 27032
rect 9905 26927 10009 26986
rect 9905 26881 9934 26927
rect 9980 26881 10009 26927
rect 9905 26822 10009 26881
rect 9905 26776 9934 26822
rect 9980 26776 10009 26822
rect 9905 26717 10009 26776
rect 9905 26671 9934 26717
rect 9980 26671 10009 26717
rect 9905 26612 10009 26671
rect 9905 26566 9934 26612
rect 9980 26566 10009 26612
rect 9905 26507 10009 26566
rect 9905 26461 9934 26507
rect 9980 26461 10009 26507
rect 9905 26402 10009 26461
rect 9905 26356 9934 26402
rect 9980 26356 10009 26402
rect 9905 26297 10009 26356
rect 9905 26251 9934 26297
rect 9980 26251 10009 26297
rect 9905 26192 10009 26251
rect 9905 26146 9934 26192
rect 9980 26146 10009 26192
rect 9905 26088 10009 26146
rect 9905 26042 9934 26088
rect 9980 26042 10009 26088
rect 9905 25984 10009 26042
rect 9905 25938 9934 25984
rect 9980 25938 10009 25984
rect 9905 25880 10009 25938
rect 9905 25834 9934 25880
rect 9980 25834 10009 25880
rect 9905 25776 10009 25834
rect 9905 25730 9934 25776
rect 9980 25730 10009 25776
rect 9905 25672 10009 25730
rect 9905 25626 9934 25672
rect 9980 25626 10009 25672
rect 9905 25568 10009 25626
rect 9905 25522 9934 25568
rect 9980 25522 10009 25568
rect 9905 25464 10009 25522
rect 9905 25418 9934 25464
rect 9980 25418 10009 25464
rect 9905 25360 10009 25418
rect 9905 25314 9934 25360
rect 9980 25314 10009 25360
rect 9905 25256 10009 25314
rect 9905 25210 9934 25256
rect 9980 25210 10009 25256
rect 9905 25197 10009 25210
rect 10129 27452 10233 27465
rect 10129 27406 10158 27452
rect 10204 27406 10233 27452
rect 10129 27347 10233 27406
rect 10129 27301 10158 27347
rect 10204 27301 10233 27347
rect 10129 27242 10233 27301
rect 10129 27196 10158 27242
rect 10204 27196 10233 27242
rect 10129 27137 10233 27196
rect 10129 27091 10158 27137
rect 10204 27091 10233 27137
rect 10129 27032 10233 27091
rect 10129 26986 10158 27032
rect 10204 26986 10233 27032
rect 10129 26927 10233 26986
rect 10129 26881 10158 26927
rect 10204 26881 10233 26927
rect 10129 26822 10233 26881
rect 10129 26776 10158 26822
rect 10204 26776 10233 26822
rect 10129 26717 10233 26776
rect 10129 26671 10158 26717
rect 10204 26671 10233 26717
rect 10129 26612 10233 26671
rect 10129 26566 10158 26612
rect 10204 26566 10233 26612
rect 10129 26507 10233 26566
rect 10129 26461 10158 26507
rect 10204 26461 10233 26507
rect 10129 26402 10233 26461
rect 10129 26356 10158 26402
rect 10204 26356 10233 26402
rect 10129 26297 10233 26356
rect 10129 26251 10158 26297
rect 10204 26251 10233 26297
rect 10129 26192 10233 26251
rect 10129 26146 10158 26192
rect 10204 26146 10233 26192
rect 10129 26088 10233 26146
rect 10129 26042 10158 26088
rect 10204 26042 10233 26088
rect 10129 25984 10233 26042
rect 10129 25938 10158 25984
rect 10204 25938 10233 25984
rect 10129 25880 10233 25938
rect 10129 25834 10158 25880
rect 10204 25834 10233 25880
rect 10129 25776 10233 25834
rect 10129 25730 10158 25776
rect 10204 25730 10233 25776
rect 10129 25672 10233 25730
rect 10129 25626 10158 25672
rect 10204 25626 10233 25672
rect 10129 25568 10233 25626
rect 10129 25522 10158 25568
rect 10204 25522 10233 25568
rect 10129 25464 10233 25522
rect 10129 25418 10158 25464
rect 10204 25418 10233 25464
rect 10129 25360 10233 25418
rect 10129 25314 10158 25360
rect 10204 25314 10233 25360
rect 10129 25256 10233 25314
rect 10129 25210 10158 25256
rect 10204 25210 10233 25256
rect 10129 25197 10233 25210
rect 10353 27452 10457 27465
rect 10353 27406 10382 27452
rect 10428 27406 10457 27452
rect 10353 27347 10457 27406
rect 10353 27301 10382 27347
rect 10428 27301 10457 27347
rect 10353 27242 10457 27301
rect 10353 27196 10382 27242
rect 10428 27196 10457 27242
rect 10353 27137 10457 27196
rect 10353 27091 10382 27137
rect 10428 27091 10457 27137
rect 10353 27032 10457 27091
rect 10353 26986 10382 27032
rect 10428 26986 10457 27032
rect 10353 26927 10457 26986
rect 10353 26881 10382 26927
rect 10428 26881 10457 26927
rect 10353 26822 10457 26881
rect 10353 26776 10382 26822
rect 10428 26776 10457 26822
rect 10353 26717 10457 26776
rect 10353 26671 10382 26717
rect 10428 26671 10457 26717
rect 10353 26612 10457 26671
rect 10353 26566 10382 26612
rect 10428 26566 10457 26612
rect 10353 26507 10457 26566
rect 10353 26461 10382 26507
rect 10428 26461 10457 26507
rect 10353 26402 10457 26461
rect 10353 26356 10382 26402
rect 10428 26356 10457 26402
rect 10353 26297 10457 26356
rect 10353 26251 10382 26297
rect 10428 26251 10457 26297
rect 10353 26192 10457 26251
rect 10353 26146 10382 26192
rect 10428 26146 10457 26192
rect 10353 26088 10457 26146
rect 10353 26042 10382 26088
rect 10428 26042 10457 26088
rect 10353 25984 10457 26042
rect 10353 25938 10382 25984
rect 10428 25938 10457 25984
rect 10353 25880 10457 25938
rect 10353 25834 10382 25880
rect 10428 25834 10457 25880
rect 10353 25776 10457 25834
rect 10353 25730 10382 25776
rect 10428 25730 10457 25776
rect 10353 25672 10457 25730
rect 10353 25626 10382 25672
rect 10428 25626 10457 25672
rect 10353 25568 10457 25626
rect 10353 25522 10382 25568
rect 10428 25522 10457 25568
rect 10353 25464 10457 25522
rect 10353 25418 10382 25464
rect 10428 25418 10457 25464
rect 10353 25360 10457 25418
rect 10353 25314 10382 25360
rect 10428 25314 10457 25360
rect 10353 25256 10457 25314
rect 10353 25210 10382 25256
rect 10428 25210 10457 25256
rect 10353 25197 10457 25210
rect 10577 27452 10681 27465
rect 10577 27406 10606 27452
rect 10652 27406 10681 27452
rect 10577 27347 10681 27406
rect 10577 27301 10606 27347
rect 10652 27301 10681 27347
rect 10577 27242 10681 27301
rect 10577 27196 10606 27242
rect 10652 27196 10681 27242
rect 10577 27137 10681 27196
rect 10577 27091 10606 27137
rect 10652 27091 10681 27137
rect 10577 27032 10681 27091
rect 10577 26986 10606 27032
rect 10652 26986 10681 27032
rect 10577 26927 10681 26986
rect 10577 26881 10606 26927
rect 10652 26881 10681 26927
rect 10577 26822 10681 26881
rect 10577 26776 10606 26822
rect 10652 26776 10681 26822
rect 10577 26717 10681 26776
rect 10577 26671 10606 26717
rect 10652 26671 10681 26717
rect 10577 26612 10681 26671
rect 10577 26566 10606 26612
rect 10652 26566 10681 26612
rect 10577 26507 10681 26566
rect 10577 26461 10606 26507
rect 10652 26461 10681 26507
rect 10577 26402 10681 26461
rect 10577 26356 10606 26402
rect 10652 26356 10681 26402
rect 10577 26297 10681 26356
rect 10577 26251 10606 26297
rect 10652 26251 10681 26297
rect 10577 26192 10681 26251
rect 10577 26146 10606 26192
rect 10652 26146 10681 26192
rect 10577 26088 10681 26146
rect 10577 26042 10606 26088
rect 10652 26042 10681 26088
rect 10577 25984 10681 26042
rect 10577 25938 10606 25984
rect 10652 25938 10681 25984
rect 10577 25880 10681 25938
rect 10577 25834 10606 25880
rect 10652 25834 10681 25880
rect 10577 25776 10681 25834
rect 10577 25730 10606 25776
rect 10652 25730 10681 25776
rect 10577 25672 10681 25730
rect 10577 25626 10606 25672
rect 10652 25626 10681 25672
rect 10577 25568 10681 25626
rect 10577 25522 10606 25568
rect 10652 25522 10681 25568
rect 10577 25464 10681 25522
rect 10577 25418 10606 25464
rect 10652 25418 10681 25464
rect 10577 25360 10681 25418
rect 10577 25314 10606 25360
rect 10652 25314 10681 25360
rect 10577 25256 10681 25314
rect 10577 25210 10606 25256
rect 10652 25210 10681 25256
rect 10577 25197 10681 25210
rect 10801 27452 10905 27465
rect 10801 27406 10830 27452
rect 10876 27406 10905 27452
rect 10801 27347 10905 27406
rect 10801 27301 10830 27347
rect 10876 27301 10905 27347
rect 10801 27242 10905 27301
rect 10801 27196 10830 27242
rect 10876 27196 10905 27242
rect 10801 27137 10905 27196
rect 10801 27091 10830 27137
rect 10876 27091 10905 27137
rect 10801 27032 10905 27091
rect 10801 26986 10830 27032
rect 10876 26986 10905 27032
rect 10801 26927 10905 26986
rect 10801 26881 10830 26927
rect 10876 26881 10905 26927
rect 10801 26822 10905 26881
rect 10801 26776 10830 26822
rect 10876 26776 10905 26822
rect 10801 26717 10905 26776
rect 10801 26671 10830 26717
rect 10876 26671 10905 26717
rect 10801 26612 10905 26671
rect 10801 26566 10830 26612
rect 10876 26566 10905 26612
rect 10801 26507 10905 26566
rect 10801 26461 10830 26507
rect 10876 26461 10905 26507
rect 10801 26402 10905 26461
rect 10801 26356 10830 26402
rect 10876 26356 10905 26402
rect 10801 26297 10905 26356
rect 10801 26251 10830 26297
rect 10876 26251 10905 26297
rect 10801 26192 10905 26251
rect 10801 26146 10830 26192
rect 10876 26146 10905 26192
rect 10801 26088 10905 26146
rect 10801 26042 10830 26088
rect 10876 26042 10905 26088
rect 10801 25984 10905 26042
rect 10801 25938 10830 25984
rect 10876 25938 10905 25984
rect 10801 25880 10905 25938
rect 10801 25834 10830 25880
rect 10876 25834 10905 25880
rect 10801 25776 10905 25834
rect 10801 25730 10830 25776
rect 10876 25730 10905 25776
rect 10801 25672 10905 25730
rect 10801 25626 10830 25672
rect 10876 25626 10905 25672
rect 10801 25568 10905 25626
rect 10801 25522 10830 25568
rect 10876 25522 10905 25568
rect 10801 25464 10905 25522
rect 10801 25418 10830 25464
rect 10876 25418 10905 25464
rect 10801 25360 10905 25418
rect 10801 25314 10830 25360
rect 10876 25314 10905 25360
rect 10801 25256 10905 25314
rect 10801 25210 10830 25256
rect 10876 25210 10905 25256
rect 10801 25197 10905 25210
rect 11025 27452 11129 27465
rect 11025 27406 11054 27452
rect 11100 27406 11129 27452
rect 11025 27347 11129 27406
rect 11025 27301 11054 27347
rect 11100 27301 11129 27347
rect 11025 27242 11129 27301
rect 11025 27196 11054 27242
rect 11100 27196 11129 27242
rect 11025 27137 11129 27196
rect 11025 27091 11054 27137
rect 11100 27091 11129 27137
rect 11025 27032 11129 27091
rect 11025 26986 11054 27032
rect 11100 26986 11129 27032
rect 11025 26927 11129 26986
rect 11025 26881 11054 26927
rect 11100 26881 11129 26927
rect 11025 26822 11129 26881
rect 11025 26776 11054 26822
rect 11100 26776 11129 26822
rect 11025 26717 11129 26776
rect 11025 26671 11054 26717
rect 11100 26671 11129 26717
rect 11025 26612 11129 26671
rect 11025 26566 11054 26612
rect 11100 26566 11129 26612
rect 11025 26507 11129 26566
rect 11025 26461 11054 26507
rect 11100 26461 11129 26507
rect 11025 26402 11129 26461
rect 11025 26356 11054 26402
rect 11100 26356 11129 26402
rect 11025 26297 11129 26356
rect 11025 26251 11054 26297
rect 11100 26251 11129 26297
rect 11025 26192 11129 26251
rect 11025 26146 11054 26192
rect 11100 26146 11129 26192
rect 11025 26088 11129 26146
rect 11025 26042 11054 26088
rect 11100 26042 11129 26088
rect 11025 25984 11129 26042
rect 11025 25938 11054 25984
rect 11100 25938 11129 25984
rect 11025 25880 11129 25938
rect 11025 25834 11054 25880
rect 11100 25834 11129 25880
rect 11025 25776 11129 25834
rect 11025 25730 11054 25776
rect 11100 25730 11129 25776
rect 11025 25672 11129 25730
rect 11025 25626 11054 25672
rect 11100 25626 11129 25672
rect 11025 25568 11129 25626
rect 11025 25522 11054 25568
rect 11100 25522 11129 25568
rect 11025 25464 11129 25522
rect 11025 25418 11054 25464
rect 11100 25418 11129 25464
rect 11025 25360 11129 25418
rect 11025 25314 11054 25360
rect 11100 25314 11129 25360
rect 11025 25256 11129 25314
rect 11025 25210 11054 25256
rect 11100 25210 11129 25256
rect 11025 25197 11129 25210
rect 11249 27452 11353 27465
rect 11249 27406 11278 27452
rect 11324 27406 11353 27452
rect 11249 27347 11353 27406
rect 11249 27301 11278 27347
rect 11324 27301 11353 27347
rect 11249 27242 11353 27301
rect 11249 27196 11278 27242
rect 11324 27196 11353 27242
rect 11249 27137 11353 27196
rect 11249 27091 11278 27137
rect 11324 27091 11353 27137
rect 11249 27032 11353 27091
rect 11249 26986 11278 27032
rect 11324 26986 11353 27032
rect 11249 26927 11353 26986
rect 11249 26881 11278 26927
rect 11324 26881 11353 26927
rect 11249 26822 11353 26881
rect 11249 26776 11278 26822
rect 11324 26776 11353 26822
rect 11249 26717 11353 26776
rect 11249 26671 11278 26717
rect 11324 26671 11353 26717
rect 11249 26612 11353 26671
rect 11249 26566 11278 26612
rect 11324 26566 11353 26612
rect 11249 26507 11353 26566
rect 11249 26461 11278 26507
rect 11324 26461 11353 26507
rect 11249 26402 11353 26461
rect 11249 26356 11278 26402
rect 11324 26356 11353 26402
rect 11249 26297 11353 26356
rect 11249 26251 11278 26297
rect 11324 26251 11353 26297
rect 11249 26192 11353 26251
rect 11249 26146 11278 26192
rect 11324 26146 11353 26192
rect 11249 26088 11353 26146
rect 11249 26042 11278 26088
rect 11324 26042 11353 26088
rect 11249 25984 11353 26042
rect 11249 25938 11278 25984
rect 11324 25938 11353 25984
rect 11249 25880 11353 25938
rect 11249 25834 11278 25880
rect 11324 25834 11353 25880
rect 11249 25776 11353 25834
rect 11249 25730 11278 25776
rect 11324 25730 11353 25776
rect 11249 25672 11353 25730
rect 11249 25626 11278 25672
rect 11324 25626 11353 25672
rect 11249 25568 11353 25626
rect 11249 25522 11278 25568
rect 11324 25522 11353 25568
rect 11249 25464 11353 25522
rect 11249 25418 11278 25464
rect 11324 25418 11353 25464
rect 11249 25360 11353 25418
rect 11249 25314 11278 25360
rect 11324 25314 11353 25360
rect 11249 25256 11353 25314
rect 11249 25210 11278 25256
rect 11324 25210 11353 25256
rect 11249 25197 11353 25210
rect 11473 27452 11577 27465
rect 11473 27406 11502 27452
rect 11548 27406 11577 27452
rect 11473 27347 11577 27406
rect 11473 27301 11502 27347
rect 11548 27301 11577 27347
rect 11473 27242 11577 27301
rect 11473 27196 11502 27242
rect 11548 27196 11577 27242
rect 11473 27137 11577 27196
rect 11473 27091 11502 27137
rect 11548 27091 11577 27137
rect 11473 27032 11577 27091
rect 11473 26986 11502 27032
rect 11548 26986 11577 27032
rect 11473 26927 11577 26986
rect 11473 26881 11502 26927
rect 11548 26881 11577 26927
rect 11473 26822 11577 26881
rect 11473 26776 11502 26822
rect 11548 26776 11577 26822
rect 11473 26717 11577 26776
rect 11473 26671 11502 26717
rect 11548 26671 11577 26717
rect 11473 26612 11577 26671
rect 11473 26566 11502 26612
rect 11548 26566 11577 26612
rect 11473 26507 11577 26566
rect 11473 26461 11502 26507
rect 11548 26461 11577 26507
rect 11473 26402 11577 26461
rect 11473 26356 11502 26402
rect 11548 26356 11577 26402
rect 11473 26297 11577 26356
rect 11473 26251 11502 26297
rect 11548 26251 11577 26297
rect 11473 26192 11577 26251
rect 11473 26146 11502 26192
rect 11548 26146 11577 26192
rect 11473 26088 11577 26146
rect 11473 26042 11502 26088
rect 11548 26042 11577 26088
rect 11473 25984 11577 26042
rect 11473 25938 11502 25984
rect 11548 25938 11577 25984
rect 11473 25880 11577 25938
rect 11473 25834 11502 25880
rect 11548 25834 11577 25880
rect 11473 25776 11577 25834
rect 11473 25730 11502 25776
rect 11548 25730 11577 25776
rect 11473 25672 11577 25730
rect 11473 25626 11502 25672
rect 11548 25626 11577 25672
rect 11473 25568 11577 25626
rect 11473 25522 11502 25568
rect 11548 25522 11577 25568
rect 11473 25464 11577 25522
rect 11473 25418 11502 25464
rect 11548 25418 11577 25464
rect 11473 25360 11577 25418
rect 11473 25314 11502 25360
rect 11548 25314 11577 25360
rect 11473 25256 11577 25314
rect 11473 25210 11502 25256
rect 11548 25210 11577 25256
rect 11473 25197 11577 25210
rect 11697 27452 11801 27465
rect 11697 27406 11726 27452
rect 11772 27406 11801 27452
rect 11697 27347 11801 27406
rect 11697 27301 11726 27347
rect 11772 27301 11801 27347
rect 11697 27242 11801 27301
rect 11697 27196 11726 27242
rect 11772 27196 11801 27242
rect 11697 27137 11801 27196
rect 11697 27091 11726 27137
rect 11772 27091 11801 27137
rect 11697 27032 11801 27091
rect 11697 26986 11726 27032
rect 11772 26986 11801 27032
rect 11697 26927 11801 26986
rect 11697 26881 11726 26927
rect 11772 26881 11801 26927
rect 11697 26822 11801 26881
rect 11697 26776 11726 26822
rect 11772 26776 11801 26822
rect 11697 26717 11801 26776
rect 11697 26671 11726 26717
rect 11772 26671 11801 26717
rect 11697 26612 11801 26671
rect 11697 26566 11726 26612
rect 11772 26566 11801 26612
rect 11697 26507 11801 26566
rect 11697 26461 11726 26507
rect 11772 26461 11801 26507
rect 11697 26402 11801 26461
rect 11697 26356 11726 26402
rect 11772 26356 11801 26402
rect 11697 26297 11801 26356
rect 11697 26251 11726 26297
rect 11772 26251 11801 26297
rect 11697 26192 11801 26251
rect 11697 26146 11726 26192
rect 11772 26146 11801 26192
rect 11697 26088 11801 26146
rect 11697 26042 11726 26088
rect 11772 26042 11801 26088
rect 11697 25984 11801 26042
rect 11697 25938 11726 25984
rect 11772 25938 11801 25984
rect 11697 25880 11801 25938
rect 11697 25834 11726 25880
rect 11772 25834 11801 25880
rect 11697 25776 11801 25834
rect 11697 25730 11726 25776
rect 11772 25730 11801 25776
rect 11697 25672 11801 25730
rect 11697 25626 11726 25672
rect 11772 25626 11801 25672
rect 11697 25568 11801 25626
rect 11697 25522 11726 25568
rect 11772 25522 11801 25568
rect 11697 25464 11801 25522
rect 11697 25418 11726 25464
rect 11772 25418 11801 25464
rect 11697 25360 11801 25418
rect 11697 25314 11726 25360
rect 11772 25314 11801 25360
rect 11697 25256 11801 25314
rect 11697 25210 11726 25256
rect 11772 25210 11801 25256
rect 11697 25197 11801 25210
rect 11921 27452 12025 27465
rect 11921 27406 11950 27452
rect 11996 27406 12025 27452
rect 11921 27347 12025 27406
rect 11921 27301 11950 27347
rect 11996 27301 12025 27347
rect 11921 27242 12025 27301
rect 11921 27196 11950 27242
rect 11996 27196 12025 27242
rect 11921 27137 12025 27196
rect 11921 27091 11950 27137
rect 11996 27091 12025 27137
rect 11921 27032 12025 27091
rect 11921 26986 11950 27032
rect 11996 26986 12025 27032
rect 11921 26927 12025 26986
rect 11921 26881 11950 26927
rect 11996 26881 12025 26927
rect 11921 26822 12025 26881
rect 11921 26776 11950 26822
rect 11996 26776 12025 26822
rect 11921 26717 12025 26776
rect 11921 26671 11950 26717
rect 11996 26671 12025 26717
rect 11921 26612 12025 26671
rect 11921 26566 11950 26612
rect 11996 26566 12025 26612
rect 11921 26507 12025 26566
rect 11921 26461 11950 26507
rect 11996 26461 12025 26507
rect 11921 26402 12025 26461
rect 11921 26356 11950 26402
rect 11996 26356 12025 26402
rect 11921 26297 12025 26356
rect 11921 26251 11950 26297
rect 11996 26251 12025 26297
rect 11921 26192 12025 26251
rect 11921 26146 11950 26192
rect 11996 26146 12025 26192
rect 11921 26088 12025 26146
rect 11921 26042 11950 26088
rect 11996 26042 12025 26088
rect 11921 25984 12025 26042
rect 11921 25938 11950 25984
rect 11996 25938 12025 25984
rect 11921 25880 12025 25938
rect 11921 25834 11950 25880
rect 11996 25834 12025 25880
rect 11921 25776 12025 25834
rect 11921 25730 11950 25776
rect 11996 25730 12025 25776
rect 11921 25672 12025 25730
rect 11921 25626 11950 25672
rect 11996 25626 12025 25672
rect 11921 25568 12025 25626
rect 11921 25522 11950 25568
rect 11996 25522 12025 25568
rect 11921 25464 12025 25522
rect 11921 25418 11950 25464
rect 11996 25418 12025 25464
rect 11921 25360 12025 25418
rect 11921 25314 11950 25360
rect 11996 25314 12025 25360
rect 11921 25256 12025 25314
rect 11921 25210 11950 25256
rect 11996 25210 12025 25256
rect 11921 25197 12025 25210
rect 12145 27452 12249 27465
rect 12145 27406 12174 27452
rect 12220 27406 12249 27452
rect 12145 27347 12249 27406
rect 12145 27301 12174 27347
rect 12220 27301 12249 27347
rect 12145 27242 12249 27301
rect 12145 27196 12174 27242
rect 12220 27196 12249 27242
rect 12145 27137 12249 27196
rect 12145 27091 12174 27137
rect 12220 27091 12249 27137
rect 12145 27032 12249 27091
rect 12145 26986 12174 27032
rect 12220 26986 12249 27032
rect 12145 26927 12249 26986
rect 12145 26881 12174 26927
rect 12220 26881 12249 26927
rect 12145 26822 12249 26881
rect 12145 26776 12174 26822
rect 12220 26776 12249 26822
rect 12145 26717 12249 26776
rect 12145 26671 12174 26717
rect 12220 26671 12249 26717
rect 12145 26612 12249 26671
rect 12145 26566 12174 26612
rect 12220 26566 12249 26612
rect 12145 26507 12249 26566
rect 12145 26461 12174 26507
rect 12220 26461 12249 26507
rect 12145 26402 12249 26461
rect 12145 26356 12174 26402
rect 12220 26356 12249 26402
rect 12145 26297 12249 26356
rect 12145 26251 12174 26297
rect 12220 26251 12249 26297
rect 12145 26192 12249 26251
rect 12145 26146 12174 26192
rect 12220 26146 12249 26192
rect 12145 26088 12249 26146
rect 12145 26042 12174 26088
rect 12220 26042 12249 26088
rect 12145 25984 12249 26042
rect 12145 25938 12174 25984
rect 12220 25938 12249 25984
rect 12145 25880 12249 25938
rect 12145 25834 12174 25880
rect 12220 25834 12249 25880
rect 12145 25776 12249 25834
rect 12145 25730 12174 25776
rect 12220 25730 12249 25776
rect 12145 25672 12249 25730
rect 12145 25626 12174 25672
rect 12220 25626 12249 25672
rect 12145 25568 12249 25626
rect 12145 25522 12174 25568
rect 12220 25522 12249 25568
rect 12145 25464 12249 25522
rect 12145 25418 12174 25464
rect 12220 25418 12249 25464
rect 12145 25360 12249 25418
rect 12145 25314 12174 25360
rect 12220 25314 12249 25360
rect 12145 25256 12249 25314
rect 12145 25210 12174 25256
rect 12220 25210 12249 25256
rect 12145 25197 12249 25210
rect 12369 27452 12473 27465
rect 12369 27406 12398 27452
rect 12444 27406 12473 27452
rect 12369 27347 12473 27406
rect 12369 27301 12398 27347
rect 12444 27301 12473 27347
rect 12369 27242 12473 27301
rect 12369 27196 12398 27242
rect 12444 27196 12473 27242
rect 12369 27137 12473 27196
rect 12369 27091 12398 27137
rect 12444 27091 12473 27137
rect 12369 27032 12473 27091
rect 12369 26986 12398 27032
rect 12444 26986 12473 27032
rect 12369 26927 12473 26986
rect 12369 26881 12398 26927
rect 12444 26881 12473 26927
rect 12369 26822 12473 26881
rect 12369 26776 12398 26822
rect 12444 26776 12473 26822
rect 12369 26717 12473 26776
rect 12369 26671 12398 26717
rect 12444 26671 12473 26717
rect 12369 26612 12473 26671
rect 12369 26566 12398 26612
rect 12444 26566 12473 26612
rect 12369 26507 12473 26566
rect 12369 26461 12398 26507
rect 12444 26461 12473 26507
rect 12369 26402 12473 26461
rect 12369 26356 12398 26402
rect 12444 26356 12473 26402
rect 12369 26297 12473 26356
rect 12369 26251 12398 26297
rect 12444 26251 12473 26297
rect 12369 26192 12473 26251
rect 12369 26146 12398 26192
rect 12444 26146 12473 26192
rect 12369 26088 12473 26146
rect 12369 26042 12398 26088
rect 12444 26042 12473 26088
rect 12369 25984 12473 26042
rect 12369 25938 12398 25984
rect 12444 25938 12473 25984
rect 12369 25880 12473 25938
rect 12369 25834 12398 25880
rect 12444 25834 12473 25880
rect 12369 25776 12473 25834
rect 12369 25730 12398 25776
rect 12444 25730 12473 25776
rect 12369 25672 12473 25730
rect 12369 25626 12398 25672
rect 12444 25626 12473 25672
rect 12369 25568 12473 25626
rect 12369 25522 12398 25568
rect 12444 25522 12473 25568
rect 12369 25464 12473 25522
rect 12369 25418 12398 25464
rect 12444 25418 12473 25464
rect 12369 25360 12473 25418
rect 12369 25314 12398 25360
rect 12444 25314 12473 25360
rect 12369 25256 12473 25314
rect 12369 25210 12398 25256
rect 12444 25210 12473 25256
rect 12369 25197 12473 25210
rect 12593 27452 12681 27465
rect 12593 27406 12622 27452
rect 12668 27406 12681 27452
rect 12593 27347 12681 27406
rect 12593 27301 12622 27347
rect 12668 27301 12681 27347
rect 12593 27242 12681 27301
rect 12593 27196 12622 27242
rect 12668 27196 12681 27242
rect 12593 27137 12681 27196
rect 12593 27091 12622 27137
rect 12668 27091 12681 27137
rect 13268 27382 13387 27427
rect 13268 27336 13312 27382
rect 13358 27336 13387 27382
rect 13268 27178 13387 27336
rect 13268 27132 13312 27178
rect 13358 27132 13387 27178
rect 12593 27032 12681 27091
rect 13268 27086 13387 27132
rect 13507 27086 13610 27427
rect 13730 27382 13835 27427
rect 13730 27336 13760 27382
rect 13806 27336 13835 27382
rect 13730 27178 13835 27336
rect 13730 27132 13760 27178
rect 13806 27132 13835 27178
rect 13730 27086 13835 27132
rect 13955 27086 14058 27427
rect 14178 27382 14297 27427
rect 14178 27336 14208 27382
rect 14254 27336 14297 27382
rect 14178 27178 14297 27336
rect 14178 27132 14208 27178
rect 14254 27132 14297 27178
rect 14178 27086 14297 27132
rect 14775 27315 14863 27328
rect 14775 27269 14788 27315
rect 14834 27269 14863 27315
rect 14775 27159 14863 27269
rect 14775 27113 14788 27159
rect 14834 27113 14863 27159
rect 14775 27100 14863 27113
rect 14983 27315 15087 27328
rect 14983 27269 15012 27315
rect 15058 27269 15087 27315
rect 14983 27159 15087 27269
rect 14983 27113 15012 27159
rect 15058 27113 15087 27159
rect 14983 27100 15087 27113
rect 15207 27315 15295 27328
rect 15207 27269 15236 27315
rect 15282 27269 15295 27315
rect 15207 27159 15295 27269
rect 15207 27113 15236 27159
rect 15282 27113 15295 27159
rect 23753 27382 23872 27541
rect 23753 27336 23797 27382
rect 23843 27336 23872 27382
rect 15207 27100 15295 27113
rect 12593 26986 12622 27032
rect 12668 26986 12681 27032
rect 12593 26927 12681 26986
rect 12593 26881 12622 26927
rect 12668 26881 12681 26927
rect 23753 27178 23872 27336
rect 23753 27132 23797 27178
rect 23843 27132 23872 27178
rect 23753 27086 23872 27132
rect 23992 27086 24096 27541
rect 24216 27382 24320 27541
rect 24216 27336 24245 27382
rect 24291 27336 24320 27382
rect 24216 27178 24320 27336
rect 24216 27132 24245 27178
rect 24291 27132 24320 27178
rect 24216 27086 24320 27132
rect 24440 27086 24544 27541
rect 24664 27382 24783 27541
rect 25260 27429 25348 27442
rect 24664 27336 24693 27382
rect 24739 27336 24783 27382
rect 24664 27178 24783 27336
rect 25260 27383 25273 27429
rect 25319 27383 25348 27429
rect 25260 27294 25348 27383
rect 25260 27248 25273 27294
rect 25319 27248 25348 27294
rect 24664 27132 24693 27178
rect 24739 27132 24783 27178
rect 24664 27086 24783 27132
rect 25260 27159 25348 27248
rect 25260 27113 25273 27159
rect 25319 27113 25348 27159
rect 25260 27100 25348 27113
rect 25468 27429 25572 27442
rect 25468 27383 25497 27429
rect 25543 27383 25572 27429
rect 25468 27294 25572 27383
rect 25468 27248 25497 27294
rect 25543 27248 25572 27294
rect 25468 27159 25572 27248
rect 25468 27113 25497 27159
rect 25543 27113 25572 27159
rect 25468 27100 25572 27113
rect 25692 27429 25780 27442
rect 25692 27383 25721 27429
rect 25767 27383 25780 27429
rect 25692 27294 25780 27383
rect 25692 27248 25721 27294
rect 25767 27248 25780 27294
rect 25692 27159 25780 27248
rect 25692 27113 25721 27159
rect 25767 27113 25780 27159
rect 25692 27100 25780 27113
rect 12593 26822 12681 26881
rect 12593 26776 12622 26822
rect 12668 26776 12681 26822
rect 16691 26888 16779 26901
rect 16691 26842 16704 26888
rect 16750 26842 16779 26888
rect 12593 26717 12681 26776
rect 16691 26783 16779 26842
rect 12593 26671 12622 26717
rect 12668 26671 12681 26717
rect 12593 26612 12681 26671
rect 12593 26566 12622 26612
rect 12668 26566 12681 26612
rect 12593 26507 12681 26566
rect 12593 26461 12622 26507
rect 12668 26461 12681 26507
rect 12593 26402 12681 26461
rect 12593 26356 12622 26402
rect 12668 26356 12681 26402
rect 12593 26297 12681 26356
rect 12593 26251 12622 26297
rect 12668 26251 12681 26297
rect 12593 26192 12681 26251
rect 12593 26146 12622 26192
rect 12668 26146 12681 26192
rect 12593 26088 12681 26146
rect 12593 26042 12622 26088
rect 12668 26042 12681 26088
rect 12593 25984 12681 26042
rect 12593 25938 12622 25984
rect 12668 25938 12681 25984
rect 12593 25880 12681 25938
rect 12593 25834 12622 25880
rect 12668 25834 12681 25880
rect 12593 25776 12681 25834
rect 12593 25730 12622 25776
rect 12668 25730 12681 25776
rect 12593 25672 12681 25730
rect 12593 25626 12622 25672
rect 12668 25626 12681 25672
rect 12593 25568 12681 25626
rect 12593 25522 12622 25568
rect 12668 25522 12681 25568
rect 12593 25464 12681 25522
rect 12593 25418 12622 25464
rect 12668 25418 12681 25464
rect 12593 25360 12681 25418
rect 12593 25314 12622 25360
rect 12668 25314 12681 25360
rect 12593 25256 12681 25314
rect 16691 26737 16704 26783
rect 16750 26737 16779 26783
rect 16691 26678 16779 26737
rect 16691 26632 16704 26678
rect 16750 26632 16779 26678
rect 16691 26573 16779 26632
rect 16691 26527 16704 26573
rect 16750 26527 16779 26573
rect 16691 26468 16779 26527
rect 16691 26422 16704 26468
rect 16750 26422 16779 26468
rect 16691 26363 16779 26422
rect 16691 26317 16704 26363
rect 16750 26317 16779 26363
rect 16691 26258 16779 26317
rect 16691 26212 16704 26258
rect 16750 26212 16779 26258
rect 16691 26153 16779 26212
rect 16691 26107 16704 26153
rect 16750 26107 16779 26153
rect 16691 26048 16779 26107
rect 16691 26002 16704 26048
rect 16750 26002 16779 26048
rect 16691 25943 16779 26002
rect 16691 25897 16704 25943
rect 16750 25897 16779 25943
rect 16691 25838 16779 25897
rect 16691 25792 16704 25838
rect 16750 25792 16779 25838
rect 16691 25733 16779 25792
rect 16691 25687 16704 25733
rect 16750 25687 16779 25733
rect 16691 25628 16779 25687
rect 16691 25582 16704 25628
rect 16750 25582 16779 25628
rect 16691 25524 16779 25582
rect 16691 25478 16704 25524
rect 16750 25478 16779 25524
rect 16691 25420 16779 25478
rect 12593 25210 12622 25256
rect 12668 25210 12681 25256
rect 12593 25197 12681 25210
rect 6078 25002 6166 25015
rect 1804 24550 1892 24563
rect 1804 22566 1817 24550
rect 1863 22566 1892 24550
rect 1804 22509 1892 22566
rect 1804 22463 1817 22509
rect 1863 22463 1892 22509
rect 1804 22406 1892 22463
rect 1804 22360 1817 22406
rect 1863 22360 1892 22406
rect 1804 22303 1892 22360
rect 1804 22257 1817 22303
rect 1863 22257 1892 22303
rect 1804 22200 1892 22257
rect 1804 22154 1817 22200
rect 1863 22154 1892 22200
rect 1804 22097 1892 22154
rect 1804 22051 1817 22097
rect 1863 22051 1892 22097
rect 1804 21994 1892 22051
rect 1804 21948 1817 21994
rect 1863 21948 1892 21994
rect 1804 21891 1892 21948
rect 1804 21845 1817 21891
rect 1863 21845 1892 21891
rect 1804 21788 1892 21845
rect 1804 21742 1817 21788
rect 1863 21742 1892 21788
rect 1804 21685 1892 21742
rect 1804 21639 1817 21685
rect 1863 21639 1892 21685
rect 1804 21582 1892 21639
rect 1804 21536 1817 21582
rect 1863 21536 1892 21582
rect 1804 21523 1892 21536
rect 2012 24550 2116 24563
rect 2012 22566 2041 24550
rect 2087 22566 2116 24550
rect 2012 22509 2116 22566
rect 2012 22463 2041 22509
rect 2087 22463 2116 22509
rect 2012 22406 2116 22463
rect 2012 22360 2041 22406
rect 2087 22360 2116 22406
rect 2012 22303 2116 22360
rect 2012 22257 2041 22303
rect 2087 22257 2116 22303
rect 2012 22200 2116 22257
rect 2012 22154 2041 22200
rect 2087 22154 2116 22200
rect 2012 22097 2116 22154
rect 2012 22051 2041 22097
rect 2087 22051 2116 22097
rect 2012 21994 2116 22051
rect 2012 21948 2041 21994
rect 2087 21948 2116 21994
rect 2012 21891 2116 21948
rect 2012 21845 2041 21891
rect 2087 21845 2116 21891
rect 2012 21788 2116 21845
rect 2012 21742 2041 21788
rect 2087 21742 2116 21788
rect 2012 21685 2116 21742
rect 2012 21639 2041 21685
rect 2087 21639 2116 21685
rect 2012 21582 2116 21639
rect 2012 21536 2041 21582
rect 2087 21536 2116 21582
rect 2012 21523 2116 21536
rect 2236 24550 2324 24563
rect 2236 22566 2265 24550
rect 2311 22566 2324 24550
rect 2236 22509 2324 22566
rect 2236 22463 2265 22509
rect 2311 22463 2324 22509
rect 2236 22406 2324 22463
rect 2236 22360 2265 22406
rect 2311 22360 2324 22406
rect 2236 22303 2324 22360
rect 2236 22257 2265 22303
rect 2311 22257 2324 22303
rect 2236 22200 2324 22257
rect 2236 22154 2265 22200
rect 2311 22154 2324 22200
rect 2236 22097 2324 22154
rect 2236 22051 2265 22097
rect 2311 22051 2324 22097
rect 2236 21994 2324 22051
rect 2832 24550 2920 24563
rect 2832 22566 2845 24550
rect 2891 22566 2920 24550
rect 2832 22509 2920 22566
rect 2832 22463 2845 22509
rect 2891 22463 2920 22509
rect 2832 22406 2920 22463
rect 2832 22360 2845 22406
rect 2891 22360 2920 22406
rect 2832 22303 2920 22360
rect 2832 22257 2845 22303
rect 2891 22257 2920 22303
rect 2832 22200 2920 22257
rect 2832 22154 2845 22200
rect 2891 22154 2920 22200
rect 2832 22097 2920 22154
rect 2832 22051 2845 22097
rect 2891 22051 2920 22097
rect 2236 21948 2265 21994
rect 2311 21948 2324 21994
rect 2236 21891 2324 21948
rect 2236 21845 2265 21891
rect 2311 21845 2324 21891
rect 2236 21788 2324 21845
rect 2236 21742 2265 21788
rect 2311 21742 2324 21788
rect 2236 21685 2324 21742
rect 2236 21639 2265 21685
rect 2311 21639 2324 21685
rect 2832 21994 2920 22051
rect 2832 21948 2845 21994
rect 2891 21948 2920 21994
rect 2832 21891 2920 21948
rect 2832 21845 2845 21891
rect 2891 21845 2920 21891
rect 2832 21788 2920 21845
rect 2832 21742 2845 21788
rect 2891 21742 2920 21788
rect 2832 21685 2920 21742
rect 2236 21582 2324 21639
rect 2236 21536 2265 21582
rect 2311 21536 2324 21582
rect 2236 21523 2324 21536
rect 2832 21639 2845 21685
rect 2891 21639 2920 21685
rect 2832 21582 2920 21639
rect 2832 21536 2845 21582
rect 2891 21536 2920 21582
rect 2832 21523 2920 21536
rect 3040 24550 3144 24563
rect 3040 22566 3069 24550
rect 3115 22566 3144 24550
rect 3040 22509 3144 22566
rect 3040 22463 3069 22509
rect 3115 22463 3144 22509
rect 3040 22406 3144 22463
rect 3040 22360 3069 22406
rect 3115 22360 3144 22406
rect 3040 22303 3144 22360
rect 3040 22257 3069 22303
rect 3115 22257 3144 22303
rect 3040 22200 3144 22257
rect 3040 22154 3069 22200
rect 3115 22154 3144 22200
rect 3040 22097 3144 22154
rect 3040 22051 3069 22097
rect 3115 22051 3144 22097
rect 3040 21994 3144 22051
rect 3040 21948 3069 21994
rect 3115 21948 3144 21994
rect 3040 21891 3144 21948
rect 3040 21845 3069 21891
rect 3115 21845 3144 21891
rect 3040 21788 3144 21845
rect 3040 21742 3069 21788
rect 3115 21742 3144 21788
rect 3040 21685 3144 21742
rect 3040 21639 3069 21685
rect 3115 21639 3144 21685
rect 3040 21582 3144 21639
rect 3040 21536 3069 21582
rect 3115 21536 3144 21582
rect 3040 21523 3144 21536
rect 3264 24550 3352 24563
rect 3264 22566 3293 24550
rect 3339 22566 3352 24550
rect 3264 22509 3352 22566
rect 3264 22463 3293 22509
rect 3339 22463 3352 22509
rect 3264 22406 3352 22463
rect 3264 22360 3293 22406
rect 3339 22360 3352 22406
rect 3264 22303 3352 22360
rect 3264 22257 3293 22303
rect 3339 22257 3352 22303
rect 3264 22200 3352 22257
rect 3264 22154 3293 22200
rect 3339 22154 3352 22200
rect 3264 22097 3352 22154
rect 3264 22051 3293 22097
rect 3339 22051 3352 22097
rect 3264 21994 3352 22051
rect 3264 21948 3293 21994
rect 3339 21948 3352 21994
rect 3264 21891 3352 21948
rect 3264 21845 3293 21891
rect 3339 21845 3352 21891
rect 3264 21788 3352 21845
rect 3264 21742 3293 21788
rect 3339 21742 3352 21788
rect 3264 21685 3352 21742
rect 3264 21639 3293 21685
rect 3339 21639 3352 21685
rect 3264 21582 3352 21639
rect 3264 21536 3293 21582
rect 3339 21536 3352 21582
rect 3264 21523 3352 21536
rect 3596 24550 3684 24563
rect 3596 22566 3609 24550
rect 3655 22566 3684 24550
rect 3596 22509 3684 22566
rect 3596 22463 3609 22509
rect 3655 22463 3684 22509
rect 3596 22406 3684 22463
rect 3596 22360 3609 22406
rect 3655 22360 3684 22406
rect 3596 22303 3684 22360
rect 3596 22257 3609 22303
rect 3655 22257 3684 22303
rect 3596 22200 3684 22257
rect 3596 22154 3609 22200
rect 3655 22154 3684 22200
rect 3596 22097 3684 22154
rect 3596 22051 3609 22097
rect 3655 22051 3684 22097
rect 3596 21994 3684 22051
rect 3596 21948 3609 21994
rect 3655 21948 3684 21994
rect 3596 21891 3684 21948
rect 3596 21845 3609 21891
rect 3655 21845 3684 21891
rect 3596 21788 3684 21845
rect 3596 21742 3609 21788
rect 3655 21742 3684 21788
rect 3596 21685 3684 21742
rect 3596 21639 3609 21685
rect 3655 21639 3684 21685
rect 3596 21582 3684 21639
rect 3596 21536 3609 21582
rect 3655 21536 3684 21582
rect 3596 21523 3684 21536
rect 3804 24550 3908 24563
rect 3804 22566 3833 24550
rect 3879 22566 3908 24550
rect 3804 22509 3908 22566
rect 3804 22463 3833 22509
rect 3879 22463 3908 22509
rect 3804 22406 3908 22463
rect 3804 22360 3833 22406
rect 3879 22360 3908 22406
rect 3804 22303 3908 22360
rect 3804 22257 3833 22303
rect 3879 22257 3908 22303
rect 3804 22200 3908 22257
rect 3804 22154 3833 22200
rect 3879 22154 3908 22200
rect 3804 22097 3908 22154
rect 3804 22051 3833 22097
rect 3879 22051 3908 22097
rect 3804 21994 3908 22051
rect 3804 21948 3833 21994
rect 3879 21948 3908 21994
rect 3804 21891 3908 21948
rect 3804 21845 3833 21891
rect 3879 21845 3908 21891
rect 3804 21788 3908 21845
rect 3804 21742 3833 21788
rect 3879 21742 3908 21788
rect 3804 21685 3908 21742
rect 3804 21639 3833 21685
rect 3879 21639 3908 21685
rect 3804 21582 3908 21639
rect 3804 21536 3833 21582
rect 3879 21536 3908 21582
rect 3804 21523 3908 21536
rect 4028 24550 4116 24563
rect 4028 22566 4057 24550
rect 4103 22566 4116 24550
rect 4028 22509 4116 22566
rect 4028 22463 4057 22509
rect 4103 22463 4116 22509
rect 4028 22406 4116 22463
rect 4028 22360 4057 22406
rect 4103 22360 4116 22406
rect 4028 22303 4116 22360
rect 4028 22257 4057 22303
rect 4103 22257 4116 22303
rect 4028 22200 4116 22257
rect 4028 22154 4057 22200
rect 4103 22154 4116 22200
rect 4028 22097 4116 22154
rect 4028 22051 4057 22097
rect 4103 22051 4116 22097
rect 4028 21994 4116 22051
rect 4624 24550 4712 24563
rect 4624 22566 4637 24550
rect 4683 22566 4712 24550
rect 4624 22509 4712 22566
rect 4624 22463 4637 22509
rect 4683 22463 4712 22509
rect 4624 22406 4712 22463
rect 4624 22360 4637 22406
rect 4683 22360 4712 22406
rect 4624 22303 4712 22360
rect 4624 22257 4637 22303
rect 4683 22257 4712 22303
rect 4624 22200 4712 22257
rect 4624 22154 4637 22200
rect 4683 22154 4712 22200
rect 4624 22097 4712 22154
rect 4624 22051 4637 22097
rect 4683 22051 4712 22097
rect 4028 21948 4057 21994
rect 4103 21948 4116 21994
rect 4028 21891 4116 21948
rect 4028 21845 4057 21891
rect 4103 21845 4116 21891
rect 4028 21788 4116 21845
rect 4028 21742 4057 21788
rect 4103 21742 4116 21788
rect 4028 21685 4116 21742
rect 4028 21639 4057 21685
rect 4103 21639 4116 21685
rect 4624 21994 4712 22051
rect 4624 21948 4637 21994
rect 4683 21948 4712 21994
rect 4624 21891 4712 21948
rect 4624 21845 4637 21891
rect 4683 21845 4712 21891
rect 4624 21788 4712 21845
rect 4624 21742 4637 21788
rect 4683 21742 4712 21788
rect 4624 21685 4712 21742
rect 4028 21582 4116 21639
rect 4028 21536 4057 21582
rect 4103 21536 4116 21582
rect 4028 21523 4116 21536
rect 4624 21639 4637 21685
rect 4683 21639 4712 21685
rect 4624 21582 4712 21639
rect 4624 21536 4637 21582
rect 4683 21536 4712 21582
rect 4624 21523 4712 21536
rect 4832 24550 4936 24563
rect 4832 22566 4861 24550
rect 4907 22566 4936 24550
rect 4832 22509 4936 22566
rect 4832 22463 4861 22509
rect 4907 22463 4936 22509
rect 4832 22406 4936 22463
rect 4832 22360 4861 22406
rect 4907 22360 4936 22406
rect 4832 22303 4936 22360
rect 4832 22257 4861 22303
rect 4907 22257 4936 22303
rect 4832 22200 4936 22257
rect 4832 22154 4861 22200
rect 4907 22154 4936 22200
rect 4832 22097 4936 22154
rect 4832 22051 4861 22097
rect 4907 22051 4936 22097
rect 4832 21994 4936 22051
rect 4832 21948 4861 21994
rect 4907 21948 4936 21994
rect 4832 21891 4936 21948
rect 4832 21845 4861 21891
rect 4907 21845 4936 21891
rect 4832 21788 4936 21845
rect 4832 21742 4861 21788
rect 4907 21742 4936 21788
rect 4832 21685 4936 21742
rect 4832 21639 4861 21685
rect 4907 21639 4936 21685
rect 4832 21582 4936 21639
rect 4832 21536 4861 21582
rect 4907 21536 4936 21582
rect 4832 21523 4936 21536
rect 5056 24550 5144 24563
rect 5056 22566 5085 24550
rect 5131 22566 5144 24550
rect 5056 22509 5144 22566
rect 5056 22463 5085 22509
rect 5131 22463 5144 22509
rect 5056 22406 5144 22463
rect 5056 22360 5085 22406
rect 5131 22360 5144 22406
rect 5056 22303 5144 22360
rect 5056 22257 5085 22303
rect 5131 22257 5144 22303
rect 5056 22200 5144 22257
rect 5056 22154 5085 22200
rect 5131 22154 5144 22200
rect 5056 22097 5144 22154
rect 5056 22051 5085 22097
rect 5131 22051 5144 22097
rect 5056 21994 5144 22051
rect 5056 21948 5085 21994
rect 5131 21948 5144 21994
rect 5056 21891 5144 21948
rect 5056 21845 5085 21891
rect 5131 21845 5144 21891
rect 5056 21788 5144 21845
rect 5056 21742 5085 21788
rect 5131 21742 5144 21788
rect 5056 21685 5144 21742
rect 5056 21639 5085 21685
rect 5131 21639 5144 21685
rect 5056 21582 5144 21639
rect 5056 21536 5085 21582
rect 5131 21536 5144 21582
rect 5056 21523 5144 21536
rect 6078 21490 6091 25002
rect 6137 21490 6166 25002
rect 6078 21477 6166 21490
rect 6286 25002 6374 25015
rect 6286 21490 6315 25002
rect 6361 21490 6374 25002
rect 6592 25003 6680 25016
rect 6592 23427 6605 25003
rect 6651 23427 6680 25003
rect 6592 23370 6680 23427
rect 6592 23324 6605 23370
rect 6651 23324 6680 23370
rect 6592 23267 6680 23324
rect 6592 23221 6605 23267
rect 6651 23221 6680 23267
rect 6592 23164 6680 23221
rect 6592 23118 6605 23164
rect 6651 23118 6680 23164
rect 6592 23061 6680 23118
rect 6592 23015 6605 23061
rect 6651 23015 6680 23061
rect 6592 22958 6680 23015
rect 6592 22912 6605 22958
rect 6651 22912 6680 22958
rect 6592 22855 6680 22912
rect 6592 22809 6605 22855
rect 6651 22809 6680 22855
rect 6592 22752 6680 22809
rect 6592 22706 6605 22752
rect 6651 22706 6680 22752
rect 6592 22649 6680 22706
rect 6592 22603 6605 22649
rect 6651 22603 6680 22649
rect 6592 22546 6680 22603
rect 6592 22500 6605 22546
rect 6651 22500 6680 22546
rect 6592 22443 6680 22500
rect 6592 22397 6605 22443
rect 6651 22397 6680 22443
rect 6592 22384 6680 22397
rect 6800 25003 6888 25016
rect 6800 23427 6829 25003
rect 6875 23427 6888 25003
rect 7769 25002 7857 25015
rect 6800 23370 6888 23427
rect 6800 23324 6829 23370
rect 6875 23324 6888 23370
rect 6800 23267 6888 23324
rect 6800 23221 6829 23267
rect 6875 23221 6888 23267
rect 6800 23164 6888 23221
rect 6800 23118 6829 23164
rect 6875 23118 6888 23164
rect 6800 23061 6888 23118
rect 6800 23015 6829 23061
rect 6875 23015 6888 23061
rect 6800 22958 6888 23015
rect 6800 22912 6829 22958
rect 6875 22912 6888 22958
rect 6800 22855 6888 22912
rect 6800 22809 6829 22855
rect 6875 22809 6888 22855
rect 6800 22752 6888 22809
rect 6800 22706 6829 22752
rect 6875 22706 6888 22752
rect 6800 22649 6888 22706
rect 6800 22603 6829 22649
rect 6875 22603 6888 22649
rect 6800 22546 6888 22603
rect 6800 22500 6829 22546
rect 6875 22500 6888 22546
rect 6800 22443 6888 22500
rect 6800 22397 6829 22443
rect 6875 22397 6888 22443
rect 6800 22384 6888 22397
rect 6286 21477 6374 21490
rect 7769 21490 7782 25002
rect 7828 21490 7857 25002
rect 7769 21477 7857 21490
rect 7977 25002 8065 25015
rect 7977 21490 8006 25002
rect 8052 21490 8065 25002
rect 8283 25003 8371 25016
rect 8283 23427 8296 25003
rect 8342 23427 8371 25003
rect 8283 23370 8371 23427
rect 8283 23324 8296 23370
rect 8342 23324 8371 23370
rect 8283 23267 8371 23324
rect 8283 23221 8296 23267
rect 8342 23221 8371 23267
rect 8283 23164 8371 23221
rect 8283 23118 8296 23164
rect 8342 23118 8371 23164
rect 8283 23061 8371 23118
rect 8283 23015 8296 23061
rect 8342 23015 8371 23061
rect 8283 22958 8371 23015
rect 8283 22912 8296 22958
rect 8342 22912 8371 22958
rect 8283 22855 8371 22912
rect 8283 22809 8296 22855
rect 8342 22809 8371 22855
rect 8283 22752 8371 22809
rect 8283 22706 8296 22752
rect 8342 22706 8371 22752
rect 8283 22649 8371 22706
rect 8283 22603 8296 22649
rect 8342 22603 8371 22649
rect 8283 22546 8371 22603
rect 8283 22500 8296 22546
rect 8342 22500 8371 22546
rect 8283 22443 8371 22500
rect 8283 22397 8296 22443
rect 8342 22397 8371 22443
rect 8283 22384 8371 22397
rect 8491 25003 8579 25016
rect 8491 23427 8520 25003
rect 8566 23427 8579 25003
rect 13457 25002 13545 25015
rect 8491 23370 8579 23427
rect 8491 23324 8520 23370
rect 8566 23324 8579 23370
rect 8491 23267 8579 23324
rect 8491 23221 8520 23267
rect 8566 23221 8579 23267
rect 8491 23164 8579 23221
rect 8491 23118 8520 23164
rect 8566 23118 8579 23164
rect 8491 23061 8579 23118
rect 8491 23015 8520 23061
rect 8566 23015 8579 23061
rect 8491 22958 8579 23015
rect 8491 22912 8520 22958
rect 8566 22912 8579 22958
rect 8491 22855 8579 22912
rect 8491 22809 8520 22855
rect 8566 22809 8579 22855
rect 8491 22752 8579 22809
rect 8491 22706 8520 22752
rect 8566 22706 8579 22752
rect 8491 22649 8579 22706
rect 8491 22603 8520 22649
rect 8566 22603 8579 22649
rect 8491 22546 8579 22603
rect 8491 22500 8520 22546
rect 8566 22500 8579 22546
rect 8491 22443 8579 22500
rect 8491 22397 8520 22443
rect 8566 22397 8579 22443
rect 8491 22384 8579 22397
rect 9183 24550 9271 24563
rect 9183 22566 9196 24550
rect 9242 22566 9271 24550
rect 9183 22509 9271 22566
rect 9183 22463 9196 22509
rect 9242 22463 9271 22509
rect 9183 22406 9271 22463
rect 9183 22360 9196 22406
rect 9242 22360 9271 22406
rect 9183 22303 9271 22360
rect 9183 22257 9196 22303
rect 9242 22257 9271 22303
rect 9183 22200 9271 22257
rect 9183 22154 9196 22200
rect 9242 22154 9271 22200
rect 9183 22097 9271 22154
rect 9183 22051 9196 22097
rect 9242 22051 9271 22097
rect 9183 21994 9271 22051
rect 9183 21948 9196 21994
rect 9242 21948 9271 21994
rect 9183 21891 9271 21948
rect 9183 21845 9196 21891
rect 9242 21845 9271 21891
rect 9183 21788 9271 21845
rect 9183 21742 9196 21788
rect 9242 21742 9271 21788
rect 9183 21685 9271 21742
rect 9183 21639 9196 21685
rect 9242 21639 9271 21685
rect 9183 21582 9271 21639
rect 9183 21536 9196 21582
rect 9242 21536 9271 21582
rect 9183 21523 9271 21536
rect 9391 24550 9495 24563
rect 9391 22566 9420 24550
rect 9466 22566 9495 24550
rect 9391 22509 9495 22566
rect 9391 22463 9420 22509
rect 9466 22463 9495 22509
rect 9391 22406 9495 22463
rect 9391 22360 9420 22406
rect 9466 22360 9495 22406
rect 9391 22303 9495 22360
rect 9391 22257 9420 22303
rect 9466 22257 9495 22303
rect 9391 22200 9495 22257
rect 9391 22154 9420 22200
rect 9466 22154 9495 22200
rect 9391 22097 9495 22154
rect 9391 22051 9420 22097
rect 9466 22051 9495 22097
rect 9391 21994 9495 22051
rect 9391 21948 9420 21994
rect 9466 21948 9495 21994
rect 9391 21891 9495 21948
rect 9391 21845 9420 21891
rect 9466 21845 9495 21891
rect 9391 21788 9495 21845
rect 9391 21742 9420 21788
rect 9466 21742 9495 21788
rect 9391 21685 9495 21742
rect 9391 21639 9420 21685
rect 9466 21639 9495 21685
rect 9391 21582 9495 21639
rect 9391 21536 9420 21582
rect 9466 21536 9495 21582
rect 9391 21523 9495 21536
rect 9615 24550 9703 24563
rect 9615 22566 9644 24550
rect 9690 22566 9703 24550
rect 9615 22509 9703 22566
rect 9615 22463 9644 22509
rect 9690 22463 9703 22509
rect 9615 22406 9703 22463
rect 9615 22360 9644 22406
rect 9690 22360 9703 22406
rect 9615 22303 9703 22360
rect 9615 22257 9644 22303
rect 9690 22257 9703 22303
rect 9615 22200 9703 22257
rect 9615 22154 9644 22200
rect 9690 22154 9703 22200
rect 9615 22097 9703 22154
rect 9615 22051 9644 22097
rect 9690 22051 9703 22097
rect 9615 21994 9703 22051
rect 10211 24550 10299 24563
rect 10211 22566 10224 24550
rect 10270 22566 10299 24550
rect 10211 22509 10299 22566
rect 10211 22463 10224 22509
rect 10270 22463 10299 22509
rect 10211 22406 10299 22463
rect 10211 22360 10224 22406
rect 10270 22360 10299 22406
rect 10211 22303 10299 22360
rect 10211 22257 10224 22303
rect 10270 22257 10299 22303
rect 10211 22200 10299 22257
rect 10211 22154 10224 22200
rect 10270 22154 10299 22200
rect 10211 22097 10299 22154
rect 10211 22051 10224 22097
rect 10270 22051 10299 22097
rect 9615 21948 9644 21994
rect 9690 21948 9703 21994
rect 9615 21891 9703 21948
rect 9615 21845 9644 21891
rect 9690 21845 9703 21891
rect 9615 21788 9703 21845
rect 9615 21742 9644 21788
rect 9690 21742 9703 21788
rect 9615 21685 9703 21742
rect 9615 21639 9644 21685
rect 9690 21639 9703 21685
rect 10211 21994 10299 22051
rect 10211 21948 10224 21994
rect 10270 21948 10299 21994
rect 10211 21891 10299 21948
rect 10211 21845 10224 21891
rect 10270 21845 10299 21891
rect 10211 21788 10299 21845
rect 10211 21742 10224 21788
rect 10270 21742 10299 21788
rect 10211 21685 10299 21742
rect 9615 21582 9703 21639
rect 9615 21536 9644 21582
rect 9690 21536 9703 21582
rect 9615 21523 9703 21536
rect 10211 21639 10224 21685
rect 10270 21639 10299 21685
rect 10211 21582 10299 21639
rect 10211 21536 10224 21582
rect 10270 21536 10299 21582
rect 10211 21523 10299 21536
rect 10419 24550 10523 24563
rect 10419 22566 10448 24550
rect 10494 22566 10523 24550
rect 10419 22509 10523 22566
rect 10419 22463 10448 22509
rect 10494 22463 10523 22509
rect 10419 22406 10523 22463
rect 10419 22360 10448 22406
rect 10494 22360 10523 22406
rect 10419 22303 10523 22360
rect 10419 22257 10448 22303
rect 10494 22257 10523 22303
rect 10419 22200 10523 22257
rect 10419 22154 10448 22200
rect 10494 22154 10523 22200
rect 10419 22097 10523 22154
rect 10419 22051 10448 22097
rect 10494 22051 10523 22097
rect 10419 21994 10523 22051
rect 10419 21948 10448 21994
rect 10494 21948 10523 21994
rect 10419 21891 10523 21948
rect 10419 21845 10448 21891
rect 10494 21845 10523 21891
rect 10419 21788 10523 21845
rect 10419 21742 10448 21788
rect 10494 21742 10523 21788
rect 10419 21685 10523 21742
rect 10419 21639 10448 21685
rect 10494 21639 10523 21685
rect 10419 21582 10523 21639
rect 10419 21536 10448 21582
rect 10494 21536 10523 21582
rect 10419 21523 10523 21536
rect 10643 24550 10731 24563
rect 10643 22566 10672 24550
rect 10718 22566 10731 24550
rect 10643 22509 10731 22566
rect 10643 22463 10672 22509
rect 10718 22463 10731 22509
rect 10643 22406 10731 22463
rect 10643 22360 10672 22406
rect 10718 22360 10731 22406
rect 10643 22303 10731 22360
rect 10643 22257 10672 22303
rect 10718 22257 10731 22303
rect 10643 22200 10731 22257
rect 10643 22154 10672 22200
rect 10718 22154 10731 22200
rect 10643 22097 10731 22154
rect 10643 22051 10672 22097
rect 10718 22051 10731 22097
rect 10643 21994 10731 22051
rect 10643 21948 10672 21994
rect 10718 21948 10731 21994
rect 10643 21891 10731 21948
rect 10643 21845 10672 21891
rect 10718 21845 10731 21891
rect 10643 21788 10731 21845
rect 10643 21742 10672 21788
rect 10718 21742 10731 21788
rect 10643 21685 10731 21742
rect 10643 21639 10672 21685
rect 10718 21639 10731 21685
rect 10643 21582 10731 21639
rect 10643 21536 10672 21582
rect 10718 21536 10731 21582
rect 10643 21523 10731 21536
rect 10975 24550 11063 24563
rect 10975 22566 10988 24550
rect 11034 22566 11063 24550
rect 10975 22509 11063 22566
rect 10975 22463 10988 22509
rect 11034 22463 11063 22509
rect 10975 22406 11063 22463
rect 10975 22360 10988 22406
rect 11034 22360 11063 22406
rect 10975 22303 11063 22360
rect 10975 22257 10988 22303
rect 11034 22257 11063 22303
rect 10975 22200 11063 22257
rect 10975 22154 10988 22200
rect 11034 22154 11063 22200
rect 10975 22097 11063 22154
rect 10975 22051 10988 22097
rect 11034 22051 11063 22097
rect 10975 21994 11063 22051
rect 10975 21948 10988 21994
rect 11034 21948 11063 21994
rect 10975 21891 11063 21948
rect 10975 21845 10988 21891
rect 11034 21845 11063 21891
rect 10975 21788 11063 21845
rect 10975 21742 10988 21788
rect 11034 21742 11063 21788
rect 10975 21685 11063 21742
rect 10975 21639 10988 21685
rect 11034 21639 11063 21685
rect 10975 21582 11063 21639
rect 10975 21536 10988 21582
rect 11034 21536 11063 21582
rect 10975 21523 11063 21536
rect 11183 24550 11287 24563
rect 11183 22566 11212 24550
rect 11258 22566 11287 24550
rect 11183 22509 11287 22566
rect 11183 22463 11212 22509
rect 11258 22463 11287 22509
rect 11183 22406 11287 22463
rect 11183 22360 11212 22406
rect 11258 22360 11287 22406
rect 11183 22303 11287 22360
rect 11183 22257 11212 22303
rect 11258 22257 11287 22303
rect 11183 22200 11287 22257
rect 11183 22154 11212 22200
rect 11258 22154 11287 22200
rect 11183 22097 11287 22154
rect 11183 22051 11212 22097
rect 11258 22051 11287 22097
rect 11183 21994 11287 22051
rect 11183 21948 11212 21994
rect 11258 21948 11287 21994
rect 11183 21891 11287 21948
rect 11183 21845 11212 21891
rect 11258 21845 11287 21891
rect 11183 21788 11287 21845
rect 11183 21742 11212 21788
rect 11258 21742 11287 21788
rect 11183 21685 11287 21742
rect 11183 21639 11212 21685
rect 11258 21639 11287 21685
rect 11183 21582 11287 21639
rect 11183 21536 11212 21582
rect 11258 21536 11287 21582
rect 11183 21523 11287 21536
rect 11407 24550 11495 24563
rect 11407 22566 11436 24550
rect 11482 22566 11495 24550
rect 11407 22509 11495 22566
rect 11407 22463 11436 22509
rect 11482 22463 11495 22509
rect 11407 22406 11495 22463
rect 11407 22360 11436 22406
rect 11482 22360 11495 22406
rect 11407 22303 11495 22360
rect 11407 22257 11436 22303
rect 11482 22257 11495 22303
rect 11407 22200 11495 22257
rect 11407 22154 11436 22200
rect 11482 22154 11495 22200
rect 11407 22097 11495 22154
rect 11407 22051 11436 22097
rect 11482 22051 11495 22097
rect 11407 21994 11495 22051
rect 12003 24550 12091 24563
rect 12003 22566 12016 24550
rect 12062 22566 12091 24550
rect 12003 22509 12091 22566
rect 12003 22463 12016 22509
rect 12062 22463 12091 22509
rect 12003 22406 12091 22463
rect 12003 22360 12016 22406
rect 12062 22360 12091 22406
rect 12003 22303 12091 22360
rect 12003 22257 12016 22303
rect 12062 22257 12091 22303
rect 12003 22200 12091 22257
rect 12003 22154 12016 22200
rect 12062 22154 12091 22200
rect 12003 22097 12091 22154
rect 12003 22051 12016 22097
rect 12062 22051 12091 22097
rect 11407 21948 11436 21994
rect 11482 21948 11495 21994
rect 11407 21891 11495 21948
rect 11407 21845 11436 21891
rect 11482 21845 11495 21891
rect 11407 21788 11495 21845
rect 11407 21742 11436 21788
rect 11482 21742 11495 21788
rect 11407 21685 11495 21742
rect 11407 21639 11436 21685
rect 11482 21639 11495 21685
rect 12003 21994 12091 22051
rect 12003 21948 12016 21994
rect 12062 21948 12091 21994
rect 12003 21891 12091 21948
rect 12003 21845 12016 21891
rect 12062 21845 12091 21891
rect 12003 21788 12091 21845
rect 12003 21742 12016 21788
rect 12062 21742 12091 21788
rect 12003 21685 12091 21742
rect 11407 21582 11495 21639
rect 11407 21536 11436 21582
rect 11482 21536 11495 21582
rect 11407 21523 11495 21536
rect 12003 21639 12016 21685
rect 12062 21639 12091 21685
rect 12003 21582 12091 21639
rect 12003 21536 12016 21582
rect 12062 21536 12091 21582
rect 12003 21523 12091 21536
rect 12211 24550 12315 24563
rect 12211 22566 12240 24550
rect 12286 22566 12315 24550
rect 12211 22509 12315 22566
rect 12211 22463 12240 22509
rect 12286 22463 12315 22509
rect 12211 22406 12315 22463
rect 12211 22360 12240 22406
rect 12286 22360 12315 22406
rect 12211 22303 12315 22360
rect 12211 22257 12240 22303
rect 12286 22257 12315 22303
rect 12211 22200 12315 22257
rect 12211 22154 12240 22200
rect 12286 22154 12315 22200
rect 12211 22097 12315 22154
rect 12211 22051 12240 22097
rect 12286 22051 12315 22097
rect 12211 21994 12315 22051
rect 12211 21948 12240 21994
rect 12286 21948 12315 21994
rect 12211 21891 12315 21948
rect 12211 21845 12240 21891
rect 12286 21845 12315 21891
rect 12211 21788 12315 21845
rect 12211 21742 12240 21788
rect 12286 21742 12315 21788
rect 12211 21685 12315 21742
rect 12211 21639 12240 21685
rect 12286 21639 12315 21685
rect 12211 21582 12315 21639
rect 12211 21536 12240 21582
rect 12286 21536 12315 21582
rect 12211 21523 12315 21536
rect 12435 24550 12523 24563
rect 12435 22566 12464 24550
rect 12510 22566 12523 24550
rect 12435 22509 12523 22566
rect 12435 22463 12464 22509
rect 12510 22463 12523 22509
rect 12435 22406 12523 22463
rect 12435 22360 12464 22406
rect 12510 22360 12523 22406
rect 12435 22303 12523 22360
rect 12435 22257 12464 22303
rect 12510 22257 12523 22303
rect 12435 22200 12523 22257
rect 12435 22154 12464 22200
rect 12510 22154 12523 22200
rect 12435 22097 12523 22154
rect 12435 22051 12464 22097
rect 12510 22051 12523 22097
rect 12435 21994 12523 22051
rect 12435 21948 12464 21994
rect 12510 21948 12523 21994
rect 12435 21891 12523 21948
rect 12435 21845 12464 21891
rect 12510 21845 12523 21891
rect 12435 21788 12523 21845
rect 12435 21742 12464 21788
rect 12510 21742 12523 21788
rect 12435 21685 12523 21742
rect 12435 21639 12464 21685
rect 12510 21639 12523 21685
rect 12435 21582 12523 21639
rect 12435 21536 12464 21582
rect 12510 21536 12523 21582
rect 12435 21523 12523 21536
rect 7977 21477 8065 21490
rect 13457 21490 13470 25002
rect 13516 21490 13545 25002
rect 13457 21477 13545 21490
rect 13665 25002 13753 25015
rect 13665 21490 13694 25002
rect 13740 21490 13753 25002
rect 13971 25003 14059 25016
rect 13971 23427 13984 25003
rect 14030 23427 14059 25003
rect 13971 23370 14059 23427
rect 13971 23324 13984 23370
rect 14030 23324 14059 23370
rect 13971 23267 14059 23324
rect 13971 23221 13984 23267
rect 14030 23221 14059 23267
rect 13971 23164 14059 23221
rect 13971 23118 13984 23164
rect 14030 23118 14059 23164
rect 13971 23061 14059 23118
rect 13971 23015 13984 23061
rect 14030 23015 14059 23061
rect 13971 22958 14059 23015
rect 13971 22912 13984 22958
rect 14030 22912 14059 22958
rect 13971 22855 14059 22912
rect 13971 22809 13984 22855
rect 14030 22809 14059 22855
rect 13971 22752 14059 22809
rect 13971 22706 13984 22752
rect 14030 22706 14059 22752
rect 13971 22649 14059 22706
rect 13971 22603 13984 22649
rect 14030 22603 14059 22649
rect 13971 22546 14059 22603
rect 13971 22500 13984 22546
rect 14030 22500 14059 22546
rect 13971 22443 14059 22500
rect 13971 22397 13984 22443
rect 14030 22397 14059 22443
rect 13971 22384 14059 22397
rect 14179 25003 14267 25016
rect 16691 25374 16704 25420
rect 16750 25374 16779 25420
rect 16691 25316 16779 25374
rect 16691 25270 16704 25316
rect 16750 25270 16779 25316
rect 16691 25212 16779 25270
rect 16691 25166 16704 25212
rect 16750 25166 16779 25212
rect 16691 25108 16779 25166
rect 16691 25062 16704 25108
rect 16750 25062 16779 25108
rect 14179 23427 14208 25003
rect 14254 23427 14267 25003
rect 15148 25002 15236 25015
rect 14179 23370 14267 23427
rect 14179 23324 14208 23370
rect 14254 23324 14267 23370
rect 14179 23267 14267 23324
rect 14179 23221 14208 23267
rect 14254 23221 14267 23267
rect 14179 23164 14267 23221
rect 14179 23118 14208 23164
rect 14254 23118 14267 23164
rect 14179 23061 14267 23118
rect 14179 23015 14208 23061
rect 14254 23015 14267 23061
rect 14179 22958 14267 23015
rect 14179 22912 14208 22958
rect 14254 22912 14267 22958
rect 14179 22855 14267 22912
rect 14179 22809 14208 22855
rect 14254 22809 14267 22855
rect 14179 22752 14267 22809
rect 14179 22706 14208 22752
rect 14254 22706 14267 22752
rect 14179 22649 14267 22706
rect 14179 22603 14208 22649
rect 14254 22603 14267 22649
rect 14179 22546 14267 22603
rect 14179 22500 14208 22546
rect 14254 22500 14267 22546
rect 14179 22443 14267 22500
rect 14179 22397 14208 22443
rect 14254 22397 14267 22443
rect 14179 22384 14267 22397
rect 13665 21477 13753 21490
rect 15148 21490 15161 25002
rect 15207 21490 15236 25002
rect 15148 21477 15236 21490
rect 15356 25002 15444 25015
rect 15356 21490 15385 25002
rect 15431 21490 15444 25002
rect 15662 25003 15750 25016
rect 15662 23427 15675 25003
rect 15721 23427 15750 25003
rect 15662 23370 15750 23427
rect 15662 23324 15675 23370
rect 15721 23324 15750 23370
rect 15662 23267 15750 23324
rect 15662 23221 15675 23267
rect 15721 23221 15750 23267
rect 15662 23164 15750 23221
rect 15662 23118 15675 23164
rect 15721 23118 15750 23164
rect 15662 23061 15750 23118
rect 15662 23015 15675 23061
rect 15721 23015 15750 23061
rect 15662 22958 15750 23015
rect 15662 22912 15675 22958
rect 15721 22912 15750 22958
rect 15662 22855 15750 22912
rect 15662 22809 15675 22855
rect 15721 22809 15750 22855
rect 15662 22752 15750 22809
rect 15662 22706 15675 22752
rect 15721 22706 15750 22752
rect 15662 22649 15750 22706
rect 15662 22603 15675 22649
rect 15721 22603 15750 22649
rect 15662 22546 15750 22603
rect 15662 22500 15675 22546
rect 15721 22500 15750 22546
rect 15662 22443 15750 22500
rect 15662 22397 15675 22443
rect 15721 22397 15750 22443
rect 15662 22384 15750 22397
rect 15870 25003 15958 25016
rect 15870 23427 15899 25003
rect 15945 23427 15958 25003
rect 16691 25004 16779 25062
rect 16691 24958 16704 25004
rect 16750 24958 16779 25004
rect 16691 24900 16779 24958
rect 16691 24854 16704 24900
rect 16750 24854 16779 24900
rect 16691 24796 16779 24854
rect 16691 24750 16704 24796
rect 16750 24750 16779 24796
rect 16691 24692 16779 24750
rect 16691 24646 16704 24692
rect 16750 24646 16779 24692
rect 16691 24633 16779 24646
rect 16899 26888 17003 26901
rect 16899 26842 16928 26888
rect 16974 26842 17003 26888
rect 16899 26783 17003 26842
rect 16899 26737 16928 26783
rect 16974 26737 17003 26783
rect 16899 26678 17003 26737
rect 16899 26632 16928 26678
rect 16974 26632 17003 26678
rect 16899 26573 17003 26632
rect 16899 26527 16928 26573
rect 16974 26527 17003 26573
rect 16899 26468 17003 26527
rect 16899 26422 16928 26468
rect 16974 26422 17003 26468
rect 16899 26363 17003 26422
rect 16899 26317 16928 26363
rect 16974 26317 17003 26363
rect 16899 26258 17003 26317
rect 16899 26212 16928 26258
rect 16974 26212 17003 26258
rect 16899 26153 17003 26212
rect 16899 26107 16928 26153
rect 16974 26107 17003 26153
rect 16899 26048 17003 26107
rect 16899 26002 16928 26048
rect 16974 26002 17003 26048
rect 16899 25943 17003 26002
rect 16899 25897 16928 25943
rect 16974 25897 17003 25943
rect 16899 25838 17003 25897
rect 16899 25792 16928 25838
rect 16974 25792 17003 25838
rect 16899 25733 17003 25792
rect 16899 25687 16928 25733
rect 16974 25687 17003 25733
rect 16899 25628 17003 25687
rect 16899 25582 16928 25628
rect 16974 25582 17003 25628
rect 16899 25524 17003 25582
rect 16899 25478 16928 25524
rect 16974 25478 17003 25524
rect 16899 25420 17003 25478
rect 16899 25374 16928 25420
rect 16974 25374 17003 25420
rect 16899 25316 17003 25374
rect 16899 25270 16928 25316
rect 16974 25270 17003 25316
rect 16899 25212 17003 25270
rect 16899 25166 16928 25212
rect 16974 25166 17003 25212
rect 16899 25108 17003 25166
rect 16899 25062 16928 25108
rect 16974 25062 17003 25108
rect 16899 25004 17003 25062
rect 16899 24958 16928 25004
rect 16974 24958 17003 25004
rect 16899 24900 17003 24958
rect 16899 24854 16928 24900
rect 16974 24854 17003 24900
rect 16899 24796 17003 24854
rect 16899 24750 16928 24796
rect 16974 24750 17003 24796
rect 16899 24692 17003 24750
rect 16899 24646 16928 24692
rect 16974 24646 17003 24692
rect 16899 24633 17003 24646
rect 17123 26888 17227 26901
rect 17123 26842 17152 26888
rect 17198 26842 17227 26888
rect 17123 26783 17227 26842
rect 17123 26737 17152 26783
rect 17198 26737 17227 26783
rect 17123 26678 17227 26737
rect 17123 26632 17152 26678
rect 17198 26632 17227 26678
rect 17123 26573 17227 26632
rect 17123 26527 17152 26573
rect 17198 26527 17227 26573
rect 17123 26468 17227 26527
rect 17123 26422 17152 26468
rect 17198 26422 17227 26468
rect 17123 26363 17227 26422
rect 17123 26317 17152 26363
rect 17198 26317 17227 26363
rect 17123 26258 17227 26317
rect 17123 26212 17152 26258
rect 17198 26212 17227 26258
rect 17123 26153 17227 26212
rect 17123 26107 17152 26153
rect 17198 26107 17227 26153
rect 17123 26048 17227 26107
rect 17123 26002 17152 26048
rect 17198 26002 17227 26048
rect 17123 25943 17227 26002
rect 17123 25897 17152 25943
rect 17198 25897 17227 25943
rect 17123 25838 17227 25897
rect 17123 25792 17152 25838
rect 17198 25792 17227 25838
rect 17123 25733 17227 25792
rect 17123 25687 17152 25733
rect 17198 25687 17227 25733
rect 17123 25628 17227 25687
rect 17123 25582 17152 25628
rect 17198 25582 17227 25628
rect 17123 25524 17227 25582
rect 17123 25478 17152 25524
rect 17198 25478 17227 25524
rect 17123 25420 17227 25478
rect 17123 25374 17152 25420
rect 17198 25374 17227 25420
rect 17123 25316 17227 25374
rect 17123 25270 17152 25316
rect 17198 25270 17227 25316
rect 17123 25212 17227 25270
rect 17123 25166 17152 25212
rect 17198 25166 17227 25212
rect 17123 25108 17227 25166
rect 17123 25062 17152 25108
rect 17198 25062 17227 25108
rect 17123 25004 17227 25062
rect 17123 24958 17152 25004
rect 17198 24958 17227 25004
rect 17123 24900 17227 24958
rect 17123 24854 17152 24900
rect 17198 24854 17227 24900
rect 17123 24796 17227 24854
rect 17123 24750 17152 24796
rect 17198 24750 17227 24796
rect 17123 24692 17227 24750
rect 17123 24646 17152 24692
rect 17198 24646 17227 24692
rect 17123 24633 17227 24646
rect 17347 26888 17451 26901
rect 17347 26842 17376 26888
rect 17422 26842 17451 26888
rect 17347 26783 17451 26842
rect 17347 26737 17376 26783
rect 17422 26737 17451 26783
rect 17347 26678 17451 26737
rect 17347 26632 17376 26678
rect 17422 26632 17451 26678
rect 17347 26573 17451 26632
rect 17347 26527 17376 26573
rect 17422 26527 17451 26573
rect 17347 26468 17451 26527
rect 17347 26422 17376 26468
rect 17422 26422 17451 26468
rect 17347 26363 17451 26422
rect 17347 26317 17376 26363
rect 17422 26317 17451 26363
rect 17347 26258 17451 26317
rect 17347 26212 17376 26258
rect 17422 26212 17451 26258
rect 17347 26153 17451 26212
rect 17347 26107 17376 26153
rect 17422 26107 17451 26153
rect 17347 26048 17451 26107
rect 17347 26002 17376 26048
rect 17422 26002 17451 26048
rect 17347 25943 17451 26002
rect 17347 25897 17376 25943
rect 17422 25897 17451 25943
rect 17347 25838 17451 25897
rect 17347 25792 17376 25838
rect 17422 25792 17451 25838
rect 17347 25733 17451 25792
rect 17347 25687 17376 25733
rect 17422 25687 17451 25733
rect 17347 25628 17451 25687
rect 17347 25582 17376 25628
rect 17422 25582 17451 25628
rect 17347 25524 17451 25582
rect 17347 25478 17376 25524
rect 17422 25478 17451 25524
rect 17347 25420 17451 25478
rect 17347 25374 17376 25420
rect 17422 25374 17451 25420
rect 17347 25316 17451 25374
rect 17347 25270 17376 25316
rect 17422 25270 17451 25316
rect 17347 25212 17451 25270
rect 17347 25166 17376 25212
rect 17422 25166 17451 25212
rect 17347 25108 17451 25166
rect 17347 25062 17376 25108
rect 17422 25062 17451 25108
rect 17347 25004 17451 25062
rect 17347 24958 17376 25004
rect 17422 24958 17451 25004
rect 17347 24900 17451 24958
rect 17347 24854 17376 24900
rect 17422 24854 17451 24900
rect 17347 24796 17451 24854
rect 17347 24750 17376 24796
rect 17422 24750 17451 24796
rect 17347 24692 17451 24750
rect 17347 24646 17376 24692
rect 17422 24646 17451 24692
rect 17347 24633 17451 24646
rect 17571 26888 17675 26901
rect 17571 26842 17600 26888
rect 17646 26842 17675 26888
rect 17571 26783 17675 26842
rect 17571 26737 17600 26783
rect 17646 26737 17675 26783
rect 17571 26678 17675 26737
rect 17571 26632 17600 26678
rect 17646 26632 17675 26678
rect 17571 26573 17675 26632
rect 17571 26527 17600 26573
rect 17646 26527 17675 26573
rect 17571 26468 17675 26527
rect 17571 26422 17600 26468
rect 17646 26422 17675 26468
rect 17571 26363 17675 26422
rect 17571 26317 17600 26363
rect 17646 26317 17675 26363
rect 17571 26258 17675 26317
rect 17571 26212 17600 26258
rect 17646 26212 17675 26258
rect 17571 26153 17675 26212
rect 17571 26107 17600 26153
rect 17646 26107 17675 26153
rect 17571 26048 17675 26107
rect 17571 26002 17600 26048
rect 17646 26002 17675 26048
rect 17571 25943 17675 26002
rect 17571 25897 17600 25943
rect 17646 25897 17675 25943
rect 17571 25838 17675 25897
rect 17571 25792 17600 25838
rect 17646 25792 17675 25838
rect 17571 25733 17675 25792
rect 17571 25687 17600 25733
rect 17646 25687 17675 25733
rect 17571 25628 17675 25687
rect 17571 25582 17600 25628
rect 17646 25582 17675 25628
rect 17571 25524 17675 25582
rect 17571 25478 17600 25524
rect 17646 25478 17675 25524
rect 17571 25420 17675 25478
rect 17571 25374 17600 25420
rect 17646 25374 17675 25420
rect 17571 25316 17675 25374
rect 17571 25270 17600 25316
rect 17646 25270 17675 25316
rect 17571 25212 17675 25270
rect 17571 25166 17600 25212
rect 17646 25166 17675 25212
rect 17571 25108 17675 25166
rect 17571 25062 17600 25108
rect 17646 25062 17675 25108
rect 17571 25004 17675 25062
rect 17571 24958 17600 25004
rect 17646 24958 17675 25004
rect 17571 24900 17675 24958
rect 17571 24854 17600 24900
rect 17646 24854 17675 24900
rect 17571 24796 17675 24854
rect 17571 24750 17600 24796
rect 17646 24750 17675 24796
rect 17571 24692 17675 24750
rect 17571 24646 17600 24692
rect 17646 24646 17675 24692
rect 17571 24633 17675 24646
rect 17795 26888 17899 26901
rect 17795 26842 17824 26888
rect 17870 26842 17899 26888
rect 17795 26783 17899 26842
rect 17795 26737 17824 26783
rect 17870 26737 17899 26783
rect 17795 26678 17899 26737
rect 17795 26632 17824 26678
rect 17870 26632 17899 26678
rect 17795 26573 17899 26632
rect 17795 26527 17824 26573
rect 17870 26527 17899 26573
rect 17795 26468 17899 26527
rect 17795 26422 17824 26468
rect 17870 26422 17899 26468
rect 17795 26363 17899 26422
rect 17795 26317 17824 26363
rect 17870 26317 17899 26363
rect 17795 26258 17899 26317
rect 17795 26212 17824 26258
rect 17870 26212 17899 26258
rect 17795 26153 17899 26212
rect 17795 26107 17824 26153
rect 17870 26107 17899 26153
rect 17795 26048 17899 26107
rect 17795 26002 17824 26048
rect 17870 26002 17899 26048
rect 17795 25943 17899 26002
rect 17795 25897 17824 25943
rect 17870 25897 17899 25943
rect 17795 25838 17899 25897
rect 17795 25792 17824 25838
rect 17870 25792 17899 25838
rect 17795 25733 17899 25792
rect 17795 25687 17824 25733
rect 17870 25687 17899 25733
rect 17795 25628 17899 25687
rect 17795 25582 17824 25628
rect 17870 25582 17899 25628
rect 17795 25524 17899 25582
rect 17795 25478 17824 25524
rect 17870 25478 17899 25524
rect 17795 25420 17899 25478
rect 17795 25374 17824 25420
rect 17870 25374 17899 25420
rect 17795 25316 17899 25374
rect 17795 25270 17824 25316
rect 17870 25270 17899 25316
rect 17795 25212 17899 25270
rect 17795 25166 17824 25212
rect 17870 25166 17899 25212
rect 17795 25108 17899 25166
rect 17795 25062 17824 25108
rect 17870 25062 17899 25108
rect 17795 25004 17899 25062
rect 17795 24958 17824 25004
rect 17870 24958 17899 25004
rect 17795 24900 17899 24958
rect 17795 24854 17824 24900
rect 17870 24854 17899 24900
rect 17795 24796 17899 24854
rect 17795 24750 17824 24796
rect 17870 24750 17899 24796
rect 17795 24692 17899 24750
rect 17795 24646 17824 24692
rect 17870 24646 17899 24692
rect 17795 24633 17899 24646
rect 18019 26888 18107 26901
rect 18019 26842 18048 26888
rect 18094 26842 18107 26888
rect 18019 26783 18107 26842
rect 18019 26737 18048 26783
rect 18094 26737 18107 26783
rect 18019 26678 18107 26737
rect 18019 26632 18048 26678
rect 18094 26632 18107 26678
rect 18019 26573 18107 26632
rect 18019 26527 18048 26573
rect 18094 26527 18107 26573
rect 18019 26468 18107 26527
rect 18019 26422 18048 26468
rect 18094 26422 18107 26468
rect 18019 26363 18107 26422
rect 18019 26317 18048 26363
rect 18094 26317 18107 26363
rect 18019 26258 18107 26317
rect 18019 26212 18048 26258
rect 18094 26212 18107 26258
rect 18019 26153 18107 26212
rect 18019 26107 18048 26153
rect 18094 26107 18107 26153
rect 18019 26048 18107 26107
rect 18019 26002 18048 26048
rect 18094 26002 18107 26048
rect 18019 25943 18107 26002
rect 18019 25897 18048 25943
rect 18094 25897 18107 25943
rect 18019 25838 18107 25897
rect 18019 25792 18048 25838
rect 18094 25792 18107 25838
rect 18019 25733 18107 25792
rect 18019 25687 18048 25733
rect 18094 25687 18107 25733
rect 18019 25628 18107 25687
rect 18019 25582 18048 25628
rect 18094 25582 18107 25628
rect 18019 25524 18107 25582
rect 18019 25478 18048 25524
rect 18094 25478 18107 25524
rect 18019 25420 18107 25478
rect 18019 25374 18048 25420
rect 18094 25374 18107 25420
rect 18019 25316 18107 25374
rect 18019 25270 18048 25316
rect 18094 25270 18107 25316
rect 18019 25212 18107 25270
rect 18019 25166 18048 25212
rect 18094 25166 18107 25212
rect 18019 25108 18107 25166
rect 18019 25062 18048 25108
rect 18094 25062 18107 25108
rect 18019 25004 18107 25062
rect 18019 24958 18048 25004
rect 18094 24958 18107 25004
rect 18019 24900 18107 24958
rect 18019 24854 18048 24900
rect 18094 24854 18107 24900
rect 18019 24796 18107 24854
rect 18019 24750 18048 24796
rect 18094 24750 18107 24796
rect 18019 24692 18107 24750
rect 18019 24646 18048 24692
rect 18094 24646 18107 24692
rect 18019 24633 18107 24646
rect 18325 26888 18413 26901
rect 18325 26842 18338 26888
rect 18384 26842 18413 26888
rect 18325 26783 18413 26842
rect 18325 26737 18338 26783
rect 18384 26737 18413 26783
rect 18325 26678 18413 26737
rect 18325 26632 18338 26678
rect 18384 26632 18413 26678
rect 18325 26573 18413 26632
rect 18325 26527 18338 26573
rect 18384 26527 18413 26573
rect 18325 26468 18413 26527
rect 18325 26422 18338 26468
rect 18384 26422 18413 26468
rect 18325 26363 18413 26422
rect 18325 26317 18338 26363
rect 18384 26317 18413 26363
rect 18325 26258 18413 26317
rect 18325 26212 18338 26258
rect 18384 26212 18413 26258
rect 18325 26153 18413 26212
rect 18325 26107 18338 26153
rect 18384 26107 18413 26153
rect 18325 26048 18413 26107
rect 18325 26002 18338 26048
rect 18384 26002 18413 26048
rect 18325 25943 18413 26002
rect 18325 25897 18338 25943
rect 18384 25897 18413 25943
rect 18325 25838 18413 25897
rect 18325 25792 18338 25838
rect 18384 25792 18413 25838
rect 18325 25733 18413 25792
rect 18325 25687 18338 25733
rect 18384 25687 18413 25733
rect 18325 25628 18413 25687
rect 18325 25582 18338 25628
rect 18384 25582 18413 25628
rect 18325 25524 18413 25582
rect 18325 25478 18338 25524
rect 18384 25478 18413 25524
rect 18325 25420 18413 25478
rect 18325 25374 18338 25420
rect 18384 25374 18413 25420
rect 18325 25316 18413 25374
rect 18325 25270 18338 25316
rect 18384 25270 18413 25316
rect 18325 25212 18413 25270
rect 18325 25166 18338 25212
rect 18384 25166 18413 25212
rect 18325 25108 18413 25166
rect 18325 25062 18338 25108
rect 18384 25062 18413 25108
rect 18325 25004 18413 25062
rect 18325 24958 18338 25004
rect 18384 24958 18413 25004
rect 18325 24900 18413 24958
rect 18325 24854 18338 24900
rect 18384 24854 18413 24900
rect 18325 24796 18413 24854
rect 18325 24750 18338 24796
rect 18384 24750 18413 24796
rect 18325 24692 18413 24750
rect 18325 24646 18338 24692
rect 18384 24646 18413 24692
rect 18325 24633 18413 24646
rect 18533 26888 18637 26901
rect 18533 26842 18562 26888
rect 18608 26842 18637 26888
rect 18533 26783 18637 26842
rect 18533 26737 18562 26783
rect 18608 26737 18637 26783
rect 18533 26678 18637 26737
rect 18533 26632 18562 26678
rect 18608 26632 18637 26678
rect 18533 26573 18637 26632
rect 18533 26527 18562 26573
rect 18608 26527 18637 26573
rect 18533 26468 18637 26527
rect 18533 26422 18562 26468
rect 18608 26422 18637 26468
rect 18533 26363 18637 26422
rect 18533 26317 18562 26363
rect 18608 26317 18637 26363
rect 18533 26258 18637 26317
rect 18533 26212 18562 26258
rect 18608 26212 18637 26258
rect 18533 26153 18637 26212
rect 18533 26107 18562 26153
rect 18608 26107 18637 26153
rect 18533 26048 18637 26107
rect 18533 26002 18562 26048
rect 18608 26002 18637 26048
rect 18533 25943 18637 26002
rect 18533 25897 18562 25943
rect 18608 25897 18637 25943
rect 18533 25838 18637 25897
rect 18533 25792 18562 25838
rect 18608 25792 18637 25838
rect 18533 25733 18637 25792
rect 18533 25687 18562 25733
rect 18608 25687 18637 25733
rect 18533 25628 18637 25687
rect 18533 25582 18562 25628
rect 18608 25582 18637 25628
rect 18533 25524 18637 25582
rect 18533 25478 18562 25524
rect 18608 25478 18637 25524
rect 18533 25420 18637 25478
rect 18533 25374 18562 25420
rect 18608 25374 18637 25420
rect 18533 25316 18637 25374
rect 18533 25270 18562 25316
rect 18608 25270 18637 25316
rect 18533 25212 18637 25270
rect 18533 25166 18562 25212
rect 18608 25166 18637 25212
rect 18533 25108 18637 25166
rect 18533 25062 18562 25108
rect 18608 25062 18637 25108
rect 18533 25004 18637 25062
rect 18533 24958 18562 25004
rect 18608 24958 18637 25004
rect 18533 24900 18637 24958
rect 18533 24854 18562 24900
rect 18608 24854 18637 24900
rect 18533 24796 18637 24854
rect 18533 24750 18562 24796
rect 18608 24750 18637 24796
rect 18533 24692 18637 24750
rect 18533 24646 18562 24692
rect 18608 24646 18637 24692
rect 18533 24633 18637 24646
rect 18757 26888 18861 26901
rect 18757 26842 18786 26888
rect 18832 26842 18861 26888
rect 18757 26783 18861 26842
rect 18757 26737 18786 26783
rect 18832 26737 18861 26783
rect 18757 26678 18861 26737
rect 18757 26632 18786 26678
rect 18832 26632 18861 26678
rect 18757 26573 18861 26632
rect 18757 26527 18786 26573
rect 18832 26527 18861 26573
rect 18757 26468 18861 26527
rect 18757 26422 18786 26468
rect 18832 26422 18861 26468
rect 18757 26363 18861 26422
rect 18757 26317 18786 26363
rect 18832 26317 18861 26363
rect 18757 26258 18861 26317
rect 18757 26212 18786 26258
rect 18832 26212 18861 26258
rect 18757 26153 18861 26212
rect 18757 26107 18786 26153
rect 18832 26107 18861 26153
rect 18757 26048 18861 26107
rect 18757 26002 18786 26048
rect 18832 26002 18861 26048
rect 18757 25943 18861 26002
rect 18757 25897 18786 25943
rect 18832 25897 18861 25943
rect 18757 25838 18861 25897
rect 18757 25792 18786 25838
rect 18832 25792 18861 25838
rect 18757 25733 18861 25792
rect 18757 25687 18786 25733
rect 18832 25687 18861 25733
rect 18757 25628 18861 25687
rect 18757 25582 18786 25628
rect 18832 25582 18861 25628
rect 18757 25524 18861 25582
rect 18757 25478 18786 25524
rect 18832 25478 18861 25524
rect 18757 25420 18861 25478
rect 18757 25374 18786 25420
rect 18832 25374 18861 25420
rect 18757 25316 18861 25374
rect 18757 25270 18786 25316
rect 18832 25270 18861 25316
rect 18757 25212 18861 25270
rect 18757 25166 18786 25212
rect 18832 25166 18861 25212
rect 18757 25108 18861 25166
rect 18757 25062 18786 25108
rect 18832 25062 18861 25108
rect 18757 25004 18861 25062
rect 18757 24958 18786 25004
rect 18832 24958 18861 25004
rect 18757 24900 18861 24958
rect 18757 24854 18786 24900
rect 18832 24854 18861 24900
rect 18757 24796 18861 24854
rect 18757 24750 18786 24796
rect 18832 24750 18861 24796
rect 18757 24692 18861 24750
rect 18757 24646 18786 24692
rect 18832 24646 18861 24692
rect 18757 24633 18861 24646
rect 18981 26888 19085 26901
rect 18981 26842 19010 26888
rect 19056 26842 19085 26888
rect 18981 26783 19085 26842
rect 18981 26737 19010 26783
rect 19056 26737 19085 26783
rect 18981 26678 19085 26737
rect 18981 26632 19010 26678
rect 19056 26632 19085 26678
rect 18981 26573 19085 26632
rect 18981 26527 19010 26573
rect 19056 26527 19085 26573
rect 18981 26468 19085 26527
rect 18981 26422 19010 26468
rect 19056 26422 19085 26468
rect 18981 26363 19085 26422
rect 18981 26317 19010 26363
rect 19056 26317 19085 26363
rect 18981 26258 19085 26317
rect 18981 26212 19010 26258
rect 19056 26212 19085 26258
rect 18981 26153 19085 26212
rect 18981 26107 19010 26153
rect 19056 26107 19085 26153
rect 18981 26048 19085 26107
rect 18981 26002 19010 26048
rect 19056 26002 19085 26048
rect 18981 25943 19085 26002
rect 18981 25897 19010 25943
rect 19056 25897 19085 25943
rect 18981 25838 19085 25897
rect 18981 25792 19010 25838
rect 19056 25792 19085 25838
rect 18981 25733 19085 25792
rect 18981 25687 19010 25733
rect 19056 25687 19085 25733
rect 18981 25628 19085 25687
rect 18981 25582 19010 25628
rect 19056 25582 19085 25628
rect 18981 25524 19085 25582
rect 18981 25478 19010 25524
rect 19056 25478 19085 25524
rect 18981 25420 19085 25478
rect 18981 25374 19010 25420
rect 19056 25374 19085 25420
rect 18981 25316 19085 25374
rect 18981 25270 19010 25316
rect 19056 25270 19085 25316
rect 18981 25212 19085 25270
rect 18981 25166 19010 25212
rect 19056 25166 19085 25212
rect 18981 25108 19085 25166
rect 18981 25062 19010 25108
rect 19056 25062 19085 25108
rect 18981 25004 19085 25062
rect 18981 24958 19010 25004
rect 19056 24958 19085 25004
rect 18981 24900 19085 24958
rect 18981 24854 19010 24900
rect 19056 24854 19085 24900
rect 18981 24796 19085 24854
rect 18981 24750 19010 24796
rect 19056 24750 19085 24796
rect 18981 24692 19085 24750
rect 18981 24646 19010 24692
rect 19056 24646 19085 24692
rect 18981 24633 19085 24646
rect 19205 26888 19309 26901
rect 19205 26842 19234 26888
rect 19280 26842 19309 26888
rect 19205 26783 19309 26842
rect 19205 26737 19234 26783
rect 19280 26737 19309 26783
rect 19205 26678 19309 26737
rect 19205 26632 19234 26678
rect 19280 26632 19309 26678
rect 19205 26573 19309 26632
rect 19205 26527 19234 26573
rect 19280 26527 19309 26573
rect 19205 26468 19309 26527
rect 19205 26422 19234 26468
rect 19280 26422 19309 26468
rect 19205 26363 19309 26422
rect 19205 26317 19234 26363
rect 19280 26317 19309 26363
rect 19205 26258 19309 26317
rect 19205 26212 19234 26258
rect 19280 26212 19309 26258
rect 19205 26153 19309 26212
rect 19205 26107 19234 26153
rect 19280 26107 19309 26153
rect 19205 26048 19309 26107
rect 19205 26002 19234 26048
rect 19280 26002 19309 26048
rect 19205 25943 19309 26002
rect 19205 25897 19234 25943
rect 19280 25897 19309 25943
rect 19205 25838 19309 25897
rect 19205 25792 19234 25838
rect 19280 25792 19309 25838
rect 19205 25733 19309 25792
rect 19205 25687 19234 25733
rect 19280 25687 19309 25733
rect 19205 25628 19309 25687
rect 19205 25582 19234 25628
rect 19280 25582 19309 25628
rect 19205 25524 19309 25582
rect 19205 25478 19234 25524
rect 19280 25478 19309 25524
rect 19205 25420 19309 25478
rect 19205 25374 19234 25420
rect 19280 25374 19309 25420
rect 19205 25316 19309 25374
rect 19205 25270 19234 25316
rect 19280 25270 19309 25316
rect 19205 25212 19309 25270
rect 19205 25166 19234 25212
rect 19280 25166 19309 25212
rect 19205 25108 19309 25166
rect 19205 25062 19234 25108
rect 19280 25062 19309 25108
rect 19205 25004 19309 25062
rect 19205 24958 19234 25004
rect 19280 24958 19309 25004
rect 19205 24900 19309 24958
rect 19205 24854 19234 24900
rect 19280 24854 19309 24900
rect 19205 24796 19309 24854
rect 19205 24750 19234 24796
rect 19280 24750 19309 24796
rect 19205 24692 19309 24750
rect 19205 24646 19234 24692
rect 19280 24646 19309 24692
rect 19205 24633 19309 24646
rect 19429 26888 19533 26901
rect 19429 26842 19458 26888
rect 19504 26842 19533 26888
rect 19429 26783 19533 26842
rect 19429 26737 19458 26783
rect 19504 26737 19533 26783
rect 19429 26678 19533 26737
rect 19429 26632 19458 26678
rect 19504 26632 19533 26678
rect 19429 26573 19533 26632
rect 19429 26527 19458 26573
rect 19504 26527 19533 26573
rect 19429 26468 19533 26527
rect 19429 26422 19458 26468
rect 19504 26422 19533 26468
rect 19429 26363 19533 26422
rect 19429 26317 19458 26363
rect 19504 26317 19533 26363
rect 19429 26258 19533 26317
rect 19429 26212 19458 26258
rect 19504 26212 19533 26258
rect 19429 26153 19533 26212
rect 19429 26107 19458 26153
rect 19504 26107 19533 26153
rect 19429 26048 19533 26107
rect 19429 26002 19458 26048
rect 19504 26002 19533 26048
rect 19429 25943 19533 26002
rect 19429 25897 19458 25943
rect 19504 25897 19533 25943
rect 19429 25838 19533 25897
rect 19429 25792 19458 25838
rect 19504 25792 19533 25838
rect 19429 25733 19533 25792
rect 19429 25687 19458 25733
rect 19504 25687 19533 25733
rect 19429 25628 19533 25687
rect 19429 25582 19458 25628
rect 19504 25582 19533 25628
rect 19429 25524 19533 25582
rect 19429 25478 19458 25524
rect 19504 25478 19533 25524
rect 19429 25420 19533 25478
rect 19429 25374 19458 25420
rect 19504 25374 19533 25420
rect 19429 25316 19533 25374
rect 19429 25270 19458 25316
rect 19504 25270 19533 25316
rect 19429 25212 19533 25270
rect 19429 25166 19458 25212
rect 19504 25166 19533 25212
rect 19429 25108 19533 25166
rect 19429 25062 19458 25108
rect 19504 25062 19533 25108
rect 19429 25004 19533 25062
rect 19429 24958 19458 25004
rect 19504 24958 19533 25004
rect 19429 24900 19533 24958
rect 19429 24854 19458 24900
rect 19504 24854 19533 24900
rect 19429 24796 19533 24854
rect 19429 24750 19458 24796
rect 19504 24750 19533 24796
rect 19429 24692 19533 24750
rect 19429 24646 19458 24692
rect 19504 24646 19533 24692
rect 19429 24633 19533 24646
rect 19653 26888 19741 26901
rect 19653 26842 19682 26888
rect 19728 26842 19741 26888
rect 19653 26783 19741 26842
rect 19653 26737 19682 26783
rect 19728 26737 19741 26783
rect 19653 26678 19741 26737
rect 19653 26632 19682 26678
rect 19728 26632 19741 26678
rect 19653 26573 19741 26632
rect 19653 26527 19682 26573
rect 19728 26527 19741 26573
rect 19653 26468 19741 26527
rect 19653 26422 19682 26468
rect 19728 26422 19741 26468
rect 19653 26363 19741 26422
rect 19653 26317 19682 26363
rect 19728 26317 19741 26363
rect 19653 26258 19741 26317
rect 19653 26212 19682 26258
rect 19728 26212 19741 26258
rect 19653 26153 19741 26212
rect 19653 26107 19682 26153
rect 19728 26107 19741 26153
rect 19653 26048 19741 26107
rect 19653 26002 19682 26048
rect 19728 26002 19741 26048
rect 19653 25943 19741 26002
rect 19653 25897 19682 25943
rect 19728 25897 19741 25943
rect 19653 25838 19741 25897
rect 19653 25792 19682 25838
rect 19728 25792 19741 25838
rect 19653 25733 19741 25792
rect 19653 25687 19682 25733
rect 19728 25687 19741 25733
rect 19653 25628 19741 25687
rect 19653 25582 19682 25628
rect 19728 25582 19741 25628
rect 19653 25524 19741 25582
rect 19653 25478 19682 25524
rect 19728 25478 19741 25524
rect 19653 25420 19741 25478
rect 19653 25374 19682 25420
rect 19728 25374 19741 25420
rect 19653 25316 19741 25374
rect 19653 25270 19682 25316
rect 19728 25270 19741 25316
rect 19653 25212 19741 25270
rect 19653 25166 19682 25212
rect 19728 25166 19741 25212
rect 19653 25108 19741 25166
rect 19653 25062 19682 25108
rect 19728 25062 19741 25108
rect 19653 25004 19741 25062
rect 19653 24958 19682 25004
rect 19728 24958 19741 25004
rect 19653 24900 19741 24958
rect 19653 24854 19682 24900
rect 19728 24854 19741 24900
rect 19653 24796 19741 24854
rect 19653 24750 19682 24796
rect 19728 24750 19741 24796
rect 19653 24692 19741 24750
rect 19653 24646 19682 24692
rect 19728 24646 19741 24692
rect 19653 24633 19741 24646
rect 19958 26888 20046 26901
rect 19958 26842 19971 26888
rect 20017 26842 20046 26888
rect 19958 26783 20046 26842
rect 19958 26737 19971 26783
rect 20017 26737 20046 26783
rect 19958 26678 20046 26737
rect 19958 26632 19971 26678
rect 20017 26632 20046 26678
rect 19958 26573 20046 26632
rect 19958 26527 19971 26573
rect 20017 26527 20046 26573
rect 19958 26468 20046 26527
rect 19958 26422 19971 26468
rect 20017 26422 20046 26468
rect 19958 26363 20046 26422
rect 19958 26317 19971 26363
rect 20017 26317 20046 26363
rect 19958 26258 20046 26317
rect 19958 26212 19971 26258
rect 20017 26212 20046 26258
rect 19958 26153 20046 26212
rect 19958 26107 19971 26153
rect 20017 26107 20046 26153
rect 19958 26048 20046 26107
rect 19958 26002 19971 26048
rect 20017 26002 20046 26048
rect 19958 25943 20046 26002
rect 19958 25897 19971 25943
rect 20017 25897 20046 25943
rect 19958 25838 20046 25897
rect 19958 25792 19971 25838
rect 20017 25792 20046 25838
rect 19958 25733 20046 25792
rect 19958 25687 19971 25733
rect 20017 25687 20046 25733
rect 19958 25628 20046 25687
rect 19958 25582 19971 25628
rect 20017 25582 20046 25628
rect 19958 25524 20046 25582
rect 19958 25478 19971 25524
rect 20017 25478 20046 25524
rect 19958 25420 20046 25478
rect 19958 25374 19971 25420
rect 20017 25374 20046 25420
rect 19958 25316 20046 25374
rect 19958 25270 19971 25316
rect 20017 25270 20046 25316
rect 19958 25212 20046 25270
rect 19958 25166 19971 25212
rect 20017 25166 20046 25212
rect 19958 25108 20046 25166
rect 19958 25062 19971 25108
rect 20017 25062 20046 25108
rect 19958 25004 20046 25062
rect 19958 24958 19971 25004
rect 20017 24958 20046 25004
rect 19958 24900 20046 24958
rect 19958 24854 19971 24900
rect 20017 24854 20046 24900
rect 19958 24796 20046 24854
rect 19958 24750 19971 24796
rect 20017 24750 20046 24796
rect 19958 24692 20046 24750
rect 19958 24646 19971 24692
rect 20017 24646 20046 24692
rect 19958 24633 20046 24646
rect 20166 26888 20270 26901
rect 20166 26842 20195 26888
rect 20241 26842 20270 26888
rect 20166 26783 20270 26842
rect 20166 26737 20195 26783
rect 20241 26737 20270 26783
rect 20166 26678 20270 26737
rect 20166 26632 20195 26678
rect 20241 26632 20270 26678
rect 20166 26573 20270 26632
rect 20166 26527 20195 26573
rect 20241 26527 20270 26573
rect 20166 26468 20270 26527
rect 20166 26422 20195 26468
rect 20241 26422 20270 26468
rect 20166 26363 20270 26422
rect 20166 26317 20195 26363
rect 20241 26317 20270 26363
rect 20166 26258 20270 26317
rect 20166 26212 20195 26258
rect 20241 26212 20270 26258
rect 20166 26153 20270 26212
rect 20166 26107 20195 26153
rect 20241 26107 20270 26153
rect 20166 26048 20270 26107
rect 20166 26002 20195 26048
rect 20241 26002 20270 26048
rect 20166 25943 20270 26002
rect 20166 25897 20195 25943
rect 20241 25897 20270 25943
rect 20166 25838 20270 25897
rect 20166 25792 20195 25838
rect 20241 25792 20270 25838
rect 20166 25733 20270 25792
rect 20166 25687 20195 25733
rect 20241 25687 20270 25733
rect 20166 25628 20270 25687
rect 20166 25582 20195 25628
rect 20241 25582 20270 25628
rect 20166 25524 20270 25582
rect 20166 25478 20195 25524
rect 20241 25478 20270 25524
rect 20166 25420 20270 25478
rect 20166 25374 20195 25420
rect 20241 25374 20270 25420
rect 20166 25316 20270 25374
rect 20166 25270 20195 25316
rect 20241 25270 20270 25316
rect 20166 25212 20270 25270
rect 20166 25166 20195 25212
rect 20241 25166 20270 25212
rect 20166 25108 20270 25166
rect 20166 25062 20195 25108
rect 20241 25062 20270 25108
rect 20166 25004 20270 25062
rect 20166 24958 20195 25004
rect 20241 24958 20270 25004
rect 20166 24900 20270 24958
rect 20166 24854 20195 24900
rect 20241 24854 20270 24900
rect 20166 24796 20270 24854
rect 20166 24750 20195 24796
rect 20241 24750 20270 24796
rect 20166 24692 20270 24750
rect 20166 24646 20195 24692
rect 20241 24646 20270 24692
rect 20166 24633 20270 24646
rect 20390 26888 20494 26901
rect 20390 26842 20419 26888
rect 20465 26842 20494 26888
rect 20390 26783 20494 26842
rect 20390 26737 20419 26783
rect 20465 26737 20494 26783
rect 20390 26678 20494 26737
rect 20390 26632 20419 26678
rect 20465 26632 20494 26678
rect 20390 26573 20494 26632
rect 20390 26527 20419 26573
rect 20465 26527 20494 26573
rect 20390 26468 20494 26527
rect 20390 26422 20419 26468
rect 20465 26422 20494 26468
rect 20390 26363 20494 26422
rect 20390 26317 20419 26363
rect 20465 26317 20494 26363
rect 20390 26258 20494 26317
rect 20390 26212 20419 26258
rect 20465 26212 20494 26258
rect 20390 26153 20494 26212
rect 20390 26107 20419 26153
rect 20465 26107 20494 26153
rect 20390 26048 20494 26107
rect 20390 26002 20419 26048
rect 20465 26002 20494 26048
rect 20390 25943 20494 26002
rect 20390 25897 20419 25943
rect 20465 25897 20494 25943
rect 20390 25838 20494 25897
rect 20390 25792 20419 25838
rect 20465 25792 20494 25838
rect 20390 25733 20494 25792
rect 20390 25687 20419 25733
rect 20465 25687 20494 25733
rect 20390 25628 20494 25687
rect 20390 25582 20419 25628
rect 20465 25582 20494 25628
rect 20390 25524 20494 25582
rect 20390 25478 20419 25524
rect 20465 25478 20494 25524
rect 20390 25420 20494 25478
rect 20390 25374 20419 25420
rect 20465 25374 20494 25420
rect 20390 25316 20494 25374
rect 20390 25270 20419 25316
rect 20465 25270 20494 25316
rect 20390 25212 20494 25270
rect 20390 25166 20419 25212
rect 20465 25166 20494 25212
rect 20390 25108 20494 25166
rect 20390 25062 20419 25108
rect 20465 25062 20494 25108
rect 20390 25004 20494 25062
rect 20390 24958 20419 25004
rect 20465 24958 20494 25004
rect 20390 24900 20494 24958
rect 20390 24854 20419 24900
rect 20465 24854 20494 24900
rect 20390 24796 20494 24854
rect 20390 24750 20419 24796
rect 20465 24750 20494 24796
rect 20390 24692 20494 24750
rect 20390 24646 20419 24692
rect 20465 24646 20494 24692
rect 20390 24633 20494 24646
rect 20614 26888 20718 26901
rect 20614 26842 20643 26888
rect 20689 26842 20718 26888
rect 20614 26783 20718 26842
rect 20614 26737 20643 26783
rect 20689 26737 20718 26783
rect 20614 26678 20718 26737
rect 20614 26632 20643 26678
rect 20689 26632 20718 26678
rect 20614 26573 20718 26632
rect 20614 26527 20643 26573
rect 20689 26527 20718 26573
rect 20614 26468 20718 26527
rect 20614 26422 20643 26468
rect 20689 26422 20718 26468
rect 20614 26363 20718 26422
rect 20614 26317 20643 26363
rect 20689 26317 20718 26363
rect 20614 26258 20718 26317
rect 20614 26212 20643 26258
rect 20689 26212 20718 26258
rect 20614 26153 20718 26212
rect 20614 26107 20643 26153
rect 20689 26107 20718 26153
rect 20614 26048 20718 26107
rect 20614 26002 20643 26048
rect 20689 26002 20718 26048
rect 20614 25943 20718 26002
rect 20614 25897 20643 25943
rect 20689 25897 20718 25943
rect 20614 25838 20718 25897
rect 20614 25792 20643 25838
rect 20689 25792 20718 25838
rect 20614 25733 20718 25792
rect 20614 25687 20643 25733
rect 20689 25687 20718 25733
rect 20614 25628 20718 25687
rect 20614 25582 20643 25628
rect 20689 25582 20718 25628
rect 20614 25524 20718 25582
rect 20614 25478 20643 25524
rect 20689 25478 20718 25524
rect 20614 25420 20718 25478
rect 20614 25374 20643 25420
rect 20689 25374 20718 25420
rect 20614 25316 20718 25374
rect 20614 25270 20643 25316
rect 20689 25270 20718 25316
rect 20614 25212 20718 25270
rect 20614 25166 20643 25212
rect 20689 25166 20718 25212
rect 20614 25108 20718 25166
rect 20614 25062 20643 25108
rect 20689 25062 20718 25108
rect 20614 25004 20718 25062
rect 20614 24958 20643 25004
rect 20689 24958 20718 25004
rect 20614 24900 20718 24958
rect 20614 24854 20643 24900
rect 20689 24854 20718 24900
rect 20614 24796 20718 24854
rect 20614 24750 20643 24796
rect 20689 24750 20718 24796
rect 20614 24692 20718 24750
rect 20614 24646 20643 24692
rect 20689 24646 20718 24692
rect 20614 24633 20718 24646
rect 20838 26888 20942 26901
rect 20838 26842 20867 26888
rect 20913 26842 20942 26888
rect 20838 26783 20942 26842
rect 20838 26737 20867 26783
rect 20913 26737 20942 26783
rect 20838 26678 20942 26737
rect 20838 26632 20867 26678
rect 20913 26632 20942 26678
rect 20838 26573 20942 26632
rect 20838 26527 20867 26573
rect 20913 26527 20942 26573
rect 20838 26468 20942 26527
rect 20838 26422 20867 26468
rect 20913 26422 20942 26468
rect 20838 26363 20942 26422
rect 20838 26317 20867 26363
rect 20913 26317 20942 26363
rect 20838 26258 20942 26317
rect 20838 26212 20867 26258
rect 20913 26212 20942 26258
rect 20838 26153 20942 26212
rect 20838 26107 20867 26153
rect 20913 26107 20942 26153
rect 20838 26048 20942 26107
rect 20838 26002 20867 26048
rect 20913 26002 20942 26048
rect 20838 25943 20942 26002
rect 20838 25897 20867 25943
rect 20913 25897 20942 25943
rect 20838 25838 20942 25897
rect 20838 25792 20867 25838
rect 20913 25792 20942 25838
rect 20838 25733 20942 25792
rect 20838 25687 20867 25733
rect 20913 25687 20942 25733
rect 20838 25628 20942 25687
rect 20838 25582 20867 25628
rect 20913 25582 20942 25628
rect 20838 25524 20942 25582
rect 20838 25478 20867 25524
rect 20913 25478 20942 25524
rect 20838 25420 20942 25478
rect 20838 25374 20867 25420
rect 20913 25374 20942 25420
rect 20838 25316 20942 25374
rect 20838 25270 20867 25316
rect 20913 25270 20942 25316
rect 20838 25212 20942 25270
rect 20838 25166 20867 25212
rect 20913 25166 20942 25212
rect 20838 25108 20942 25166
rect 20838 25062 20867 25108
rect 20913 25062 20942 25108
rect 20838 25004 20942 25062
rect 20838 24958 20867 25004
rect 20913 24958 20942 25004
rect 20838 24900 20942 24958
rect 20838 24854 20867 24900
rect 20913 24854 20942 24900
rect 20838 24796 20942 24854
rect 20838 24750 20867 24796
rect 20913 24750 20942 24796
rect 20838 24692 20942 24750
rect 20838 24646 20867 24692
rect 20913 24646 20942 24692
rect 20838 24633 20942 24646
rect 21062 26888 21166 26901
rect 21062 26842 21091 26888
rect 21137 26842 21166 26888
rect 21062 26783 21166 26842
rect 21062 26737 21091 26783
rect 21137 26737 21166 26783
rect 21062 26678 21166 26737
rect 21062 26632 21091 26678
rect 21137 26632 21166 26678
rect 21062 26573 21166 26632
rect 21062 26527 21091 26573
rect 21137 26527 21166 26573
rect 21062 26468 21166 26527
rect 21062 26422 21091 26468
rect 21137 26422 21166 26468
rect 21062 26363 21166 26422
rect 21062 26317 21091 26363
rect 21137 26317 21166 26363
rect 21062 26258 21166 26317
rect 21062 26212 21091 26258
rect 21137 26212 21166 26258
rect 21062 26153 21166 26212
rect 21062 26107 21091 26153
rect 21137 26107 21166 26153
rect 21062 26048 21166 26107
rect 21062 26002 21091 26048
rect 21137 26002 21166 26048
rect 21062 25943 21166 26002
rect 21062 25897 21091 25943
rect 21137 25897 21166 25943
rect 21062 25838 21166 25897
rect 21062 25792 21091 25838
rect 21137 25792 21166 25838
rect 21062 25733 21166 25792
rect 21062 25687 21091 25733
rect 21137 25687 21166 25733
rect 21062 25628 21166 25687
rect 21062 25582 21091 25628
rect 21137 25582 21166 25628
rect 21062 25524 21166 25582
rect 21062 25478 21091 25524
rect 21137 25478 21166 25524
rect 21062 25420 21166 25478
rect 21062 25374 21091 25420
rect 21137 25374 21166 25420
rect 21062 25316 21166 25374
rect 21062 25270 21091 25316
rect 21137 25270 21166 25316
rect 21062 25212 21166 25270
rect 21062 25166 21091 25212
rect 21137 25166 21166 25212
rect 21062 25108 21166 25166
rect 21062 25062 21091 25108
rect 21137 25062 21166 25108
rect 21062 25004 21166 25062
rect 21062 24958 21091 25004
rect 21137 24958 21166 25004
rect 21062 24900 21166 24958
rect 21062 24854 21091 24900
rect 21137 24854 21166 24900
rect 21062 24796 21166 24854
rect 21062 24750 21091 24796
rect 21137 24750 21166 24796
rect 21062 24692 21166 24750
rect 21062 24646 21091 24692
rect 21137 24646 21166 24692
rect 21062 24633 21166 24646
rect 21286 26888 21374 26901
rect 21286 26842 21315 26888
rect 21361 26842 21374 26888
rect 21286 26783 21374 26842
rect 21286 26737 21315 26783
rect 21361 26737 21374 26783
rect 21286 26678 21374 26737
rect 21286 26632 21315 26678
rect 21361 26632 21374 26678
rect 21286 26573 21374 26632
rect 21286 26527 21315 26573
rect 21361 26527 21374 26573
rect 21286 26468 21374 26527
rect 21286 26422 21315 26468
rect 21361 26422 21374 26468
rect 21286 26363 21374 26422
rect 21286 26317 21315 26363
rect 21361 26317 21374 26363
rect 21286 26258 21374 26317
rect 21286 26212 21315 26258
rect 21361 26212 21374 26258
rect 21286 26153 21374 26212
rect 21286 26107 21315 26153
rect 21361 26107 21374 26153
rect 21286 26048 21374 26107
rect 21286 26002 21315 26048
rect 21361 26002 21374 26048
rect 21286 25943 21374 26002
rect 21286 25897 21315 25943
rect 21361 25897 21374 25943
rect 21286 25838 21374 25897
rect 21286 25792 21315 25838
rect 21361 25792 21374 25838
rect 21286 25733 21374 25792
rect 21286 25687 21315 25733
rect 21361 25687 21374 25733
rect 21286 25628 21374 25687
rect 21286 25582 21315 25628
rect 21361 25582 21374 25628
rect 21286 25524 21374 25582
rect 21286 25478 21315 25524
rect 21361 25478 21374 25524
rect 21286 25420 21374 25478
rect 21286 25374 21315 25420
rect 21361 25374 21374 25420
rect 21286 25316 21374 25374
rect 21286 25270 21315 25316
rect 21361 25270 21374 25316
rect 21286 25212 21374 25270
rect 21286 25166 21315 25212
rect 21361 25166 21374 25212
rect 21286 25108 21374 25166
rect 21286 25062 21315 25108
rect 21361 25062 21374 25108
rect 21286 25004 21374 25062
rect 21286 24958 21315 25004
rect 21361 24958 21374 25004
rect 21286 24900 21374 24958
rect 21286 24854 21315 24900
rect 21361 24854 21374 24900
rect 21286 24796 21374 24854
rect 21286 24750 21315 24796
rect 21361 24750 21374 24796
rect 21286 24692 21374 24750
rect 21286 24646 21315 24692
rect 21361 24646 21374 24692
rect 21286 24633 21374 24646
rect 21592 26888 21680 26901
rect 21592 26842 21605 26888
rect 21651 26842 21680 26888
rect 21592 26783 21680 26842
rect 21592 26737 21605 26783
rect 21651 26737 21680 26783
rect 21592 26678 21680 26737
rect 21592 26632 21605 26678
rect 21651 26632 21680 26678
rect 21592 26573 21680 26632
rect 21592 26527 21605 26573
rect 21651 26527 21680 26573
rect 21592 26468 21680 26527
rect 21592 26422 21605 26468
rect 21651 26422 21680 26468
rect 21592 26363 21680 26422
rect 21592 26317 21605 26363
rect 21651 26317 21680 26363
rect 21592 26258 21680 26317
rect 21592 26212 21605 26258
rect 21651 26212 21680 26258
rect 21592 26153 21680 26212
rect 21592 26107 21605 26153
rect 21651 26107 21680 26153
rect 21592 26048 21680 26107
rect 21592 26002 21605 26048
rect 21651 26002 21680 26048
rect 21592 25943 21680 26002
rect 21592 25897 21605 25943
rect 21651 25897 21680 25943
rect 21592 25838 21680 25897
rect 21592 25792 21605 25838
rect 21651 25792 21680 25838
rect 21592 25733 21680 25792
rect 21592 25687 21605 25733
rect 21651 25687 21680 25733
rect 21592 25628 21680 25687
rect 21592 25582 21605 25628
rect 21651 25582 21680 25628
rect 21592 25524 21680 25582
rect 21592 25478 21605 25524
rect 21651 25478 21680 25524
rect 21592 25420 21680 25478
rect 21592 25374 21605 25420
rect 21651 25374 21680 25420
rect 21592 25316 21680 25374
rect 21592 25270 21605 25316
rect 21651 25270 21680 25316
rect 21592 25212 21680 25270
rect 21592 25166 21605 25212
rect 21651 25166 21680 25212
rect 21592 25108 21680 25166
rect 21592 25062 21605 25108
rect 21651 25062 21680 25108
rect 21592 25004 21680 25062
rect 21592 24958 21605 25004
rect 21651 24958 21680 25004
rect 21592 24900 21680 24958
rect 21592 24854 21605 24900
rect 21651 24854 21680 24900
rect 21592 24796 21680 24854
rect 21592 24750 21605 24796
rect 21651 24750 21680 24796
rect 21592 24692 21680 24750
rect 21592 24646 21605 24692
rect 21651 24646 21680 24692
rect 21592 24633 21680 24646
rect 21800 26888 21904 26901
rect 21800 26842 21829 26888
rect 21875 26842 21904 26888
rect 21800 26783 21904 26842
rect 21800 26737 21829 26783
rect 21875 26737 21904 26783
rect 21800 26678 21904 26737
rect 21800 26632 21829 26678
rect 21875 26632 21904 26678
rect 21800 26573 21904 26632
rect 21800 26527 21829 26573
rect 21875 26527 21904 26573
rect 21800 26468 21904 26527
rect 21800 26422 21829 26468
rect 21875 26422 21904 26468
rect 21800 26363 21904 26422
rect 21800 26317 21829 26363
rect 21875 26317 21904 26363
rect 21800 26258 21904 26317
rect 21800 26212 21829 26258
rect 21875 26212 21904 26258
rect 21800 26153 21904 26212
rect 21800 26107 21829 26153
rect 21875 26107 21904 26153
rect 21800 26048 21904 26107
rect 21800 26002 21829 26048
rect 21875 26002 21904 26048
rect 21800 25943 21904 26002
rect 21800 25897 21829 25943
rect 21875 25897 21904 25943
rect 21800 25838 21904 25897
rect 21800 25792 21829 25838
rect 21875 25792 21904 25838
rect 21800 25733 21904 25792
rect 21800 25687 21829 25733
rect 21875 25687 21904 25733
rect 21800 25628 21904 25687
rect 21800 25582 21829 25628
rect 21875 25582 21904 25628
rect 21800 25524 21904 25582
rect 21800 25478 21829 25524
rect 21875 25478 21904 25524
rect 21800 25420 21904 25478
rect 21800 25374 21829 25420
rect 21875 25374 21904 25420
rect 21800 25316 21904 25374
rect 21800 25270 21829 25316
rect 21875 25270 21904 25316
rect 21800 25212 21904 25270
rect 21800 25166 21829 25212
rect 21875 25166 21904 25212
rect 21800 25108 21904 25166
rect 21800 25062 21829 25108
rect 21875 25062 21904 25108
rect 21800 25004 21904 25062
rect 21800 24958 21829 25004
rect 21875 24958 21904 25004
rect 21800 24900 21904 24958
rect 21800 24854 21829 24900
rect 21875 24854 21904 24900
rect 21800 24796 21904 24854
rect 21800 24750 21829 24796
rect 21875 24750 21904 24796
rect 21800 24692 21904 24750
rect 21800 24646 21829 24692
rect 21875 24646 21904 24692
rect 21800 24633 21904 24646
rect 22024 26888 22128 26901
rect 22024 26842 22053 26888
rect 22099 26842 22128 26888
rect 22024 26783 22128 26842
rect 22024 26737 22053 26783
rect 22099 26737 22128 26783
rect 22024 26678 22128 26737
rect 22024 26632 22053 26678
rect 22099 26632 22128 26678
rect 22024 26573 22128 26632
rect 22024 26527 22053 26573
rect 22099 26527 22128 26573
rect 22024 26468 22128 26527
rect 22024 26422 22053 26468
rect 22099 26422 22128 26468
rect 22024 26363 22128 26422
rect 22024 26317 22053 26363
rect 22099 26317 22128 26363
rect 22024 26258 22128 26317
rect 22024 26212 22053 26258
rect 22099 26212 22128 26258
rect 22024 26153 22128 26212
rect 22024 26107 22053 26153
rect 22099 26107 22128 26153
rect 22024 26048 22128 26107
rect 22024 26002 22053 26048
rect 22099 26002 22128 26048
rect 22024 25943 22128 26002
rect 22024 25897 22053 25943
rect 22099 25897 22128 25943
rect 22024 25838 22128 25897
rect 22024 25792 22053 25838
rect 22099 25792 22128 25838
rect 22024 25733 22128 25792
rect 22024 25687 22053 25733
rect 22099 25687 22128 25733
rect 22024 25628 22128 25687
rect 22024 25582 22053 25628
rect 22099 25582 22128 25628
rect 22024 25524 22128 25582
rect 22024 25478 22053 25524
rect 22099 25478 22128 25524
rect 22024 25420 22128 25478
rect 22024 25374 22053 25420
rect 22099 25374 22128 25420
rect 22024 25316 22128 25374
rect 22024 25270 22053 25316
rect 22099 25270 22128 25316
rect 22024 25212 22128 25270
rect 22024 25166 22053 25212
rect 22099 25166 22128 25212
rect 22024 25108 22128 25166
rect 22024 25062 22053 25108
rect 22099 25062 22128 25108
rect 22024 25004 22128 25062
rect 22024 24958 22053 25004
rect 22099 24958 22128 25004
rect 22024 24900 22128 24958
rect 22024 24854 22053 24900
rect 22099 24854 22128 24900
rect 22024 24796 22128 24854
rect 22024 24750 22053 24796
rect 22099 24750 22128 24796
rect 22024 24692 22128 24750
rect 22024 24646 22053 24692
rect 22099 24646 22128 24692
rect 22024 24633 22128 24646
rect 22248 26888 22352 26901
rect 22248 26842 22277 26888
rect 22323 26842 22352 26888
rect 22248 26783 22352 26842
rect 22248 26737 22277 26783
rect 22323 26737 22352 26783
rect 22248 26678 22352 26737
rect 22248 26632 22277 26678
rect 22323 26632 22352 26678
rect 22248 26573 22352 26632
rect 22248 26527 22277 26573
rect 22323 26527 22352 26573
rect 22248 26468 22352 26527
rect 22248 26422 22277 26468
rect 22323 26422 22352 26468
rect 22248 26363 22352 26422
rect 22248 26317 22277 26363
rect 22323 26317 22352 26363
rect 22248 26258 22352 26317
rect 22248 26212 22277 26258
rect 22323 26212 22352 26258
rect 22248 26153 22352 26212
rect 22248 26107 22277 26153
rect 22323 26107 22352 26153
rect 22248 26048 22352 26107
rect 22248 26002 22277 26048
rect 22323 26002 22352 26048
rect 22248 25943 22352 26002
rect 22248 25897 22277 25943
rect 22323 25897 22352 25943
rect 22248 25838 22352 25897
rect 22248 25792 22277 25838
rect 22323 25792 22352 25838
rect 22248 25733 22352 25792
rect 22248 25687 22277 25733
rect 22323 25687 22352 25733
rect 22248 25628 22352 25687
rect 22248 25582 22277 25628
rect 22323 25582 22352 25628
rect 22248 25524 22352 25582
rect 22248 25478 22277 25524
rect 22323 25478 22352 25524
rect 22248 25420 22352 25478
rect 22248 25374 22277 25420
rect 22323 25374 22352 25420
rect 22248 25316 22352 25374
rect 22248 25270 22277 25316
rect 22323 25270 22352 25316
rect 22248 25212 22352 25270
rect 22248 25166 22277 25212
rect 22323 25166 22352 25212
rect 22248 25108 22352 25166
rect 22248 25062 22277 25108
rect 22323 25062 22352 25108
rect 22248 25004 22352 25062
rect 22248 24958 22277 25004
rect 22323 24958 22352 25004
rect 22248 24900 22352 24958
rect 22248 24854 22277 24900
rect 22323 24854 22352 24900
rect 22248 24796 22352 24854
rect 22248 24750 22277 24796
rect 22323 24750 22352 24796
rect 22248 24692 22352 24750
rect 22248 24646 22277 24692
rect 22323 24646 22352 24692
rect 22248 24633 22352 24646
rect 22472 26888 22576 26901
rect 22472 26842 22501 26888
rect 22547 26842 22576 26888
rect 22472 26783 22576 26842
rect 22472 26737 22501 26783
rect 22547 26737 22576 26783
rect 22472 26678 22576 26737
rect 22472 26632 22501 26678
rect 22547 26632 22576 26678
rect 22472 26573 22576 26632
rect 22472 26527 22501 26573
rect 22547 26527 22576 26573
rect 22472 26468 22576 26527
rect 22472 26422 22501 26468
rect 22547 26422 22576 26468
rect 22472 26363 22576 26422
rect 22472 26317 22501 26363
rect 22547 26317 22576 26363
rect 22472 26258 22576 26317
rect 22472 26212 22501 26258
rect 22547 26212 22576 26258
rect 22472 26153 22576 26212
rect 22472 26107 22501 26153
rect 22547 26107 22576 26153
rect 22472 26048 22576 26107
rect 22472 26002 22501 26048
rect 22547 26002 22576 26048
rect 22472 25943 22576 26002
rect 22472 25897 22501 25943
rect 22547 25897 22576 25943
rect 22472 25838 22576 25897
rect 22472 25792 22501 25838
rect 22547 25792 22576 25838
rect 22472 25733 22576 25792
rect 22472 25687 22501 25733
rect 22547 25687 22576 25733
rect 22472 25628 22576 25687
rect 22472 25582 22501 25628
rect 22547 25582 22576 25628
rect 22472 25524 22576 25582
rect 22472 25478 22501 25524
rect 22547 25478 22576 25524
rect 22472 25420 22576 25478
rect 22472 25374 22501 25420
rect 22547 25374 22576 25420
rect 22472 25316 22576 25374
rect 22472 25270 22501 25316
rect 22547 25270 22576 25316
rect 22472 25212 22576 25270
rect 22472 25166 22501 25212
rect 22547 25166 22576 25212
rect 22472 25108 22576 25166
rect 22472 25062 22501 25108
rect 22547 25062 22576 25108
rect 22472 25004 22576 25062
rect 22472 24958 22501 25004
rect 22547 24958 22576 25004
rect 22472 24900 22576 24958
rect 22472 24854 22501 24900
rect 22547 24854 22576 24900
rect 22472 24796 22576 24854
rect 22472 24750 22501 24796
rect 22547 24750 22576 24796
rect 22472 24692 22576 24750
rect 22472 24646 22501 24692
rect 22547 24646 22576 24692
rect 22472 24633 22576 24646
rect 22696 26888 22800 26901
rect 22696 26842 22725 26888
rect 22771 26842 22800 26888
rect 22696 26783 22800 26842
rect 22696 26737 22725 26783
rect 22771 26737 22800 26783
rect 22696 26678 22800 26737
rect 22696 26632 22725 26678
rect 22771 26632 22800 26678
rect 22696 26573 22800 26632
rect 22696 26527 22725 26573
rect 22771 26527 22800 26573
rect 22696 26468 22800 26527
rect 22696 26422 22725 26468
rect 22771 26422 22800 26468
rect 22696 26363 22800 26422
rect 22696 26317 22725 26363
rect 22771 26317 22800 26363
rect 22696 26258 22800 26317
rect 22696 26212 22725 26258
rect 22771 26212 22800 26258
rect 22696 26153 22800 26212
rect 22696 26107 22725 26153
rect 22771 26107 22800 26153
rect 22696 26048 22800 26107
rect 22696 26002 22725 26048
rect 22771 26002 22800 26048
rect 22696 25943 22800 26002
rect 22696 25897 22725 25943
rect 22771 25897 22800 25943
rect 22696 25838 22800 25897
rect 22696 25792 22725 25838
rect 22771 25792 22800 25838
rect 22696 25733 22800 25792
rect 22696 25687 22725 25733
rect 22771 25687 22800 25733
rect 22696 25628 22800 25687
rect 22696 25582 22725 25628
rect 22771 25582 22800 25628
rect 22696 25524 22800 25582
rect 22696 25478 22725 25524
rect 22771 25478 22800 25524
rect 22696 25420 22800 25478
rect 22696 25374 22725 25420
rect 22771 25374 22800 25420
rect 22696 25316 22800 25374
rect 22696 25270 22725 25316
rect 22771 25270 22800 25316
rect 22696 25212 22800 25270
rect 22696 25166 22725 25212
rect 22771 25166 22800 25212
rect 22696 25108 22800 25166
rect 22696 25062 22725 25108
rect 22771 25062 22800 25108
rect 22696 25004 22800 25062
rect 22696 24958 22725 25004
rect 22771 24958 22800 25004
rect 22696 24900 22800 24958
rect 22696 24854 22725 24900
rect 22771 24854 22800 24900
rect 22696 24796 22800 24854
rect 22696 24750 22725 24796
rect 22771 24750 22800 24796
rect 22696 24692 22800 24750
rect 22696 24646 22725 24692
rect 22771 24646 22800 24692
rect 22696 24633 22800 24646
rect 22920 26888 23008 26901
rect 22920 26842 22949 26888
rect 22995 26842 23008 26888
rect 22920 26783 23008 26842
rect 22920 26737 22949 26783
rect 22995 26737 23008 26783
rect 22920 26678 23008 26737
rect 22920 26632 22949 26678
rect 22995 26632 23008 26678
rect 22920 26573 23008 26632
rect 22920 26527 22949 26573
rect 22995 26527 23008 26573
rect 22920 26468 23008 26527
rect 22920 26422 22949 26468
rect 22995 26422 23008 26468
rect 22920 26363 23008 26422
rect 22920 26317 22949 26363
rect 22995 26317 23008 26363
rect 22920 26258 23008 26317
rect 22920 26212 22949 26258
rect 22995 26212 23008 26258
rect 22920 26153 23008 26212
rect 22920 26107 22949 26153
rect 22995 26107 23008 26153
rect 22920 26048 23008 26107
rect 22920 26002 22949 26048
rect 22995 26002 23008 26048
rect 22920 25943 23008 26002
rect 22920 25897 22949 25943
rect 22995 25897 23008 25943
rect 22920 25838 23008 25897
rect 22920 25792 22949 25838
rect 22995 25792 23008 25838
rect 22920 25733 23008 25792
rect 22920 25687 22949 25733
rect 22995 25687 23008 25733
rect 22920 25628 23008 25687
rect 22920 25582 22949 25628
rect 22995 25582 23008 25628
rect 22920 25524 23008 25582
rect 22920 25478 22949 25524
rect 22995 25478 23008 25524
rect 22920 25420 23008 25478
rect 22920 25374 22949 25420
rect 22995 25374 23008 25420
rect 22920 25316 23008 25374
rect 22920 25270 22949 25316
rect 22995 25270 23008 25316
rect 22920 25212 23008 25270
rect 22920 25166 22949 25212
rect 22995 25166 23008 25212
rect 22920 25108 23008 25166
rect 22920 25062 22949 25108
rect 22995 25062 23008 25108
rect 22920 25004 23008 25062
rect 22920 24958 22949 25004
rect 22995 24958 23008 25004
rect 22920 24900 23008 24958
rect 22920 24854 22949 24900
rect 22995 24854 23008 24900
rect 22920 24796 23008 24854
rect 23943 25134 24031 25147
rect 23943 25088 23956 25134
rect 24002 25088 24031 25134
rect 23943 25031 24031 25088
rect 23943 24985 23956 25031
rect 24002 24985 24031 25031
rect 23943 24928 24031 24985
rect 23943 24882 23956 24928
rect 24002 24882 24031 24928
rect 23943 24825 24031 24882
rect 22920 24750 22949 24796
rect 22995 24750 23008 24796
rect 22920 24692 23008 24750
rect 22920 24646 22949 24692
rect 22995 24646 23008 24692
rect 22920 24633 23008 24646
rect 15870 23370 15958 23427
rect 15870 23324 15899 23370
rect 15945 23324 15958 23370
rect 15870 23267 15958 23324
rect 15870 23221 15899 23267
rect 15945 23221 15958 23267
rect 15870 23164 15958 23221
rect 15870 23118 15899 23164
rect 15945 23118 15958 23164
rect 15870 23061 15958 23118
rect 15870 23015 15899 23061
rect 15945 23015 15958 23061
rect 15870 22958 15958 23015
rect 15870 22912 15899 22958
rect 15945 22912 15958 22958
rect 15870 22855 15958 22912
rect 15870 22809 15899 22855
rect 15945 22809 15958 22855
rect 15870 22752 15958 22809
rect 15870 22706 15899 22752
rect 15945 22706 15958 22752
rect 15870 22649 15958 22706
rect 15870 22603 15899 22649
rect 15945 22603 15958 22649
rect 15870 22546 15958 22603
rect 15870 22500 15899 22546
rect 15945 22500 15958 22546
rect 15870 22443 15958 22500
rect 15870 22397 15899 22443
rect 15945 22397 15958 22443
rect 15870 22384 15958 22397
rect 16691 23984 16779 23997
rect 16691 21924 16704 23984
rect 16750 21924 16779 23984
rect 16691 21911 16779 21924
rect 16899 23984 17003 23997
rect 16899 21924 16928 23984
rect 16974 21924 17003 23984
rect 16899 21911 17003 21924
rect 17123 23984 17227 23997
rect 17123 21924 17152 23984
rect 17198 21924 17227 23984
rect 17123 21911 17227 21924
rect 17347 23984 17451 23997
rect 17347 21924 17376 23984
rect 17422 21924 17451 23984
rect 17347 21911 17451 21924
rect 17571 23984 17675 23997
rect 17571 21924 17600 23984
rect 17646 21924 17675 23984
rect 17571 21911 17675 21924
rect 17795 23984 17899 23997
rect 17795 21924 17824 23984
rect 17870 21924 17899 23984
rect 17795 21911 17899 21924
rect 18019 23984 18107 23997
rect 18019 21924 18048 23984
rect 18094 21924 18107 23984
rect 18019 21911 18107 21924
rect 18325 23984 18413 23997
rect 18325 21924 18338 23984
rect 18384 21924 18413 23984
rect 18325 21911 18413 21924
rect 18533 23984 18637 23997
rect 18533 21924 18562 23984
rect 18608 21924 18637 23984
rect 18533 21911 18637 21924
rect 18757 23984 18861 23997
rect 18757 21924 18786 23984
rect 18832 21924 18861 23984
rect 18757 21911 18861 21924
rect 18981 23984 19085 23997
rect 18981 21924 19010 23984
rect 19056 21924 19085 23984
rect 18981 21911 19085 21924
rect 19205 23984 19309 23997
rect 19205 21924 19234 23984
rect 19280 21924 19309 23984
rect 19205 21911 19309 21924
rect 19429 23984 19533 23997
rect 19429 21924 19458 23984
rect 19504 21924 19533 23984
rect 19429 21911 19533 21924
rect 19653 23984 19741 23997
rect 19653 21924 19682 23984
rect 19728 21924 19741 23984
rect 19653 21911 19741 21924
rect 19958 23984 20046 23997
rect 19958 21924 19971 23984
rect 20017 21924 20046 23984
rect 19958 21911 20046 21924
rect 20166 23984 20270 23997
rect 20166 21924 20195 23984
rect 20241 21924 20270 23984
rect 20166 21911 20270 21924
rect 20390 23984 20494 23997
rect 20390 21924 20419 23984
rect 20465 21924 20494 23984
rect 20390 21911 20494 21924
rect 20614 23984 20718 23997
rect 20614 21924 20643 23984
rect 20689 21924 20718 23984
rect 20614 21911 20718 21924
rect 20838 23984 20942 23997
rect 20838 21924 20867 23984
rect 20913 21924 20942 23984
rect 20838 21911 20942 21924
rect 21062 23984 21166 23997
rect 21062 21924 21091 23984
rect 21137 21924 21166 23984
rect 21062 21911 21166 21924
rect 21286 23984 21374 23997
rect 21286 21924 21315 23984
rect 21361 21924 21374 23984
rect 21286 21911 21374 21924
rect 21592 23984 21680 23997
rect 21592 21924 21605 23984
rect 21651 21924 21680 23984
rect 21592 21911 21680 21924
rect 21800 23984 21904 23997
rect 21800 21924 21829 23984
rect 21875 21924 21904 23984
rect 21800 21911 21904 21924
rect 22024 23984 22128 23997
rect 22024 21924 22053 23984
rect 22099 21924 22128 23984
rect 22024 21911 22128 21924
rect 22248 23984 22352 23997
rect 22248 21924 22277 23984
rect 22323 21924 22352 23984
rect 22248 21911 22352 21924
rect 22472 23984 22576 23997
rect 22472 21924 22501 23984
rect 22547 21924 22576 23984
rect 22472 21911 22576 21924
rect 22696 23984 22800 23997
rect 22696 21924 22725 23984
rect 22771 21924 22800 23984
rect 22696 21911 22800 21924
rect 22920 23984 23008 23997
rect 22920 21924 22949 23984
rect 22995 21924 23008 23984
rect 22920 21911 23008 21924
rect 15356 21477 15444 21490
rect 23943 24779 23956 24825
rect 24002 24779 24031 24825
rect 23943 24722 24031 24779
rect 23943 24676 23956 24722
rect 24002 24676 24031 24722
rect 23943 24619 24031 24676
rect 23943 24573 23956 24619
rect 24002 24573 24031 24619
rect 23943 24516 24031 24573
rect 23943 24470 23956 24516
rect 24002 24470 24031 24516
rect 23943 24413 24031 24470
rect 23943 24367 23956 24413
rect 24002 24367 24031 24413
rect 23943 24310 24031 24367
rect 23943 24264 23956 24310
rect 24002 24264 24031 24310
rect 23943 24207 24031 24264
rect 23943 24161 23956 24207
rect 24002 24161 24031 24207
rect 23943 24104 24031 24161
rect 23943 24058 23956 24104
rect 24002 24058 24031 24104
rect 23943 24001 24031 24058
rect 23943 23955 23956 24001
rect 24002 23955 24031 24001
rect 23943 23898 24031 23955
rect 23943 23852 23956 23898
rect 24002 23852 24031 23898
rect 23943 23795 24031 23852
rect 23943 23749 23956 23795
rect 24002 23749 24031 23795
rect 23943 23692 24031 23749
rect 23943 23646 23956 23692
rect 24002 23646 24031 23692
rect 23943 23589 24031 23646
rect 23943 23543 23956 23589
rect 24002 23543 24031 23589
rect 23943 23486 24031 23543
rect 23943 23440 23956 23486
rect 24002 23440 24031 23486
rect 23943 23383 24031 23440
rect 23943 23337 23956 23383
rect 24002 23337 24031 23383
rect 23943 23280 24031 23337
rect 23943 23234 23956 23280
rect 24002 23234 24031 23280
rect 23943 23177 24031 23234
rect 23943 23131 23956 23177
rect 24002 23131 24031 23177
rect 23943 23074 24031 23131
rect 23943 23028 23956 23074
rect 24002 23028 24031 23074
rect 23943 22971 24031 23028
rect 23943 22925 23956 22971
rect 24002 22925 24031 22971
rect 23943 22868 24031 22925
rect 23943 22822 23956 22868
rect 24002 22822 24031 22868
rect 23943 22765 24031 22822
rect 23943 22719 23956 22765
rect 24002 22719 24031 22765
rect 23943 22662 24031 22719
rect 23943 22616 23956 22662
rect 24002 22616 24031 22662
rect 23943 22559 24031 22616
rect 23943 22513 23956 22559
rect 24002 22513 24031 22559
rect 23943 22456 24031 22513
rect 23943 22410 23956 22456
rect 24002 22410 24031 22456
rect 23943 22353 24031 22410
rect 23943 22307 23956 22353
rect 24002 22307 24031 22353
rect 23943 22250 24031 22307
rect 23943 22204 23956 22250
rect 24002 22204 24031 22250
rect 23943 22147 24031 22204
rect 23943 22101 23956 22147
rect 24002 22101 24031 22147
rect 23943 22044 24031 22101
rect 23943 21998 23956 22044
rect 24002 21998 24031 22044
rect 23943 21940 24031 21998
rect 23943 21894 23956 21940
rect 24002 21894 24031 21940
rect 23943 21881 24031 21894
rect 24151 25134 24239 25147
rect 24151 25088 24180 25134
rect 24226 25088 24239 25134
rect 24151 25031 24239 25088
rect 24151 24985 24180 25031
rect 24226 24985 24239 25031
rect 24151 24928 24239 24985
rect 24151 24882 24180 24928
rect 24226 24882 24239 24928
rect 24151 24825 24239 24882
rect 24151 24779 24180 24825
rect 24226 24779 24239 24825
rect 24151 24722 24239 24779
rect 24151 24676 24180 24722
rect 24226 24676 24239 24722
rect 24151 24619 24239 24676
rect 24151 24573 24180 24619
rect 24226 24573 24239 24619
rect 24151 24516 24239 24573
rect 24151 24470 24180 24516
rect 24226 24470 24239 24516
rect 24151 24413 24239 24470
rect 24151 24367 24180 24413
rect 24226 24367 24239 24413
rect 24151 24310 24239 24367
rect 24151 24264 24180 24310
rect 24226 24264 24239 24310
rect 24151 24207 24239 24264
rect 24151 24161 24180 24207
rect 24226 24161 24239 24207
rect 24151 24104 24239 24161
rect 24151 24058 24180 24104
rect 24226 24058 24239 24104
rect 24151 24001 24239 24058
rect 24151 23955 24180 24001
rect 24226 23955 24239 24001
rect 24151 23898 24239 23955
rect 24151 23852 24180 23898
rect 24226 23852 24239 23898
rect 24151 23795 24239 23852
rect 24151 23749 24180 23795
rect 24226 23749 24239 23795
rect 24151 23692 24239 23749
rect 24151 23646 24180 23692
rect 24226 23646 24239 23692
rect 24151 23589 24239 23646
rect 24151 23543 24180 23589
rect 24226 23543 24239 23589
rect 24151 23486 24239 23543
rect 24151 23440 24180 23486
rect 24226 23440 24239 23486
rect 24151 23383 24239 23440
rect 24151 23337 24180 23383
rect 24226 23337 24239 23383
rect 24151 23280 24239 23337
rect 24151 23234 24180 23280
rect 24226 23234 24239 23280
rect 24151 23177 24239 23234
rect 24151 23131 24180 23177
rect 24226 23131 24239 23177
rect 24151 23074 24239 23131
rect 24151 23028 24180 23074
rect 24226 23028 24239 23074
rect 24151 22971 24239 23028
rect 24151 22925 24180 22971
rect 24226 22925 24239 22971
rect 24151 22868 24239 22925
rect 24151 22822 24180 22868
rect 24226 22822 24239 22868
rect 24151 22765 24239 22822
rect 24151 22719 24180 22765
rect 24226 22719 24239 22765
rect 24151 22662 24239 22719
rect 24151 22616 24180 22662
rect 24226 22616 24239 22662
rect 24151 22559 24239 22616
rect 24151 22513 24180 22559
rect 24226 22513 24239 22559
rect 24151 22456 24239 22513
rect 24151 22410 24180 22456
rect 24226 22410 24239 22456
rect 24151 22353 24239 22410
rect 24151 22307 24180 22353
rect 24226 22307 24239 22353
rect 24151 22250 24239 22307
rect 24151 22204 24180 22250
rect 24226 22204 24239 22250
rect 24151 22147 24239 22204
rect 24151 22101 24180 22147
rect 24226 22101 24239 22147
rect 24151 22044 24239 22101
rect 24151 21998 24180 22044
rect 24226 21998 24239 22044
rect 24151 21940 24239 21998
rect 24151 21894 24180 21940
rect 24226 21894 24239 21940
rect 24151 21881 24239 21894
rect 24457 25134 24545 25147
rect 24457 25088 24470 25134
rect 24516 25088 24545 25134
rect 24457 25031 24545 25088
rect 24457 24985 24470 25031
rect 24516 24985 24545 25031
rect 24457 24928 24545 24985
rect 24457 24882 24470 24928
rect 24516 24882 24545 24928
rect 24457 24825 24545 24882
rect 24457 24779 24470 24825
rect 24516 24779 24545 24825
rect 24457 24722 24545 24779
rect 24457 24676 24470 24722
rect 24516 24676 24545 24722
rect 24457 24619 24545 24676
rect 24457 24573 24470 24619
rect 24516 24573 24545 24619
rect 24457 24516 24545 24573
rect 24457 24470 24470 24516
rect 24516 24470 24545 24516
rect 24457 24413 24545 24470
rect 24457 24367 24470 24413
rect 24516 24367 24545 24413
rect 24457 24310 24545 24367
rect 24457 24264 24470 24310
rect 24516 24264 24545 24310
rect 24457 24207 24545 24264
rect 24457 24161 24470 24207
rect 24516 24161 24545 24207
rect 24457 24104 24545 24161
rect 24457 24058 24470 24104
rect 24516 24058 24545 24104
rect 24457 24001 24545 24058
rect 24457 23955 24470 24001
rect 24516 23955 24545 24001
rect 24457 23898 24545 23955
rect 24457 23852 24470 23898
rect 24516 23852 24545 23898
rect 24457 23795 24545 23852
rect 24457 23749 24470 23795
rect 24516 23749 24545 23795
rect 24457 23692 24545 23749
rect 24457 23646 24470 23692
rect 24516 23646 24545 23692
rect 24457 23589 24545 23646
rect 24457 23543 24470 23589
rect 24516 23543 24545 23589
rect 24457 23486 24545 23543
rect 24457 23440 24470 23486
rect 24516 23440 24545 23486
rect 24457 23383 24545 23440
rect 24457 23337 24470 23383
rect 24516 23337 24545 23383
rect 24457 23280 24545 23337
rect 24457 23234 24470 23280
rect 24516 23234 24545 23280
rect 24457 23177 24545 23234
rect 24457 23131 24470 23177
rect 24516 23131 24545 23177
rect 24457 23074 24545 23131
rect 24457 23028 24470 23074
rect 24516 23028 24545 23074
rect 24457 22971 24545 23028
rect 24457 22925 24470 22971
rect 24516 22925 24545 22971
rect 24457 22868 24545 22925
rect 24457 22822 24470 22868
rect 24516 22822 24545 22868
rect 24457 22765 24545 22822
rect 24457 22719 24470 22765
rect 24516 22719 24545 22765
rect 24457 22662 24545 22719
rect 24457 22616 24470 22662
rect 24516 22616 24545 22662
rect 24457 22559 24545 22616
rect 24457 22513 24470 22559
rect 24516 22513 24545 22559
rect 24457 22456 24545 22513
rect 24457 22410 24470 22456
rect 24516 22410 24545 22456
rect 24457 22353 24545 22410
rect 24457 22307 24470 22353
rect 24516 22307 24545 22353
rect 24457 22250 24545 22307
rect 24457 22204 24470 22250
rect 24516 22204 24545 22250
rect 24457 22147 24545 22204
rect 24457 22101 24470 22147
rect 24516 22101 24545 22147
rect 24457 22044 24545 22101
rect 24457 21998 24470 22044
rect 24516 21998 24545 22044
rect 24457 21940 24545 21998
rect 24457 21894 24470 21940
rect 24516 21894 24545 21940
rect 24457 21881 24545 21894
rect 24665 25134 24753 25147
rect 24665 25088 24694 25134
rect 24740 25088 24753 25134
rect 24665 25031 24753 25088
rect 24665 24985 24694 25031
rect 24740 24985 24753 25031
rect 24665 24928 24753 24985
rect 24665 24882 24694 24928
rect 24740 24882 24753 24928
rect 24665 24825 24753 24882
rect 24665 24779 24694 24825
rect 24740 24779 24753 24825
rect 25633 25134 25721 25147
rect 25633 25088 25646 25134
rect 25692 25088 25721 25134
rect 25633 25031 25721 25088
rect 25633 24985 25646 25031
rect 25692 24985 25721 25031
rect 25633 24928 25721 24985
rect 25633 24882 25646 24928
rect 25692 24882 25721 24928
rect 25633 24825 25721 24882
rect 24665 24722 24753 24779
rect 24665 24676 24694 24722
rect 24740 24676 24753 24722
rect 24665 24619 24753 24676
rect 24665 24573 24694 24619
rect 24740 24573 24753 24619
rect 24665 24516 24753 24573
rect 24665 24470 24694 24516
rect 24740 24470 24753 24516
rect 24665 24413 24753 24470
rect 24665 24367 24694 24413
rect 24740 24367 24753 24413
rect 24665 24310 24753 24367
rect 24665 24264 24694 24310
rect 24740 24264 24753 24310
rect 24665 24207 24753 24264
rect 24665 24161 24694 24207
rect 24740 24161 24753 24207
rect 24665 24104 24753 24161
rect 24665 24058 24694 24104
rect 24740 24058 24753 24104
rect 24665 24001 24753 24058
rect 24665 23955 24694 24001
rect 24740 23955 24753 24001
rect 24665 23898 24753 23955
rect 24665 23852 24694 23898
rect 24740 23852 24753 23898
rect 24665 23795 24753 23852
rect 24665 23749 24694 23795
rect 24740 23749 24753 23795
rect 24665 23692 24753 23749
rect 24665 23646 24694 23692
rect 24740 23646 24753 23692
rect 24665 23589 24753 23646
rect 24665 23543 24694 23589
rect 24740 23543 24753 23589
rect 24665 23486 24753 23543
rect 24665 23440 24694 23486
rect 24740 23440 24753 23486
rect 24665 23383 24753 23440
rect 24665 23337 24694 23383
rect 24740 23337 24753 23383
rect 24665 23280 24753 23337
rect 24665 23234 24694 23280
rect 24740 23234 24753 23280
rect 24665 23177 24753 23234
rect 24665 23131 24694 23177
rect 24740 23131 24753 23177
rect 24665 23074 24753 23131
rect 24665 23028 24694 23074
rect 24740 23028 24753 23074
rect 24665 22971 24753 23028
rect 24665 22925 24694 22971
rect 24740 22925 24753 22971
rect 24665 22868 24753 22925
rect 24665 22822 24694 22868
rect 24740 22822 24753 22868
rect 24665 22765 24753 22822
rect 24665 22719 24694 22765
rect 24740 22719 24753 22765
rect 24665 22662 24753 22719
rect 24665 22616 24694 22662
rect 24740 22616 24753 22662
rect 24665 22559 24753 22616
rect 24665 22513 24694 22559
rect 24740 22513 24753 22559
rect 24665 22456 24753 22513
rect 24665 22410 24694 22456
rect 24740 22410 24753 22456
rect 24665 22353 24753 22410
rect 24665 22307 24694 22353
rect 24740 22307 24753 22353
rect 24665 22250 24753 22307
rect 24665 22204 24694 22250
rect 24740 22204 24753 22250
rect 24665 22147 24753 22204
rect 24665 22101 24694 22147
rect 24740 22101 24753 22147
rect 24665 22044 24753 22101
rect 24665 21998 24694 22044
rect 24740 21998 24753 22044
rect 24665 21940 24753 21998
rect 24665 21894 24694 21940
rect 24740 21894 24753 21940
rect 24665 21881 24753 21894
rect 25633 24779 25646 24825
rect 25692 24779 25721 24825
rect 25633 24722 25721 24779
rect 25633 24676 25646 24722
rect 25692 24676 25721 24722
rect 25633 24619 25721 24676
rect 25633 24573 25646 24619
rect 25692 24573 25721 24619
rect 25633 24516 25721 24573
rect 25633 24470 25646 24516
rect 25692 24470 25721 24516
rect 25633 24413 25721 24470
rect 25633 24367 25646 24413
rect 25692 24367 25721 24413
rect 25633 24310 25721 24367
rect 25633 24264 25646 24310
rect 25692 24264 25721 24310
rect 25633 24207 25721 24264
rect 25633 24161 25646 24207
rect 25692 24161 25721 24207
rect 25633 24104 25721 24161
rect 25633 24058 25646 24104
rect 25692 24058 25721 24104
rect 25633 24001 25721 24058
rect 25633 23955 25646 24001
rect 25692 23955 25721 24001
rect 25633 23898 25721 23955
rect 25633 23852 25646 23898
rect 25692 23852 25721 23898
rect 25633 23795 25721 23852
rect 25633 23749 25646 23795
rect 25692 23749 25721 23795
rect 25633 23692 25721 23749
rect 25633 23646 25646 23692
rect 25692 23646 25721 23692
rect 25633 23589 25721 23646
rect 25633 23543 25646 23589
rect 25692 23543 25721 23589
rect 25633 23486 25721 23543
rect 25633 23440 25646 23486
rect 25692 23440 25721 23486
rect 25633 23383 25721 23440
rect 25633 23337 25646 23383
rect 25692 23337 25721 23383
rect 25633 23280 25721 23337
rect 25633 23234 25646 23280
rect 25692 23234 25721 23280
rect 25633 23177 25721 23234
rect 25633 23131 25646 23177
rect 25692 23131 25721 23177
rect 25633 23074 25721 23131
rect 25633 23028 25646 23074
rect 25692 23028 25721 23074
rect 25633 22971 25721 23028
rect 25633 22925 25646 22971
rect 25692 22925 25721 22971
rect 25633 22868 25721 22925
rect 25633 22822 25646 22868
rect 25692 22822 25721 22868
rect 25633 22765 25721 22822
rect 25633 22719 25646 22765
rect 25692 22719 25721 22765
rect 25633 22662 25721 22719
rect 25633 22616 25646 22662
rect 25692 22616 25721 22662
rect 25633 22559 25721 22616
rect 25633 22513 25646 22559
rect 25692 22513 25721 22559
rect 25633 22456 25721 22513
rect 25633 22410 25646 22456
rect 25692 22410 25721 22456
rect 25633 22353 25721 22410
rect 25633 22307 25646 22353
rect 25692 22307 25721 22353
rect 25633 22250 25721 22307
rect 25633 22204 25646 22250
rect 25692 22204 25721 22250
rect 25633 22147 25721 22204
rect 25633 22101 25646 22147
rect 25692 22101 25721 22147
rect 25633 22044 25721 22101
rect 25633 21998 25646 22044
rect 25692 21998 25721 22044
rect 25633 21940 25721 21998
rect 25633 21894 25646 21940
rect 25692 21894 25721 21940
rect 25633 21881 25721 21894
rect 25841 25134 25929 25147
rect 25841 25088 25870 25134
rect 25916 25088 25929 25134
rect 25841 25031 25929 25088
rect 25841 24985 25870 25031
rect 25916 24985 25929 25031
rect 25841 24928 25929 24985
rect 25841 24882 25870 24928
rect 25916 24882 25929 24928
rect 25841 24825 25929 24882
rect 25841 24779 25870 24825
rect 25916 24779 25929 24825
rect 25841 24722 25929 24779
rect 25841 24676 25870 24722
rect 25916 24676 25929 24722
rect 25841 24619 25929 24676
rect 25841 24573 25870 24619
rect 25916 24573 25929 24619
rect 25841 24516 25929 24573
rect 25841 24470 25870 24516
rect 25916 24470 25929 24516
rect 25841 24413 25929 24470
rect 25841 24367 25870 24413
rect 25916 24367 25929 24413
rect 25841 24310 25929 24367
rect 25841 24264 25870 24310
rect 25916 24264 25929 24310
rect 25841 24207 25929 24264
rect 25841 24161 25870 24207
rect 25916 24161 25929 24207
rect 25841 24104 25929 24161
rect 25841 24058 25870 24104
rect 25916 24058 25929 24104
rect 25841 24001 25929 24058
rect 25841 23955 25870 24001
rect 25916 23955 25929 24001
rect 25841 23898 25929 23955
rect 25841 23852 25870 23898
rect 25916 23852 25929 23898
rect 25841 23795 25929 23852
rect 25841 23749 25870 23795
rect 25916 23749 25929 23795
rect 25841 23692 25929 23749
rect 25841 23646 25870 23692
rect 25916 23646 25929 23692
rect 25841 23589 25929 23646
rect 25841 23543 25870 23589
rect 25916 23543 25929 23589
rect 25841 23486 25929 23543
rect 25841 23440 25870 23486
rect 25916 23440 25929 23486
rect 25841 23383 25929 23440
rect 25841 23337 25870 23383
rect 25916 23337 25929 23383
rect 25841 23280 25929 23337
rect 25841 23234 25870 23280
rect 25916 23234 25929 23280
rect 25841 23177 25929 23234
rect 25841 23131 25870 23177
rect 25916 23131 25929 23177
rect 25841 23074 25929 23131
rect 25841 23028 25870 23074
rect 25916 23028 25929 23074
rect 25841 22971 25929 23028
rect 25841 22925 25870 22971
rect 25916 22925 25929 22971
rect 25841 22868 25929 22925
rect 25841 22822 25870 22868
rect 25916 22822 25929 22868
rect 25841 22765 25929 22822
rect 25841 22719 25870 22765
rect 25916 22719 25929 22765
rect 25841 22662 25929 22719
rect 25841 22616 25870 22662
rect 25916 22616 25929 22662
rect 25841 22559 25929 22616
rect 25841 22513 25870 22559
rect 25916 22513 25929 22559
rect 25841 22456 25929 22513
rect 25841 22410 25870 22456
rect 25916 22410 25929 22456
rect 25841 22353 25929 22410
rect 25841 22307 25870 22353
rect 25916 22307 25929 22353
rect 25841 22250 25929 22307
rect 25841 22204 25870 22250
rect 25916 22204 25929 22250
rect 25841 22147 25929 22204
rect 25841 22101 25870 22147
rect 25916 22101 25929 22147
rect 25841 22044 25929 22101
rect 25841 21998 25870 22044
rect 25916 21998 25929 22044
rect 25841 21940 25929 21998
rect 25841 21894 25870 21940
rect 25916 21894 25929 21940
rect 25841 21881 25929 21894
rect 26147 25134 26235 25147
rect 26147 25088 26160 25134
rect 26206 25088 26235 25134
rect 26147 25031 26235 25088
rect 26147 24985 26160 25031
rect 26206 24985 26235 25031
rect 26147 24928 26235 24985
rect 26147 24882 26160 24928
rect 26206 24882 26235 24928
rect 26147 24825 26235 24882
rect 26147 24779 26160 24825
rect 26206 24779 26235 24825
rect 26147 24722 26235 24779
rect 26147 24676 26160 24722
rect 26206 24676 26235 24722
rect 26147 24619 26235 24676
rect 26147 24573 26160 24619
rect 26206 24573 26235 24619
rect 26147 24516 26235 24573
rect 26147 24470 26160 24516
rect 26206 24470 26235 24516
rect 26147 24413 26235 24470
rect 26147 24367 26160 24413
rect 26206 24367 26235 24413
rect 26147 24310 26235 24367
rect 26147 24264 26160 24310
rect 26206 24264 26235 24310
rect 26147 24207 26235 24264
rect 26147 24161 26160 24207
rect 26206 24161 26235 24207
rect 26147 24104 26235 24161
rect 26147 24058 26160 24104
rect 26206 24058 26235 24104
rect 26147 24001 26235 24058
rect 26147 23955 26160 24001
rect 26206 23955 26235 24001
rect 26147 23898 26235 23955
rect 26147 23852 26160 23898
rect 26206 23852 26235 23898
rect 26147 23795 26235 23852
rect 26147 23749 26160 23795
rect 26206 23749 26235 23795
rect 26147 23692 26235 23749
rect 26147 23646 26160 23692
rect 26206 23646 26235 23692
rect 26147 23589 26235 23646
rect 26147 23543 26160 23589
rect 26206 23543 26235 23589
rect 26147 23486 26235 23543
rect 26147 23440 26160 23486
rect 26206 23440 26235 23486
rect 26147 23383 26235 23440
rect 26147 23337 26160 23383
rect 26206 23337 26235 23383
rect 26147 23280 26235 23337
rect 26147 23234 26160 23280
rect 26206 23234 26235 23280
rect 26147 23177 26235 23234
rect 26147 23131 26160 23177
rect 26206 23131 26235 23177
rect 26147 23074 26235 23131
rect 26147 23028 26160 23074
rect 26206 23028 26235 23074
rect 26147 22971 26235 23028
rect 26147 22925 26160 22971
rect 26206 22925 26235 22971
rect 26147 22868 26235 22925
rect 26147 22822 26160 22868
rect 26206 22822 26235 22868
rect 26147 22765 26235 22822
rect 26147 22719 26160 22765
rect 26206 22719 26235 22765
rect 26147 22662 26235 22719
rect 26147 22616 26160 22662
rect 26206 22616 26235 22662
rect 26147 22559 26235 22616
rect 26147 22513 26160 22559
rect 26206 22513 26235 22559
rect 26147 22456 26235 22513
rect 26147 22410 26160 22456
rect 26206 22410 26235 22456
rect 26147 22353 26235 22410
rect 26147 22307 26160 22353
rect 26206 22307 26235 22353
rect 26147 22250 26235 22307
rect 26147 22204 26160 22250
rect 26206 22204 26235 22250
rect 26147 22147 26235 22204
rect 26147 22101 26160 22147
rect 26206 22101 26235 22147
rect 26147 22044 26235 22101
rect 26147 21998 26160 22044
rect 26206 21998 26235 22044
rect 26147 21940 26235 21998
rect 26147 21894 26160 21940
rect 26206 21894 26235 21940
rect 26147 21881 26235 21894
rect 26355 25134 26443 25147
rect 26355 25088 26384 25134
rect 26430 25088 26443 25134
rect 26355 25031 26443 25088
rect 26355 24985 26384 25031
rect 26430 24985 26443 25031
rect 26355 24928 26443 24985
rect 26355 24882 26384 24928
rect 26430 24882 26443 24928
rect 26355 24825 26443 24882
rect 26355 24779 26384 24825
rect 26430 24779 26443 24825
rect 27324 25134 27412 25147
rect 27324 25088 27337 25134
rect 27383 25088 27412 25134
rect 27324 25031 27412 25088
rect 27324 24985 27337 25031
rect 27383 24985 27412 25031
rect 27324 24928 27412 24985
rect 27324 24882 27337 24928
rect 27383 24882 27412 24928
rect 27324 24825 27412 24882
rect 26355 24722 26443 24779
rect 26355 24676 26384 24722
rect 26430 24676 26443 24722
rect 26355 24619 26443 24676
rect 26355 24573 26384 24619
rect 26430 24573 26443 24619
rect 26355 24516 26443 24573
rect 26355 24470 26384 24516
rect 26430 24470 26443 24516
rect 26355 24413 26443 24470
rect 26355 24367 26384 24413
rect 26430 24367 26443 24413
rect 26355 24310 26443 24367
rect 26355 24264 26384 24310
rect 26430 24264 26443 24310
rect 26355 24207 26443 24264
rect 26355 24161 26384 24207
rect 26430 24161 26443 24207
rect 26355 24104 26443 24161
rect 26355 24058 26384 24104
rect 26430 24058 26443 24104
rect 26355 24001 26443 24058
rect 26355 23955 26384 24001
rect 26430 23955 26443 24001
rect 26355 23898 26443 23955
rect 26355 23852 26384 23898
rect 26430 23852 26443 23898
rect 26355 23795 26443 23852
rect 26355 23749 26384 23795
rect 26430 23749 26443 23795
rect 26355 23692 26443 23749
rect 26355 23646 26384 23692
rect 26430 23646 26443 23692
rect 26355 23589 26443 23646
rect 26355 23543 26384 23589
rect 26430 23543 26443 23589
rect 26355 23486 26443 23543
rect 26355 23440 26384 23486
rect 26430 23440 26443 23486
rect 26355 23383 26443 23440
rect 26355 23337 26384 23383
rect 26430 23337 26443 23383
rect 26355 23280 26443 23337
rect 26355 23234 26384 23280
rect 26430 23234 26443 23280
rect 26355 23177 26443 23234
rect 26355 23131 26384 23177
rect 26430 23131 26443 23177
rect 26355 23074 26443 23131
rect 26355 23028 26384 23074
rect 26430 23028 26443 23074
rect 26355 22971 26443 23028
rect 26355 22925 26384 22971
rect 26430 22925 26443 22971
rect 26355 22868 26443 22925
rect 26355 22822 26384 22868
rect 26430 22822 26443 22868
rect 26355 22765 26443 22822
rect 26355 22719 26384 22765
rect 26430 22719 26443 22765
rect 26355 22662 26443 22719
rect 26355 22616 26384 22662
rect 26430 22616 26443 22662
rect 26355 22559 26443 22616
rect 26355 22513 26384 22559
rect 26430 22513 26443 22559
rect 26355 22456 26443 22513
rect 26355 22410 26384 22456
rect 26430 22410 26443 22456
rect 26355 22353 26443 22410
rect 26355 22307 26384 22353
rect 26430 22307 26443 22353
rect 26355 22250 26443 22307
rect 26355 22204 26384 22250
rect 26430 22204 26443 22250
rect 26355 22147 26443 22204
rect 26355 22101 26384 22147
rect 26430 22101 26443 22147
rect 26355 22044 26443 22101
rect 26355 21998 26384 22044
rect 26430 21998 26443 22044
rect 26355 21940 26443 21998
rect 26355 21894 26384 21940
rect 26430 21894 26443 21940
rect 26355 21881 26443 21894
rect 27324 24779 27337 24825
rect 27383 24779 27412 24825
rect 27324 24722 27412 24779
rect 27324 24676 27337 24722
rect 27383 24676 27412 24722
rect 27324 24619 27412 24676
rect 27324 24573 27337 24619
rect 27383 24573 27412 24619
rect 27324 24516 27412 24573
rect 27324 24470 27337 24516
rect 27383 24470 27412 24516
rect 27324 24413 27412 24470
rect 27324 24367 27337 24413
rect 27383 24367 27412 24413
rect 27324 24310 27412 24367
rect 27324 24264 27337 24310
rect 27383 24264 27412 24310
rect 27324 24207 27412 24264
rect 27324 24161 27337 24207
rect 27383 24161 27412 24207
rect 27324 24104 27412 24161
rect 27324 24058 27337 24104
rect 27383 24058 27412 24104
rect 27324 24001 27412 24058
rect 27324 23955 27337 24001
rect 27383 23955 27412 24001
rect 27324 23898 27412 23955
rect 27324 23852 27337 23898
rect 27383 23852 27412 23898
rect 27324 23795 27412 23852
rect 27324 23749 27337 23795
rect 27383 23749 27412 23795
rect 27324 23692 27412 23749
rect 27324 23646 27337 23692
rect 27383 23646 27412 23692
rect 27324 23589 27412 23646
rect 27324 23543 27337 23589
rect 27383 23543 27412 23589
rect 27324 23486 27412 23543
rect 27324 23440 27337 23486
rect 27383 23440 27412 23486
rect 27324 23383 27412 23440
rect 27324 23337 27337 23383
rect 27383 23337 27412 23383
rect 27324 23280 27412 23337
rect 27324 23234 27337 23280
rect 27383 23234 27412 23280
rect 27324 23177 27412 23234
rect 27324 23131 27337 23177
rect 27383 23131 27412 23177
rect 27324 23074 27412 23131
rect 27324 23028 27337 23074
rect 27383 23028 27412 23074
rect 27324 22971 27412 23028
rect 27324 22925 27337 22971
rect 27383 22925 27412 22971
rect 27324 22868 27412 22925
rect 27324 22822 27337 22868
rect 27383 22822 27412 22868
rect 27324 22765 27412 22822
rect 27324 22719 27337 22765
rect 27383 22719 27412 22765
rect 27324 22662 27412 22719
rect 27324 22616 27337 22662
rect 27383 22616 27412 22662
rect 27324 22559 27412 22616
rect 27324 22513 27337 22559
rect 27383 22513 27412 22559
rect 27324 22456 27412 22513
rect 27324 22410 27337 22456
rect 27383 22410 27412 22456
rect 27324 22353 27412 22410
rect 27324 22307 27337 22353
rect 27383 22307 27412 22353
rect 27324 22250 27412 22307
rect 27324 22204 27337 22250
rect 27383 22204 27412 22250
rect 27324 22147 27412 22204
rect 27324 22101 27337 22147
rect 27383 22101 27412 22147
rect 27324 22044 27412 22101
rect 27324 21998 27337 22044
rect 27383 21998 27412 22044
rect 27324 21940 27412 21998
rect 27324 21894 27337 21940
rect 27383 21894 27412 21940
rect 27324 21881 27412 21894
rect 27532 25134 27620 25147
rect 27532 25088 27561 25134
rect 27607 25088 27620 25134
rect 27532 25031 27620 25088
rect 27532 24985 27561 25031
rect 27607 24985 27620 25031
rect 27532 24928 27620 24985
rect 27532 24882 27561 24928
rect 27607 24882 27620 24928
rect 27532 24825 27620 24882
rect 27532 24779 27561 24825
rect 27607 24779 27620 24825
rect 27532 24722 27620 24779
rect 27532 24676 27561 24722
rect 27607 24676 27620 24722
rect 27532 24619 27620 24676
rect 27532 24573 27561 24619
rect 27607 24573 27620 24619
rect 27532 24516 27620 24573
rect 27532 24470 27561 24516
rect 27607 24470 27620 24516
rect 27532 24413 27620 24470
rect 27532 24367 27561 24413
rect 27607 24367 27620 24413
rect 27532 24310 27620 24367
rect 27532 24264 27561 24310
rect 27607 24264 27620 24310
rect 27532 24207 27620 24264
rect 27532 24161 27561 24207
rect 27607 24161 27620 24207
rect 27532 24104 27620 24161
rect 27532 24058 27561 24104
rect 27607 24058 27620 24104
rect 27532 24001 27620 24058
rect 27532 23955 27561 24001
rect 27607 23955 27620 24001
rect 27532 23898 27620 23955
rect 27532 23852 27561 23898
rect 27607 23852 27620 23898
rect 27532 23795 27620 23852
rect 27532 23749 27561 23795
rect 27607 23749 27620 23795
rect 27532 23692 27620 23749
rect 27532 23646 27561 23692
rect 27607 23646 27620 23692
rect 27532 23589 27620 23646
rect 27532 23543 27561 23589
rect 27607 23543 27620 23589
rect 27532 23486 27620 23543
rect 27532 23440 27561 23486
rect 27607 23440 27620 23486
rect 27532 23383 27620 23440
rect 27532 23337 27561 23383
rect 27607 23337 27620 23383
rect 27532 23280 27620 23337
rect 27532 23234 27561 23280
rect 27607 23234 27620 23280
rect 27532 23177 27620 23234
rect 27532 23131 27561 23177
rect 27607 23131 27620 23177
rect 27532 23074 27620 23131
rect 27532 23028 27561 23074
rect 27607 23028 27620 23074
rect 27532 22971 27620 23028
rect 27532 22925 27561 22971
rect 27607 22925 27620 22971
rect 27532 22868 27620 22925
rect 27532 22822 27561 22868
rect 27607 22822 27620 22868
rect 27532 22765 27620 22822
rect 27532 22719 27561 22765
rect 27607 22719 27620 22765
rect 27532 22662 27620 22719
rect 27532 22616 27561 22662
rect 27607 22616 27620 22662
rect 27532 22559 27620 22616
rect 27532 22513 27561 22559
rect 27607 22513 27620 22559
rect 27532 22456 27620 22513
rect 27532 22410 27561 22456
rect 27607 22410 27620 22456
rect 27532 22353 27620 22410
rect 27532 22307 27561 22353
rect 27607 22307 27620 22353
rect 27532 22250 27620 22307
rect 27532 22204 27561 22250
rect 27607 22204 27620 22250
rect 27532 22147 27620 22204
rect 27532 22101 27561 22147
rect 27607 22101 27620 22147
rect 27532 22044 27620 22101
rect 27532 21998 27561 22044
rect 27607 21998 27620 22044
rect 27532 21940 27620 21998
rect 27532 21894 27561 21940
rect 27607 21894 27620 21940
rect 27532 21881 27620 21894
rect 27838 25134 27926 25147
rect 27838 25088 27851 25134
rect 27897 25088 27926 25134
rect 27838 25031 27926 25088
rect 27838 24985 27851 25031
rect 27897 24985 27926 25031
rect 27838 24928 27926 24985
rect 27838 24882 27851 24928
rect 27897 24882 27926 24928
rect 27838 24825 27926 24882
rect 27838 24779 27851 24825
rect 27897 24779 27926 24825
rect 27838 24722 27926 24779
rect 27838 24676 27851 24722
rect 27897 24676 27926 24722
rect 27838 24619 27926 24676
rect 27838 24573 27851 24619
rect 27897 24573 27926 24619
rect 27838 24516 27926 24573
rect 27838 24470 27851 24516
rect 27897 24470 27926 24516
rect 27838 24413 27926 24470
rect 27838 24367 27851 24413
rect 27897 24367 27926 24413
rect 27838 24310 27926 24367
rect 27838 24264 27851 24310
rect 27897 24264 27926 24310
rect 27838 24207 27926 24264
rect 27838 24161 27851 24207
rect 27897 24161 27926 24207
rect 27838 24104 27926 24161
rect 27838 24058 27851 24104
rect 27897 24058 27926 24104
rect 27838 24001 27926 24058
rect 27838 23955 27851 24001
rect 27897 23955 27926 24001
rect 27838 23898 27926 23955
rect 27838 23852 27851 23898
rect 27897 23852 27926 23898
rect 27838 23795 27926 23852
rect 27838 23749 27851 23795
rect 27897 23749 27926 23795
rect 27838 23692 27926 23749
rect 27838 23646 27851 23692
rect 27897 23646 27926 23692
rect 27838 23589 27926 23646
rect 27838 23543 27851 23589
rect 27897 23543 27926 23589
rect 27838 23486 27926 23543
rect 27838 23440 27851 23486
rect 27897 23440 27926 23486
rect 27838 23383 27926 23440
rect 27838 23337 27851 23383
rect 27897 23337 27926 23383
rect 27838 23280 27926 23337
rect 27838 23234 27851 23280
rect 27897 23234 27926 23280
rect 27838 23177 27926 23234
rect 27838 23131 27851 23177
rect 27897 23131 27926 23177
rect 27838 23074 27926 23131
rect 27838 23028 27851 23074
rect 27897 23028 27926 23074
rect 27838 22971 27926 23028
rect 27838 22925 27851 22971
rect 27897 22925 27926 22971
rect 27838 22868 27926 22925
rect 27838 22822 27851 22868
rect 27897 22822 27926 22868
rect 27838 22765 27926 22822
rect 27838 22719 27851 22765
rect 27897 22719 27926 22765
rect 27838 22662 27926 22719
rect 27838 22616 27851 22662
rect 27897 22616 27926 22662
rect 27838 22559 27926 22616
rect 27838 22513 27851 22559
rect 27897 22513 27926 22559
rect 27838 22456 27926 22513
rect 27838 22410 27851 22456
rect 27897 22410 27926 22456
rect 27838 22353 27926 22410
rect 27838 22307 27851 22353
rect 27897 22307 27926 22353
rect 27838 22250 27926 22307
rect 27838 22204 27851 22250
rect 27897 22204 27926 22250
rect 27838 22147 27926 22204
rect 27838 22101 27851 22147
rect 27897 22101 27926 22147
rect 27838 22044 27926 22101
rect 27838 21998 27851 22044
rect 27897 21998 27926 22044
rect 27838 21940 27926 21998
rect 27838 21894 27851 21940
rect 27897 21894 27926 21940
rect 27838 21881 27926 21894
rect 28046 25134 28134 25147
rect 28046 25088 28075 25134
rect 28121 25088 28134 25134
rect 28046 25031 28134 25088
rect 28046 24985 28075 25031
rect 28121 24985 28134 25031
rect 28046 24928 28134 24985
rect 28046 24882 28075 24928
rect 28121 24882 28134 24928
rect 28046 24825 28134 24882
rect 28046 24779 28075 24825
rect 28121 24779 28134 24825
rect 28046 24722 28134 24779
rect 28046 24676 28075 24722
rect 28121 24676 28134 24722
rect 28046 24619 28134 24676
rect 28046 24573 28075 24619
rect 28121 24573 28134 24619
rect 28046 24516 28134 24573
rect 28046 24470 28075 24516
rect 28121 24470 28134 24516
rect 28046 24413 28134 24470
rect 28046 24367 28075 24413
rect 28121 24367 28134 24413
rect 28046 24310 28134 24367
rect 28046 24264 28075 24310
rect 28121 24264 28134 24310
rect 28046 24207 28134 24264
rect 28046 24161 28075 24207
rect 28121 24161 28134 24207
rect 28046 24104 28134 24161
rect 28046 24058 28075 24104
rect 28121 24058 28134 24104
rect 28046 24001 28134 24058
rect 28046 23955 28075 24001
rect 28121 23955 28134 24001
rect 28046 23898 28134 23955
rect 28046 23852 28075 23898
rect 28121 23852 28134 23898
rect 28046 23795 28134 23852
rect 28046 23749 28075 23795
rect 28121 23749 28134 23795
rect 28046 23692 28134 23749
rect 28046 23646 28075 23692
rect 28121 23646 28134 23692
rect 28046 23589 28134 23646
rect 28046 23543 28075 23589
rect 28121 23543 28134 23589
rect 28046 23486 28134 23543
rect 28046 23440 28075 23486
rect 28121 23440 28134 23486
rect 28046 23383 28134 23440
rect 28046 23337 28075 23383
rect 28121 23337 28134 23383
rect 28046 23280 28134 23337
rect 28046 23234 28075 23280
rect 28121 23234 28134 23280
rect 28046 23177 28134 23234
rect 28046 23131 28075 23177
rect 28121 23131 28134 23177
rect 28046 23074 28134 23131
rect 28046 23028 28075 23074
rect 28121 23028 28134 23074
rect 28046 22971 28134 23028
rect 28046 22925 28075 22971
rect 28121 22925 28134 22971
rect 28046 22868 28134 22925
rect 28046 22822 28075 22868
rect 28121 22822 28134 22868
rect 28046 22765 28134 22822
rect 28046 22719 28075 22765
rect 28121 22719 28134 22765
rect 28046 22662 28134 22719
rect 28046 22616 28075 22662
rect 28121 22616 28134 22662
rect 28046 22559 28134 22616
rect 28046 22513 28075 22559
rect 28121 22513 28134 22559
rect 28046 22456 28134 22513
rect 28046 22410 28075 22456
rect 28121 22410 28134 22456
rect 28046 22353 28134 22410
rect 28046 22307 28075 22353
rect 28121 22307 28134 22353
rect 28046 22250 28134 22307
rect 28046 22204 28075 22250
rect 28121 22204 28134 22250
rect 28046 22147 28134 22204
rect 28046 22101 28075 22147
rect 28121 22101 28134 22147
rect 28046 22044 28134 22101
rect 28046 21998 28075 22044
rect 28121 21998 28134 22044
rect 28046 21940 28134 21998
rect 28046 21894 28075 21940
rect 28121 21894 28134 21940
rect 28046 21881 28134 21894
rect 1982 16572 2070 16585
rect 1982 12598 1995 16572
rect 2041 12598 2070 16572
rect 1982 12585 2070 12598
rect 2190 16572 2278 16585
rect 2190 12598 2219 16572
rect 2265 12598 2278 16572
rect 2190 12585 2278 12598
rect 2430 16572 2518 16585
rect 2430 12598 2443 16572
rect 2489 12598 2518 16572
rect 2430 12585 2518 12598
rect 2638 16572 2742 16585
rect 2638 12598 2667 16572
rect 2713 12598 2742 16572
rect 2638 12585 2742 12598
rect 2862 16572 2966 16585
rect 2862 12598 2891 16572
rect 2937 12598 2966 16572
rect 2862 12585 2966 12598
rect 3086 16572 3190 16585
rect 3086 12598 3115 16572
rect 3161 12598 3190 16572
rect 3086 12585 3190 12598
rect 3310 16572 3398 16585
rect 3310 12598 3339 16572
rect 3385 12598 3398 16572
rect 3310 12585 3398 12598
rect 3550 16572 3638 16585
rect 3550 12598 3563 16572
rect 3609 12598 3638 16572
rect 3550 12585 3638 12598
rect 3758 16572 3862 16585
rect 3758 12598 3787 16572
rect 3833 12598 3862 16572
rect 3758 12585 3862 12598
rect 3982 16572 4086 16585
rect 3982 12598 4011 16572
rect 4057 12598 4086 16572
rect 3982 12585 4086 12598
rect 4206 16572 4310 16585
rect 4206 12598 4235 16572
rect 4281 12598 4310 16572
rect 4206 12585 4310 12598
rect 4430 16572 4518 16585
rect 4430 12598 4459 16572
rect 4505 12598 4518 16572
rect 4430 12585 4518 12598
rect 4670 16572 4758 16585
rect 4670 12598 4683 16572
rect 4729 12598 4758 16572
rect 4670 12585 4758 12598
rect 4878 16572 4982 16585
rect 4878 12598 4907 16572
rect 4953 12598 4982 16572
rect 4878 12585 4982 12598
rect 5102 16572 5206 16585
rect 5102 12598 5131 16572
rect 5177 12598 5206 16572
rect 5102 12585 5206 12598
rect 5326 16572 5430 16585
rect 5326 12598 5355 16572
rect 5401 12598 5430 16572
rect 5326 12585 5430 12598
rect 5550 16572 5638 16585
rect 5550 12598 5579 16572
rect 5625 12598 5638 16572
rect 5550 12585 5638 12598
rect 5790 16572 5878 16585
rect 5790 12598 5803 16572
rect 5849 12598 5878 16572
rect 5790 12585 5878 12598
rect 5998 16572 6102 16585
rect 5998 12598 6027 16572
rect 6073 12598 6102 16572
rect 5998 12585 6102 12598
rect 6222 16572 6326 16585
rect 6222 12598 6251 16572
rect 6297 12598 6326 16572
rect 6222 12585 6326 12598
rect 6446 16572 6550 16585
rect 6446 12598 6475 16572
rect 6521 12598 6550 16572
rect 6446 12585 6550 12598
rect 6670 16572 6758 16585
rect 6670 12598 6699 16572
rect 6745 12598 6758 16572
rect 6670 12585 6758 12598
rect 6910 16572 6998 16585
rect 6910 12598 6923 16572
rect 6969 12598 6998 16572
rect 6910 12585 6998 12598
rect 7118 16572 7222 16585
rect 7118 12598 7147 16572
rect 7193 12598 7222 16572
rect 7118 12585 7222 12598
rect 7342 16572 7446 16585
rect 7342 12598 7371 16572
rect 7417 12598 7446 16572
rect 7342 12585 7446 12598
rect 7566 16572 7670 16585
rect 7566 12598 7595 16572
rect 7641 12598 7670 16572
rect 7566 12585 7670 12598
rect 7790 16572 7878 16585
rect 7790 12598 7819 16572
rect 7865 12598 7878 16572
rect 7790 12585 7878 12598
rect 8030 16572 8118 16585
rect 8030 12598 8043 16572
rect 8089 12598 8118 16572
rect 8030 12585 8118 12598
rect 8238 16572 8342 16585
rect 8238 12598 8267 16572
rect 8313 12598 8342 16572
rect 8238 12585 8342 12598
rect 8462 16572 8566 16585
rect 8462 12598 8491 16572
rect 8537 12598 8566 16572
rect 8462 12585 8566 12598
rect 8686 16572 8790 16585
rect 8686 12598 8715 16572
rect 8761 12598 8790 16572
rect 8686 12585 8790 12598
rect 8910 16572 8998 16585
rect 8910 12598 8939 16572
rect 8985 12598 8998 16572
rect 8910 12585 8998 12598
rect 9150 16572 9238 16585
rect 9150 12598 9163 16572
rect 9209 12598 9238 16572
rect 9150 12585 9238 12598
rect 9358 16572 9462 16585
rect 9358 12598 9387 16572
rect 9433 12598 9462 16572
rect 9358 12585 9462 12598
rect 9582 16572 9686 16585
rect 9582 12598 9611 16572
rect 9657 12598 9686 16572
rect 9582 12585 9686 12598
rect 9806 16572 9910 16585
rect 9806 12598 9835 16572
rect 9881 12598 9910 16572
rect 9806 12585 9910 12598
rect 10030 16572 10118 16585
rect 10030 12598 10059 16572
rect 10105 12598 10118 16572
rect 10030 12585 10118 12598
rect 10270 16572 10358 16585
rect 10270 12598 10283 16572
rect 10329 12598 10358 16572
rect 10270 12585 10358 12598
rect 10478 16572 10582 16585
rect 10478 12598 10507 16572
rect 10553 12598 10582 16572
rect 10478 12585 10582 12598
rect 10702 16572 10806 16585
rect 10702 12598 10731 16572
rect 10777 12598 10806 16572
rect 10702 12585 10806 12598
rect 10926 16572 11030 16585
rect 10926 12598 10955 16572
rect 11001 12598 11030 16572
rect 10926 12585 11030 12598
rect 11150 16572 11238 16585
rect 11150 12598 11179 16572
rect 11225 12598 11238 16572
rect 11150 12585 11238 12598
rect 11390 16572 11478 16585
rect 11390 12598 11403 16572
rect 11449 12598 11478 16572
rect 11390 12585 11478 12598
rect 11598 16572 11702 16585
rect 11598 12598 11627 16572
rect 11673 12598 11702 16572
rect 11598 12585 11702 12598
rect 11822 16572 11926 16585
rect 11822 12598 11851 16572
rect 11897 12598 11926 16572
rect 11822 12585 11926 12598
rect 12046 16572 12150 16585
rect 12046 12598 12075 16572
rect 12121 12598 12150 16572
rect 12046 12585 12150 12598
rect 12270 16572 12358 16585
rect 12270 12598 12299 16572
rect 12345 12598 12358 16572
rect 12270 12585 12358 12598
rect 12510 16572 12598 16585
rect 12510 12598 12523 16572
rect 12569 12598 12598 16572
rect 12510 12585 12598 12598
rect 12718 16572 12822 16585
rect 12718 12598 12747 16572
rect 12793 12598 12822 16572
rect 12718 12585 12822 12598
rect 12942 16572 13046 16585
rect 12942 12598 12971 16572
rect 13017 12598 13046 16572
rect 12942 12585 13046 12598
rect 13166 16572 13270 16585
rect 13166 12598 13195 16572
rect 13241 12598 13270 16572
rect 13166 12585 13270 12598
rect 13390 16572 13478 16585
rect 13390 12598 13419 16572
rect 13465 12598 13478 16572
rect 13390 12585 13478 12598
rect 13630 16572 13718 16585
rect 13630 12598 13643 16572
rect 13689 12598 13718 16572
rect 13630 12585 13718 12598
rect 13838 16572 13942 16585
rect 13838 12598 13867 16572
rect 13913 12598 13942 16572
rect 13838 12585 13942 12598
rect 14062 16572 14166 16585
rect 14062 12598 14091 16572
rect 14137 12598 14166 16572
rect 14062 12585 14166 12598
rect 14286 16572 14390 16585
rect 14286 12598 14315 16572
rect 14361 12598 14390 16572
rect 14286 12585 14390 12598
rect 14510 16572 14598 16585
rect 14510 12598 14539 16572
rect 14585 12598 14598 16572
rect 14510 12585 14598 12598
rect 14750 16572 14838 16585
rect 14750 12598 14763 16572
rect 14809 12598 14838 16572
rect 14750 12585 14838 12598
rect 14958 16572 15062 16585
rect 14958 12598 14987 16572
rect 15033 12598 15062 16572
rect 14958 12585 15062 12598
rect 15182 16572 15286 16585
rect 15182 12598 15211 16572
rect 15257 12598 15286 16572
rect 15182 12585 15286 12598
rect 15406 16572 15510 16585
rect 15406 12598 15435 16572
rect 15481 12598 15510 16572
rect 15406 12585 15510 12598
rect 15630 16572 15718 16585
rect 15630 12598 15659 16572
rect 15705 12598 15718 16572
rect 15630 12585 15718 12598
rect 15870 16572 15958 16585
rect 15870 12598 15883 16572
rect 15929 12598 15958 16572
rect 15870 12585 15958 12598
rect 16078 16572 16182 16585
rect 16078 12598 16107 16572
rect 16153 12598 16182 16572
rect 16078 12585 16182 12598
rect 16302 16572 16406 16585
rect 16302 12598 16331 16572
rect 16377 12598 16406 16572
rect 16302 12585 16406 12598
rect 16526 16572 16630 16585
rect 16526 12598 16555 16572
rect 16601 12598 16630 16572
rect 16526 12585 16630 12598
rect 16750 16572 16838 16585
rect 16750 12598 16779 16572
rect 16825 12598 16838 16572
rect 16750 12585 16838 12598
rect 16990 16572 17078 16585
rect 16990 12598 17003 16572
rect 17049 12598 17078 16572
rect 16990 12585 17078 12598
rect 17198 16572 17302 16585
rect 17198 12598 17227 16572
rect 17273 12598 17302 16572
rect 17198 12585 17302 12598
rect 17422 16572 17526 16585
rect 17422 12598 17451 16572
rect 17497 12598 17526 16572
rect 17422 12585 17526 12598
rect 17646 16572 17750 16585
rect 17646 12598 17675 16572
rect 17721 12598 17750 16572
rect 17646 12585 17750 12598
rect 17870 16572 17958 16585
rect 17870 12598 17899 16572
rect 17945 12598 17958 16572
rect 17870 12585 17958 12598
rect 18110 16572 18198 16585
rect 18110 12598 18123 16572
rect 18169 12598 18198 16572
rect 18110 12585 18198 12598
rect 18318 16572 18422 16585
rect 18318 12598 18347 16572
rect 18393 12598 18422 16572
rect 18318 12585 18422 12598
rect 18542 16572 18646 16585
rect 18542 12598 18571 16572
rect 18617 12598 18646 16572
rect 18542 12585 18646 12598
rect 18766 16572 18870 16585
rect 18766 12598 18795 16572
rect 18841 12598 18870 16572
rect 18766 12585 18870 12598
rect 18990 16572 19078 16585
rect 18990 12598 19019 16572
rect 19065 12598 19078 16572
rect 18990 12585 19078 12598
rect 19230 16572 19318 16585
rect 19230 12598 19243 16572
rect 19289 12598 19318 16572
rect 19230 12585 19318 12598
rect 19438 16572 19542 16585
rect 19438 12598 19467 16572
rect 19513 12598 19542 16572
rect 19438 12585 19542 12598
rect 19662 16572 19766 16585
rect 19662 12598 19691 16572
rect 19737 12598 19766 16572
rect 19662 12585 19766 12598
rect 19886 16572 19974 16585
rect 19886 12598 19915 16572
rect 19961 12598 19974 16572
rect 19886 12585 19974 12598
rect 7437 8273 7525 8286
rect 7437 8227 7450 8273
rect 7496 8227 7525 8273
rect 7437 8164 7525 8227
rect 7437 8118 7450 8164
rect 7496 8118 7525 8164
rect 7437 8055 7525 8118
rect 7437 8009 7450 8055
rect 7496 8009 7525 8055
rect 2608 7964 2696 7977
rect 2608 5268 2621 7964
rect 2667 5268 2696 7964
rect 2608 5255 2696 5268
rect 2816 7964 2904 7977
rect 2816 5268 2845 7964
rect 2891 5268 2904 7964
rect 2816 5255 2904 5268
rect 3122 7964 3210 7977
rect 3122 5268 3135 7964
rect 3181 5268 3210 7964
rect 3122 5255 3210 5268
rect 3330 7964 3418 7977
rect 3330 5268 3359 7964
rect 3405 5268 3418 7964
rect 4299 7964 4387 7977
rect 3330 5255 3418 5268
rect 4299 5268 4312 7964
rect 4358 5268 4387 7964
rect 4299 5255 4387 5268
rect 4507 7964 4595 7977
rect 4507 5268 4536 7964
rect 4582 5268 4595 7964
rect 4507 5255 4595 5268
rect 4813 7964 4901 7977
rect 4813 5268 4826 7964
rect 4872 5268 4901 7964
rect 4813 5255 4901 5268
rect 5021 7964 5109 7977
rect 5021 5268 5050 7964
rect 5096 5268 5109 7964
rect 5990 7964 6078 7977
rect 5021 5255 5109 5268
rect 5990 5268 6003 7964
rect 6049 5268 6078 7964
rect 5990 5255 6078 5268
rect 6198 7964 6286 7977
rect 6198 5268 6227 7964
rect 6273 5268 6286 7964
rect 6198 5255 6286 5268
rect 6504 7964 6592 7977
rect 6504 5268 6517 7964
rect 6563 5268 6592 7964
rect 6504 5255 6592 5268
rect 6712 7964 6800 7977
rect 6712 5268 6741 7964
rect 6787 5268 6800 7964
rect 7437 7947 7525 8009
rect 7437 7901 7450 7947
rect 7496 7901 7525 7947
rect 7437 7839 7525 7901
rect 7437 7793 7450 7839
rect 7496 7793 7525 7839
rect 7437 7731 7525 7793
rect 7437 7685 7450 7731
rect 7496 7685 7525 7731
rect 7437 7623 7525 7685
rect 7437 7577 7450 7623
rect 7496 7577 7525 7623
rect 7437 7515 7525 7577
rect 7437 7469 7450 7515
rect 7496 7469 7525 7515
rect 7437 7407 7525 7469
rect 7437 7361 7450 7407
rect 7496 7361 7525 7407
rect 7437 7299 7525 7361
rect 7437 7253 7450 7299
rect 7496 7253 7525 7299
rect 7437 7191 7525 7253
rect 7437 7145 7450 7191
rect 7496 7145 7525 7191
rect 7437 7132 7525 7145
rect 7645 8273 7749 8286
rect 7645 8227 7674 8273
rect 7720 8227 7749 8273
rect 7645 8164 7749 8227
rect 7645 8118 7674 8164
rect 7720 8118 7749 8164
rect 7645 8055 7749 8118
rect 7645 8009 7674 8055
rect 7720 8009 7749 8055
rect 7645 7947 7749 8009
rect 7645 7901 7674 7947
rect 7720 7901 7749 7947
rect 7645 7839 7749 7901
rect 7645 7793 7674 7839
rect 7720 7793 7749 7839
rect 7645 7731 7749 7793
rect 7645 7685 7674 7731
rect 7720 7685 7749 7731
rect 7645 7623 7749 7685
rect 7645 7577 7674 7623
rect 7720 7577 7749 7623
rect 7645 7515 7749 7577
rect 7645 7469 7674 7515
rect 7720 7469 7749 7515
rect 7645 7407 7749 7469
rect 7645 7361 7674 7407
rect 7720 7361 7749 7407
rect 7645 7299 7749 7361
rect 7645 7253 7674 7299
rect 7720 7253 7749 7299
rect 7645 7191 7749 7253
rect 7645 7145 7674 7191
rect 7720 7145 7749 7191
rect 7645 7132 7749 7145
rect 7869 8273 7973 8286
rect 7869 8227 7898 8273
rect 7944 8227 7973 8273
rect 7869 8164 7973 8227
rect 7869 8118 7898 8164
rect 7944 8118 7973 8164
rect 7869 8055 7973 8118
rect 7869 8009 7898 8055
rect 7944 8009 7973 8055
rect 7869 7947 7973 8009
rect 7869 7901 7898 7947
rect 7944 7901 7973 7947
rect 7869 7839 7973 7901
rect 7869 7793 7898 7839
rect 7944 7793 7973 7839
rect 7869 7731 7973 7793
rect 7869 7685 7898 7731
rect 7944 7685 7973 7731
rect 7869 7623 7973 7685
rect 7869 7577 7898 7623
rect 7944 7577 7973 7623
rect 7869 7515 7973 7577
rect 7869 7469 7898 7515
rect 7944 7469 7973 7515
rect 7869 7407 7973 7469
rect 7869 7361 7898 7407
rect 7944 7361 7973 7407
rect 7869 7299 7973 7361
rect 7869 7253 7898 7299
rect 7944 7253 7973 7299
rect 7869 7191 7973 7253
rect 7869 7145 7898 7191
rect 7944 7145 7973 7191
rect 7869 7132 7973 7145
rect 8093 8273 8197 8286
rect 8093 8227 8122 8273
rect 8168 8227 8197 8273
rect 8093 8164 8197 8227
rect 8093 8118 8122 8164
rect 8168 8118 8197 8164
rect 8093 8055 8197 8118
rect 8093 8009 8122 8055
rect 8168 8009 8197 8055
rect 8093 7947 8197 8009
rect 8093 7901 8122 7947
rect 8168 7901 8197 7947
rect 8093 7839 8197 7901
rect 8093 7793 8122 7839
rect 8168 7793 8197 7839
rect 8093 7731 8197 7793
rect 8093 7685 8122 7731
rect 8168 7685 8197 7731
rect 8093 7623 8197 7685
rect 8093 7577 8122 7623
rect 8168 7577 8197 7623
rect 8093 7515 8197 7577
rect 8093 7469 8122 7515
rect 8168 7469 8197 7515
rect 8093 7407 8197 7469
rect 8093 7361 8122 7407
rect 8168 7361 8197 7407
rect 8093 7299 8197 7361
rect 8093 7253 8122 7299
rect 8168 7253 8197 7299
rect 8093 7191 8197 7253
rect 8093 7145 8122 7191
rect 8168 7145 8197 7191
rect 8093 7132 8197 7145
rect 8317 8273 8421 8286
rect 8317 8227 8346 8273
rect 8392 8227 8421 8273
rect 8317 8164 8421 8227
rect 8317 8118 8346 8164
rect 8392 8118 8421 8164
rect 8317 8055 8421 8118
rect 8317 8009 8346 8055
rect 8392 8009 8421 8055
rect 8317 7947 8421 8009
rect 8317 7901 8346 7947
rect 8392 7901 8421 7947
rect 8317 7839 8421 7901
rect 8317 7793 8346 7839
rect 8392 7793 8421 7839
rect 8317 7731 8421 7793
rect 8317 7685 8346 7731
rect 8392 7685 8421 7731
rect 8317 7623 8421 7685
rect 8317 7577 8346 7623
rect 8392 7577 8421 7623
rect 8317 7515 8421 7577
rect 8317 7469 8346 7515
rect 8392 7469 8421 7515
rect 8317 7407 8421 7469
rect 8317 7361 8346 7407
rect 8392 7361 8421 7407
rect 8317 7299 8421 7361
rect 8317 7253 8346 7299
rect 8392 7253 8421 7299
rect 8317 7191 8421 7253
rect 8317 7145 8346 7191
rect 8392 7145 8421 7191
rect 8317 7132 8421 7145
rect 8541 8273 8645 8286
rect 8541 8227 8570 8273
rect 8616 8227 8645 8273
rect 8541 8164 8645 8227
rect 8541 8118 8570 8164
rect 8616 8118 8645 8164
rect 8541 8055 8645 8118
rect 8541 8009 8570 8055
rect 8616 8009 8645 8055
rect 8541 7947 8645 8009
rect 8541 7901 8570 7947
rect 8616 7901 8645 7947
rect 8541 7839 8645 7901
rect 8541 7793 8570 7839
rect 8616 7793 8645 7839
rect 8541 7731 8645 7793
rect 8541 7685 8570 7731
rect 8616 7685 8645 7731
rect 8541 7623 8645 7685
rect 8541 7577 8570 7623
rect 8616 7577 8645 7623
rect 8541 7515 8645 7577
rect 8541 7469 8570 7515
rect 8616 7469 8645 7515
rect 8541 7407 8645 7469
rect 8541 7361 8570 7407
rect 8616 7361 8645 7407
rect 8541 7299 8645 7361
rect 8541 7253 8570 7299
rect 8616 7253 8645 7299
rect 8541 7191 8645 7253
rect 8541 7145 8570 7191
rect 8616 7145 8645 7191
rect 8541 7132 8645 7145
rect 8765 8273 8853 8286
rect 8765 8227 8794 8273
rect 8840 8227 8853 8273
rect 8765 8164 8853 8227
rect 8765 8118 8794 8164
rect 8840 8118 8853 8164
rect 8765 8055 8853 8118
rect 8765 8009 8794 8055
rect 8840 8009 8853 8055
rect 8765 7947 8853 8009
rect 8765 7901 8794 7947
rect 8840 7901 8853 7947
rect 8765 7839 8853 7901
rect 8765 7793 8794 7839
rect 8840 7793 8853 7839
rect 8765 7731 8853 7793
rect 8765 7685 8794 7731
rect 8840 7685 8853 7731
rect 8765 7623 8853 7685
rect 8765 7577 8794 7623
rect 8840 7577 8853 7623
rect 8765 7515 8853 7577
rect 8765 7469 8794 7515
rect 8840 7469 8853 7515
rect 8765 7407 8853 7469
rect 8765 7361 8794 7407
rect 8840 7361 8853 7407
rect 8765 7299 8853 7361
rect 8765 7253 8794 7299
rect 8840 7253 8853 7299
rect 8765 7191 8853 7253
rect 8765 7145 8794 7191
rect 8840 7145 8853 7191
rect 8765 7132 8853 7145
rect 9070 8273 9158 8286
rect 9070 8227 9083 8273
rect 9129 8227 9158 8273
rect 9070 8164 9158 8227
rect 9070 8118 9083 8164
rect 9129 8118 9158 8164
rect 9070 8055 9158 8118
rect 9070 8009 9083 8055
rect 9129 8009 9158 8055
rect 9070 7947 9158 8009
rect 9070 7901 9083 7947
rect 9129 7901 9158 7947
rect 9070 7839 9158 7901
rect 9070 7793 9083 7839
rect 9129 7793 9158 7839
rect 9070 7731 9158 7793
rect 9070 7685 9083 7731
rect 9129 7685 9158 7731
rect 9070 7623 9158 7685
rect 9070 7577 9083 7623
rect 9129 7577 9158 7623
rect 9070 7515 9158 7577
rect 9070 7469 9083 7515
rect 9129 7469 9158 7515
rect 9070 7407 9158 7469
rect 9070 7361 9083 7407
rect 9129 7361 9158 7407
rect 9070 7299 9158 7361
rect 9070 7253 9083 7299
rect 9129 7253 9158 7299
rect 9070 7191 9158 7253
rect 9070 7145 9083 7191
rect 9129 7145 9158 7191
rect 9070 7132 9158 7145
rect 9278 8273 9382 8286
rect 9278 8227 9307 8273
rect 9353 8227 9382 8273
rect 9278 8164 9382 8227
rect 9278 8118 9307 8164
rect 9353 8118 9382 8164
rect 9278 8055 9382 8118
rect 9278 8009 9307 8055
rect 9353 8009 9382 8055
rect 9278 7947 9382 8009
rect 9278 7901 9307 7947
rect 9353 7901 9382 7947
rect 9278 7839 9382 7901
rect 9278 7793 9307 7839
rect 9353 7793 9382 7839
rect 9278 7731 9382 7793
rect 9278 7685 9307 7731
rect 9353 7685 9382 7731
rect 9278 7623 9382 7685
rect 9278 7577 9307 7623
rect 9353 7577 9382 7623
rect 9278 7515 9382 7577
rect 9278 7469 9307 7515
rect 9353 7469 9382 7515
rect 9278 7407 9382 7469
rect 9278 7361 9307 7407
rect 9353 7361 9382 7407
rect 9278 7299 9382 7361
rect 9278 7253 9307 7299
rect 9353 7253 9382 7299
rect 9278 7191 9382 7253
rect 9278 7145 9307 7191
rect 9353 7145 9382 7191
rect 9278 7132 9382 7145
rect 9502 8273 9606 8286
rect 9502 8227 9531 8273
rect 9577 8227 9606 8273
rect 9502 8164 9606 8227
rect 9502 8118 9531 8164
rect 9577 8118 9606 8164
rect 9502 8055 9606 8118
rect 9502 8009 9531 8055
rect 9577 8009 9606 8055
rect 9502 7947 9606 8009
rect 9502 7901 9531 7947
rect 9577 7901 9606 7947
rect 9502 7839 9606 7901
rect 9502 7793 9531 7839
rect 9577 7793 9606 7839
rect 9502 7731 9606 7793
rect 9502 7685 9531 7731
rect 9577 7685 9606 7731
rect 9502 7623 9606 7685
rect 9502 7577 9531 7623
rect 9577 7577 9606 7623
rect 9502 7515 9606 7577
rect 9502 7469 9531 7515
rect 9577 7469 9606 7515
rect 9502 7407 9606 7469
rect 9502 7361 9531 7407
rect 9577 7361 9606 7407
rect 9502 7299 9606 7361
rect 9502 7253 9531 7299
rect 9577 7253 9606 7299
rect 9502 7191 9606 7253
rect 9502 7145 9531 7191
rect 9577 7145 9606 7191
rect 9502 7132 9606 7145
rect 9726 8273 9830 8286
rect 9726 8227 9755 8273
rect 9801 8227 9830 8273
rect 9726 8164 9830 8227
rect 9726 8118 9755 8164
rect 9801 8118 9830 8164
rect 9726 8055 9830 8118
rect 9726 8009 9755 8055
rect 9801 8009 9830 8055
rect 9726 7947 9830 8009
rect 9726 7901 9755 7947
rect 9801 7901 9830 7947
rect 9726 7839 9830 7901
rect 9726 7793 9755 7839
rect 9801 7793 9830 7839
rect 9726 7731 9830 7793
rect 9726 7685 9755 7731
rect 9801 7685 9830 7731
rect 9726 7623 9830 7685
rect 9726 7577 9755 7623
rect 9801 7577 9830 7623
rect 9726 7515 9830 7577
rect 9726 7469 9755 7515
rect 9801 7469 9830 7515
rect 9726 7407 9830 7469
rect 9726 7361 9755 7407
rect 9801 7361 9830 7407
rect 9726 7299 9830 7361
rect 9726 7253 9755 7299
rect 9801 7253 9830 7299
rect 9726 7191 9830 7253
rect 9726 7145 9755 7191
rect 9801 7145 9830 7191
rect 9726 7132 9830 7145
rect 9950 8273 10054 8286
rect 9950 8227 9979 8273
rect 10025 8227 10054 8273
rect 9950 8164 10054 8227
rect 9950 8118 9979 8164
rect 10025 8118 10054 8164
rect 9950 8055 10054 8118
rect 9950 8009 9979 8055
rect 10025 8009 10054 8055
rect 9950 7947 10054 8009
rect 9950 7901 9979 7947
rect 10025 7901 10054 7947
rect 9950 7839 10054 7901
rect 9950 7793 9979 7839
rect 10025 7793 10054 7839
rect 9950 7731 10054 7793
rect 9950 7685 9979 7731
rect 10025 7685 10054 7731
rect 9950 7623 10054 7685
rect 9950 7577 9979 7623
rect 10025 7577 10054 7623
rect 9950 7515 10054 7577
rect 9950 7469 9979 7515
rect 10025 7469 10054 7515
rect 9950 7407 10054 7469
rect 9950 7361 9979 7407
rect 10025 7361 10054 7407
rect 9950 7299 10054 7361
rect 9950 7253 9979 7299
rect 10025 7253 10054 7299
rect 9950 7191 10054 7253
rect 9950 7145 9979 7191
rect 10025 7145 10054 7191
rect 9950 7132 10054 7145
rect 10174 8273 10278 8286
rect 10174 8227 10203 8273
rect 10249 8227 10278 8273
rect 10174 8164 10278 8227
rect 10174 8118 10203 8164
rect 10249 8118 10278 8164
rect 10174 8055 10278 8118
rect 10174 8009 10203 8055
rect 10249 8009 10278 8055
rect 10174 7947 10278 8009
rect 10174 7901 10203 7947
rect 10249 7901 10278 7947
rect 10174 7839 10278 7901
rect 10174 7793 10203 7839
rect 10249 7793 10278 7839
rect 10174 7731 10278 7793
rect 10174 7685 10203 7731
rect 10249 7685 10278 7731
rect 10174 7623 10278 7685
rect 10174 7577 10203 7623
rect 10249 7577 10278 7623
rect 10174 7515 10278 7577
rect 10174 7469 10203 7515
rect 10249 7469 10278 7515
rect 10174 7407 10278 7469
rect 10174 7361 10203 7407
rect 10249 7361 10278 7407
rect 10174 7299 10278 7361
rect 10174 7253 10203 7299
rect 10249 7253 10278 7299
rect 10174 7191 10278 7253
rect 10174 7145 10203 7191
rect 10249 7145 10278 7191
rect 10174 7132 10278 7145
rect 10398 8273 10486 8286
rect 10398 8227 10427 8273
rect 10473 8227 10486 8273
rect 10398 8164 10486 8227
rect 10398 8118 10427 8164
rect 10473 8118 10486 8164
rect 10398 8055 10486 8118
rect 10398 8009 10427 8055
rect 10473 8009 10486 8055
rect 10398 7947 10486 8009
rect 10398 7901 10427 7947
rect 10473 7901 10486 7947
rect 10398 7839 10486 7901
rect 10398 7793 10427 7839
rect 10473 7793 10486 7839
rect 10398 7731 10486 7793
rect 10398 7685 10427 7731
rect 10473 7685 10486 7731
rect 10398 7623 10486 7685
rect 10398 7577 10427 7623
rect 10473 7577 10486 7623
rect 10398 7515 10486 7577
rect 10398 7469 10427 7515
rect 10473 7469 10486 7515
rect 10398 7407 10486 7469
rect 10398 7361 10427 7407
rect 10473 7361 10486 7407
rect 10398 7299 10486 7361
rect 10398 7253 10427 7299
rect 10473 7253 10486 7299
rect 10398 7191 10486 7253
rect 10398 7145 10427 7191
rect 10473 7145 10486 7191
rect 10398 7132 10486 7145
rect 10704 8273 10792 8286
rect 10704 8227 10717 8273
rect 10763 8227 10792 8273
rect 10704 8164 10792 8227
rect 10704 8118 10717 8164
rect 10763 8118 10792 8164
rect 10704 8055 10792 8118
rect 10704 8009 10717 8055
rect 10763 8009 10792 8055
rect 10704 7947 10792 8009
rect 10704 7901 10717 7947
rect 10763 7901 10792 7947
rect 10704 7839 10792 7901
rect 10704 7793 10717 7839
rect 10763 7793 10792 7839
rect 10704 7731 10792 7793
rect 10704 7685 10717 7731
rect 10763 7685 10792 7731
rect 10704 7623 10792 7685
rect 10704 7577 10717 7623
rect 10763 7577 10792 7623
rect 10704 7515 10792 7577
rect 10704 7469 10717 7515
rect 10763 7469 10792 7515
rect 10704 7407 10792 7469
rect 10704 7361 10717 7407
rect 10763 7361 10792 7407
rect 10704 7299 10792 7361
rect 10704 7253 10717 7299
rect 10763 7253 10792 7299
rect 10704 7191 10792 7253
rect 10704 7145 10717 7191
rect 10763 7145 10792 7191
rect 10704 7132 10792 7145
rect 10912 8273 11016 8286
rect 10912 8227 10941 8273
rect 10987 8227 11016 8273
rect 10912 8164 11016 8227
rect 10912 8118 10941 8164
rect 10987 8118 11016 8164
rect 10912 8055 11016 8118
rect 10912 8009 10941 8055
rect 10987 8009 11016 8055
rect 10912 7947 11016 8009
rect 10912 7901 10941 7947
rect 10987 7901 11016 7947
rect 10912 7839 11016 7901
rect 10912 7793 10941 7839
rect 10987 7793 11016 7839
rect 10912 7731 11016 7793
rect 10912 7685 10941 7731
rect 10987 7685 11016 7731
rect 10912 7623 11016 7685
rect 10912 7577 10941 7623
rect 10987 7577 11016 7623
rect 10912 7515 11016 7577
rect 10912 7469 10941 7515
rect 10987 7469 11016 7515
rect 10912 7407 11016 7469
rect 10912 7361 10941 7407
rect 10987 7361 11016 7407
rect 10912 7299 11016 7361
rect 10912 7253 10941 7299
rect 10987 7253 11016 7299
rect 10912 7191 11016 7253
rect 10912 7145 10941 7191
rect 10987 7145 11016 7191
rect 10912 7132 11016 7145
rect 11136 8273 11240 8286
rect 11136 8227 11165 8273
rect 11211 8227 11240 8273
rect 11136 8164 11240 8227
rect 11136 8118 11165 8164
rect 11211 8118 11240 8164
rect 11136 8055 11240 8118
rect 11136 8009 11165 8055
rect 11211 8009 11240 8055
rect 11136 7947 11240 8009
rect 11136 7901 11165 7947
rect 11211 7901 11240 7947
rect 11136 7839 11240 7901
rect 11136 7793 11165 7839
rect 11211 7793 11240 7839
rect 11136 7731 11240 7793
rect 11136 7685 11165 7731
rect 11211 7685 11240 7731
rect 11136 7623 11240 7685
rect 11136 7577 11165 7623
rect 11211 7577 11240 7623
rect 11136 7515 11240 7577
rect 11136 7469 11165 7515
rect 11211 7469 11240 7515
rect 11136 7407 11240 7469
rect 11136 7361 11165 7407
rect 11211 7361 11240 7407
rect 11136 7299 11240 7361
rect 11136 7253 11165 7299
rect 11211 7253 11240 7299
rect 11136 7191 11240 7253
rect 11136 7145 11165 7191
rect 11211 7145 11240 7191
rect 11136 7132 11240 7145
rect 11360 8273 11464 8286
rect 11360 8227 11389 8273
rect 11435 8227 11464 8273
rect 11360 8164 11464 8227
rect 11360 8118 11389 8164
rect 11435 8118 11464 8164
rect 11360 8055 11464 8118
rect 11360 8009 11389 8055
rect 11435 8009 11464 8055
rect 11360 7947 11464 8009
rect 11360 7901 11389 7947
rect 11435 7901 11464 7947
rect 11360 7839 11464 7901
rect 11360 7793 11389 7839
rect 11435 7793 11464 7839
rect 11360 7731 11464 7793
rect 11360 7685 11389 7731
rect 11435 7685 11464 7731
rect 11360 7623 11464 7685
rect 11360 7577 11389 7623
rect 11435 7577 11464 7623
rect 11360 7515 11464 7577
rect 11360 7469 11389 7515
rect 11435 7469 11464 7515
rect 11360 7407 11464 7469
rect 11360 7361 11389 7407
rect 11435 7361 11464 7407
rect 11360 7299 11464 7361
rect 11360 7253 11389 7299
rect 11435 7253 11464 7299
rect 11360 7191 11464 7253
rect 11360 7145 11389 7191
rect 11435 7145 11464 7191
rect 11360 7132 11464 7145
rect 11584 8273 11688 8286
rect 11584 8227 11613 8273
rect 11659 8227 11688 8273
rect 11584 8164 11688 8227
rect 11584 8118 11613 8164
rect 11659 8118 11688 8164
rect 11584 8055 11688 8118
rect 11584 8009 11613 8055
rect 11659 8009 11688 8055
rect 11584 7947 11688 8009
rect 11584 7901 11613 7947
rect 11659 7901 11688 7947
rect 11584 7839 11688 7901
rect 11584 7793 11613 7839
rect 11659 7793 11688 7839
rect 11584 7731 11688 7793
rect 11584 7685 11613 7731
rect 11659 7685 11688 7731
rect 11584 7623 11688 7685
rect 11584 7577 11613 7623
rect 11659 7577 11688 7623
rect 11584 7515 11688 7577
rect 11584 7469 11613 7515
rect 11659 7469 11688 7515
rect 11584 7407 11688 7469
rect 11584 7361 11613 7407
rect 11659 7361 11688 7407
rect 11584 7299 11688 7361
rect 11584 7253 11613 7299
rect 11659 7253 11688 7299
rect 11584 7191 11688 7253
rect 11584 7145 11613 7191
rect 11659 7145 11688 7191
rect 11584 7132 11688 7145
rect 11808 8273 11912 8286
rect 11808 8227 11837 8273
rect 11883 8227 11912 8273
rect 11808 8164 11912 8227
rect 11808 8118 11837 8164
rect 11883 8118 11912 8164
rect 11808 8055 11912 8118
rect 11808 8009 11837 8055
rect 11883 8009 11912 8055
rect 11808 7947 11912 8009
rect 11808 7901 11837 7947
rect 11883 7901 11912 7947
rect 11808 7839 11912 7901
rect 11808 7793 11837 7839
rect 11883 7793 11912 7839
rect 11808 7731 11912 7793
rect 11808 7685 11837 7731
rect 11883 7685 11912 7731
rect 11808 7623 11912 7685
rect 11808 7577 11837 7623
rect 11883 7577 11912 7623
rect 11808 7515 11912 7577
rect 11808 7469 11837 7515
rect 11883 7469 11912 7515
rect 11808 7407 11912 7469
rect 11808 7361 11837 7407
rect 11883 7361 11912 7407
rect 11808 7299 11912 7361
rect 11808 7253 11837 7299
rect 11883 7253 11912 7299
rect 11808 7191 11912 7253
rect 11808 7145 11837 7191
rect 11883 7145 11912 7191
rect 11808 7132 11912 7145
rect 12032 8273 12120 8286
rect 12032 8227 12061 8273
rect 12107 8227 12120 8273
rect 12032 8164 12120 8227
rect 12032 8118 12061 8164
rect 12107 8118 12120 8164
rect 12032 8055 12120 8118
rect 12032 8009 12061 8055
rect 12107 8009 12120 8055
rect 12032 7947 12120 8009
rect 12032 7901 12061 7947
rect 12107 7901 12120 7947
rect 12032 7839 12120 7901
rect 12032 7793 12061 7839
rect 12107 7793 12120 7839
rect 12032 7731 12120 7793
rect 12032 7685 12061 7731
rect 12107 7685 12120 7731
rect 12032 7623 12120 7685
rect 12032 7577 12061 7623
rect 12107 7577 12120 7623
rect 12032 7515 12120 7577
rect 12032 7469 12061 7515
rect 12107 7469 12120 7515
rect 12032 7407 12120 7469
rect 12032 7361 12061 7407
rect 12107 7361 12120 7407
rect 12032 7299 12120 7361
rect 12032 7253 12061 7299
rect 12107 7253 12120 7299
rect 12032 7191 12120 7253
rect 12032 7145 12061 7191
rect 12107 7145 12120 7191
rect 12032 7132 12120 7145
rect 12338 8273 12426 8286
rect 12338 8227 12351 8273
rect 12397 8227 12426 8273
rect 12338 8164 12426 8227
rect 12338 8118 12351 8164
rect 12397 8118 12426 8164
rect 12338 8055 12426 8118
rect 12338 8009 12351 8055
rect 12397 8009 12426 8055
rect 12338 7947 12426 8009
rect 12338 7901 12351 7947
rect 12397 7901 12426 7947
rect 12338 7839 12426 7901
rect 12338 7793 12351 7839
rect 12397 7793 12426 7839
rect 12338 7731 12426 7793
rect 12338 7685 12351 7731
rect 12397 7685 12426 7731
rect 12338 7623 12426 7685
rect 12338 7577 12351 7623
rect 12397 7577 12426 7623
rect 12338 7515 12426 7577
rect 12338 7469 12351 7515
rect 12397 7469 12426 7515
rect 12338 7407 12426 7469
rect 12338 7361 12351 7407
rect 12397 7361 12426 7407
rect 12338 7299 12426 7361
rect 12338 7253 12351 7299
rect 12397 7253 12426 7299
rect 12338 7191 12426 7253
rect 12338 7145 12351 7191
rect 12397 7145 12426 7191
rect 12338 7132 12426 7145
rect 12546 8273 12650 8286
rect 12546 8227 12575 8273
rect 12621 8227 12650 8273
rect 12546 8164 12650 8227
rect 12546 8118 12575 8164
rect 12621 8118 12650 8164
rect 12546 8055 12650 8118
rect 12546 8009 12575 8055
rect 12621 8009 12650 8055
rect 12546 7947 12650 8009
rect 12546 7901 12575 7947
rect 12621 7901 12650 7947
rect 12546 7839 12650 7901
rect 12546 7793 12575 7839
rect 12621 7793 12650 7839
rect 12546 7731 12650 7793
rect 12546 7685 12575 7731
rect 12621 7685 12650 7731
rect 12546 7623 12650 7685
rect 12546 7577 12575 7623
rect 12621 7577 12650 7623
rect 12546 7515 12650 7577
rect 12546 7469 12575 7515
rect 12621 7469 12650 7515
rect 12546 7407 12650 7469
rect 12546 7361 12575 7407
rect 12621 7361 12650 7407
rect 12546 7299 12650 7361
rect 12546 7253 12575 7299
rect 12621 7253 12650 7299
rect 12546 7191 12650 7253
rect 12546 7145 12575 7191
rect 12621 7145 12650 7191
rect 12546 7132 12650 7145
rect 12770 8273 12874 8286
rect 12770 8227 12799 8273
rect 12845 8227 12874 8273
rect 12770 8164 12874 8227
rect 12770 8118 12799 8164
rect 12845 8118 12874 8164
rect 12770 8055 12874 8118
rect 12770 8009 12799 8055
rect 12845 8009 12874 8055
rect 12770 7947 12874 8009
rect 12770 7901 12799 7947
rect 12845 7901 12874 7947
rect 12770 7839 12874 7901
rect 12770 7793 12799 7839
rect 12845 7793 12874 7839
rect 12770 7731 12874 7793
rect 12770 7685 12799 7731
rect 12845 7685 12874 7731
rect 12770 7623 12874 7685
rect 12770 7577 12799 7623
rect 12845 7577 12874 7623
rect 12770 7515 12874 7577
rect 12770 7469 12799 7515
rect 12845 7469 12874 7515
rect 12770 7407 12874 7469
rect 12770 7361 12799 7407
rect 12845 7361 12874 7407
rect 12770 7299 12874 7361
rect 12770 7253 12799 7299
rect 12845 7253 12874 7299
rect 12770 7191 12874 7253
rect 12770 7145 12799 7191
rect 12845 7145 12874 7191
rect 12770 7132 12874 7145
rect 12994 8273 13098 8286
rect 12994 8227 13023 8273
rect 13069 8227 13098 8273
rect 12994 8164 13098 8227
rect 12994 8118 13023 8164
rect 13069 8118 13098 8164
rect 12994 8055 13098 8118
rect 12994 8009 13023 8055
rect 13069 8009 13098 8055
rect 12994 7947 13098 8009
rect 12994 7901 13023 7947
rect 13069 7901 13098 7947
rect 12994 7839 13098 7901
rect 12994 7793 13023 7839
rect 13069 7793 13098 7839
rect 12994 7731 13098 7793
rect 12994 7685 13023 7731
rect 13069 7685 13098 7731
rect 12994 7623 13098 7685
rect 12994 7577 13023 7623
rect 13069 7577 13098 7623
rect 12994 7515 13098 7577
rect 12994 7469 13023 7515
rect 13069 7469 13098 7515
rect 12994 7407 13098 7469
rect 12994 7361 13023 7407
rect 13069 7361 13098 7407
rect 12994 7299 13098 7361
rect 12994 7253 13023 7299
rect 13069 7253 13098 7299
rect 12994 7191 13098 7253
rect 12994 7145 13023 7191
rect 13069 7145 13098 7191
rect 12994 7132 13098 7145
rect 13218 8273 13322 8286
rect 13218 8227 13247 8273
rect 13293 8227 13322 8273
rect 13218 8164 13322 8227
rect 13218 8118 13247 8164
rect 13293 8118 13322 8164
rect 13218 8055 13322 8118
rect 13218 8009 13247 8055
rect 13293 8009 13322 8055
rect 13218 7947 13322 8009
rect 13218 7901 13247 7947
rect 13293 7901 13322 7947
rect 13218 7839 13322 7901
rect 13218 7793 13247 7839
rect 13293 7793 13322 7839
rect 13218 7731 13322 7793
rect 13218 7685 13247 7731
rect 13293 7685 13322 7731
rect 13218 7623 13322 7685
rect 13218 7577 13247 7623
rect 13293 7577 13322 7623
rect 13218 7515 13322 7577
rect 13218 7469 13247 7515
rect 13293 7469 13322 7515
rect 13218 7407 13322 7469
rect 13218 7361 13247 7407
rect 13293 7361 13322 7407
rect 13218 7299 13322 7361
rect 13218 7253 13247 7299
rect 13293 7253 13322 7299
rect 13218 7191 13322 7253
rect 13218 7145 13247 7191
rect 13293 7145 13322 7191
rect 13218 7132 13322 7145
rect 13442 8273 13546 8286
rect 13442 8227 13471 8273
rect 13517 8227 13546 8273
rect 13442 8164 13546 8227
rect 13442 8118 13471 8164
rect 13517 8118 13546 8164
rect 13442 8055 13546 8118
rect 13442 8009 13471 8055
rect 13517 8009 13546 8055
rect 13442 7947 13546 8009
rect 13442 7901 13471 7947
rect 13517 7901 13546 7947
rect 13442 7839 13546 7901
rect 13442 7793 13471 7839
rect 13517 7793 13546 7839
rect 13442 7731 13546 7793
rect 13442 7685 13471 7731
rect 13517 7685 13546 7731
rect 13442 7623 13546 7685
rect 13442 7577 13471 7623
rect 13517 7577 13546 7623
rect 13442 7515 13546 7577
rect 13442 7469 13471 7515
rect 13517 7469 13546 7515
rect 13442 7407 13546 7469
rect 13442 7361 13471 7407
rect 13517 7361 13546 7407
rect 13442 7299 13546 7361
rect 13442 7253 13471 7299
rect 13517 7253 13546 7299
rect 13442 7191 13546 7253
rect 13442 7145 13471 7191
rect 13517 7145 13546 7191
rect 13442 7132 13546 7145
rect 13666 8273 13754 8286
rect 13666 8227 13695 8273
rect 13741 8227 13754 8273
rect 13666 8164 13754 8227
rect 13666 8118 13695 8164
rect 13741 8118 13754 8164
rect 13666 8055 13754 8118
rect 13666 8009 13695 8055
rect 13741 8009 13754 8055
rect 13666 7947 13754 8009
rect 13666 7901 13695 7947
rect 13741 7901 13754 7947
rect 13666 7839 13754 7901
rect 13666 7793 13695 7839
rect 13741 7793 13754 7839
rect 13666 7731 13754 7793
rect 13666 7685 13695 7731
rect 13741 7685 13754 7731
rect 13666 7623 13754 7685
rect 13666 7577 13695 7623
rect 13741 7577 13754 7623
rect 13666 7515 13754 7577
rect 13666 7469 13695 7515
rect 13741 7469 13754 7515
rect 13666 7407 13754 7469
rect 13666 7361 13695 7407
rect 13741 7361 13754 7407
rect 13666 7299 13754 7361
rect 13666 7253 13695 7299
rect 13741 7253 13754 7299
rect 13666 7191 13754 7253
rect 13666 7145 13695 7191
rect 13741 7145 13754 7191
rect 13666 7132 13754 7145
rect 7437 6406 7525 6419
rect 7437 6360 7450 6406
rect 7496 6360 7525 6406
rect 7437 6300 7525 6360
rect 7437 6254 7450 6300
rect 7496 6254 7525 6300
rect 7437 6194 7525 6254
rect 7437 6148 7450 6194
rect 7496 6148 7525 6194
rect 7437 6088 7525 6148
rect 7437 6042 7450 6088
rect 7496 6042 7525 6088
rect 7437 5982 7525 6042
rect 7437 5936 7450 5982
rect 7496 5936 7525 5982
rect 7437 5876 7525 5936
rect 7437 5830 7450 5876
rect 7496 5830 7525 5876
rect 7437 5770 7525 5830
rect 7437 5724 7450 5770
rect 7496 5724 7525 5770
rect 7437 5664 7525 5724
rect 7437 5618 7450 5664
rect 7496 5618 7525 5664
rect 7437 5558 7525 5618
rect 7437 5512 7450 5558
rect 7496 5512 7525 5558
rect 7437 5451 7525 5512
rect 7437 5405 7450 5451
rect 7496 5405 7525 5451
rect 7437 5344 7525 5405
rect 7437 5298 7450 5344
rect 7496 5298 7525 5344
rect 7437 5285 7525 5298
rect 7645 6406 7749 6419
rect 7645 6360 7674 6406
rect 7720 6360 7749 6406
rect 7645 6300 7749 6360
rect 7645 6254 7674 6300
rect 7720 6254 7749 6300
rect 7645 6194 7749 6254
rect 7645 6148 7674 6194
rect 7720 6148 7749 6194
rect 7645 6088 7749 6148
rect 7645 6042 7674 6088
rect 7720 6042 7749 6088
rect 7645 5982 7749 6042
rect 7645 5936 7674 5982
rect 7720 5936 7749 5982
rect 7645 5876 7749 5936
rect 7645 5830 7674 5876
rect 7720 5830 7749 5876
rect 7645 5770 7749 5830
rect 7645 5724 7674 5770
rect 7720 5724 7749 5770
rect 7645 5664 7749 5724
rect 7645 5618 7674 5664
rect 7720 5618 7749 5664
rect 7645 5558 7749 5618
rect 7645 5512 7674 5558
rect 7720 5512 7749 5558
rect 7645 5451 7749 5512
rect 7645 5405 7674 5451
rect 7720 5405 7749 5451
rect 7645 5344 7749 5405
rect 7645 5298 7674 5344
rect 7720 5298 7749 5344
rect 7645 5285 7749 5298
rect 7869 6406 7973 6419
rect 7869 6360 7898 6406
rect 7944 6360 7973 6406
rect 7869 6300 7973 6360
rect 7869 6254 7898 6300
rect 7944 6254 7973 6300
rect 7869 6194 7973 6254
rect 7869 6148 7898 6194
rect 7944 6148 7973 6194
rect 7869 6088 7973 6148
rect 7869 6042 7898 6088
rect 7944 6042 7973 6088
rect 7869 5982 7973 6042
rect 7869 5936 7898 5982
rect 7944 5936 7973 5982
rect 7869 5876 7973 5936
rect 7869 5830 7898 5876
rect 7944 5830 7973 5876
rect 7869 5770 7973 5830
rect 7869 5724 7898 5770
rect 7944 5724 7973 5770
rect 7869 5664 7973 5724
rect 7869 5618 7898 5664
rect 7944 5618 7973 5664
rect 7869 5558 7973 5618
rect 7869 5512 7898 5558
rect 7944 5512 7973 5558
rect 7869 5451 7973 5512
rect 7869 5405 7898 5451
rect 7944 5405 7973 5451
rect 7869 5344 7973 5405
rect 7869 5298 7898 5344
rect 7944 5298 7973 5344
rect 7869 5285 7973 5298
rect 8093 6406 8197 6419
rect 8093 6360 8122 6406
rect 8168 6360 8197 6406
rect 8093 6300 8197 6360
rect 8093 6254 8122 6300
rect 8168 6254 8197 6300
rect 8093 6194 8197 6254
rect 8093 6148 8122 6194
rect 8168 6148 8197 6194
rect 8093 6088 8197 6148
rect 8093 6042 8122 6088
rect 8168 6042 8197 6088
rect 8093 5982 8197 6042
rect 8093 5936 8122 5982
rect 8168 5936 8197 5982
rect 8093 5876 8197 5936
rect 8093 5830 8122 5876
rect 8168 5830 8197 5876
rect 8093 5770 8197 5830
rect 8093 5724 8122 5770
rect 8168 5724 8197 5770
rect 8093 5664 8197 5724
rect 8093 5618 8122 5664
rect 8168 5618 8197 5664
rect 8093 5558 8197 5618
rect 8093 5512 8122 5558
rect 8168 5512 8197 5558
rect 8093 5451 8197 5512
rect 8093 5405 8122 5451
rect 8168 5405 8197 5451
rect 8093 5344 8197 5405
rect 8093 5298 8122 5344
rect 8168 5298 8197 5344
rect 8093 5285 8197 5298
rect 8317 6406 8421 6419
rect 8317 6360 8346 6406
rect 8392 6360 8421 6406
rect 8317 6300 8421 6360
rect 8317 6254 8346 6300
rect 8392 6254 8421 6300
rect 8317 6194 8421 6254
rect 8317 6148 8346 6194
rect 8392 6148 8421 6194
rect 8317 6088 8421 6148
rect 8317 6042 8346 6088
rect 8392 6042 8421 6088
rect 8317 5982 8421 6042
rect 8317 5936 8346 5982
rect 8392 5936 8421 5982
rect 8317 5876 8421 5936
rect 8317 5830 8346 5876
rect 8392 5830 8421 5876
rect 8317 5770 8421 5830
rect 8317 5724 8346 5770
rect 8392 5724 8421 5770
rect 8317 5664 8421 5724
rect 8317 5618 8346 5664
rect 8392 5618 8421 5664
rect 8317 5558 8421 5618
rect 8317 5512 8346 5558
rect 8392 5512 8421 5558
rect 8317 5451 8421 5512
rect 8317 5405 8346 5451
rect 8392 5405 8421 5451
rect 8317 5344 8421 5405
rect 8317 5298 8346 5344
rect 8392 5298 8421 5344
rect 8317 5285 8421 5298
rect 8541 6406 8645 6419
rect 8541 6360 8570 6406
rect 8616 6360 8645 6406
rect 8541 6300 8645 6360
rect 8541 6254 8570 6300
rect 8616 6254 8645 6300
rect 8541 6194 8645 6254
rect 8541 6148 8570 6194
rect 8616 6148 8645 6194
rect 8541 6088 8645 6148
rect 8541 6042 8570 6088
rect 8616 6042 8645 6088
rect 8541 5982 8645 6042
rect 8541 5936 8570 5982
rect 8616 5936 8645 5982
rect 8541 5876 8645 5936
rect 8541 5830 8570 5876
rect 8616 5830 8645 5876
rect 8541 5770 8645 5830
rect 8541 5724 8570 5770
rect 8616 5724 8645 5770
rect 8541 5664 8645 5724
rect 8541 5618 8570 5664
rect 8616 5618 8645 5664
rect 8541 5558 8645 5618
rect 8541 5512 8570 5558
rect 8616 5512 8645 5558
rect 8541 5451 8645 5512
rect 8541 5405 8570 5451
rect 8616 5405 8645 5451
rect 8541 5344 8645 5405
rect 8541 5298 8570 5344
rect 8616 5298 8645 5344
rect 8541 5285 8645 5298
rect 8765 6406 8853 6419
rect 8765 6360 8794 6406
rect 8840 6360 8853 6406
rect 8765 6300 8853 6360
rect 8765 6254 8794 6300
rect 8840 6254 8853 6300
rect 8765 6194 8853 6254
rect 8765 6148 8794 6194
rect 8840 6148 8853 6194
rect 8765 6088 8853 6148
rect 8765 6042 8794 6088
rect 8840 6042 8853 6088
rect 8765 5982 8853 6042
rect 8765 5936 8794 5982
rect 8840 5936 8853 5982
rect 8765 5876 8853 5936
rect 8765 5830 8794 5876
rect 8840 5830 8853 5876
rect 8765 5770 8853 5830
rect 8765 5724 8794 5770
rect 8840 5724 8853 5770
rect 8765 5664 8853 5724
rect 8765 5618 8794 5664
rect 8840 5618 8853 5664
rect 8765 5558 8853 5618
rect 8765 5512 8794 5558
rect 8840 5512 8853 5558
rect 8765 5451 8853 5512
rect 8765 5405 8794 5451
rect 8840 5405 8853 5451
rect 8765 5344 8853 5405
rect 8765 5298 8794 5344
rect 8840 5298 8853 5344
rect 8765 5285 8853 5298
rect 9070 6406 9158 6419
rect 9070 6360 9083 6406
rect 9129 6360 9158 6406
rect 9070 6300 9158 6360
rect 9070 6254 9083 6300
rect 9129 6254 9158 6300
rect 9070 6194 9158 6254
rect 9070 6148 9083 6194
rect 9129 6148 9158 6194
rect 9070 6088 9158 6148
rect 9070 6042 9083 6088
rect 9129 6042 9158 6088
rect 9070 5982 9158 6042
rect 9070 5936 9083 5982
rect 9129 5936 9158 5982
rect 9070 5876 9158 5936
rect 9070 5830 9083 5876
rect 9129 5830 9158 5876
rect 9070 5770 9158 5830
rect 9070 5724 9083 5770
rect 9129 5724 9158 5770
rect 9070 5664 9158 5724
rect 9070 5618 9083 5664
rect 9129 5618 9158 5664
rect 9070 5558 9158 5618
rect 9070 5512 9083 5558
rect 9129 5512 9158 5558
rect 9070 5451 9158 5512
rect 9070 5405 9083 5451
rect 9129 5405 9158 5451
rect 9070 5344 9158 5405
rect 9070 5298 9083 5344
rect 9129 5298 9158 5344
rect 9070 5285 9158 5298
rect 9278 6406 9382 6419
rect 9278 6360 9307 6406
rect 9353 6360 9382 6406
rect 9278 6300 9382 6360
rect 9278 6254 9307 6300
rect 9353 6254 9382 6300
rect 9278 6194 9382 6254
rect 9278 6148 9307 6194
rect 9353 6148 9382 6194
rect 9278 6088 9382 6148
rect 9278 6042 9307 6088
rect 9353 6042 9382 6088
rect 9278 5982 9382 6042
rect 9278 5936 9307 5982
rect 9353 5936 9382 5982
rect 9278 5876 9382 5936
rect 9278 5830 9307 5876
rect 9353 5830 9382 5876
rect 9278 5770 9382 5830
rect 9278 5724 9307 5770
rect 9353 5724 9382 5770
rect 9278 5664 9382 5724
rect 9278 5618 9307 5664
rect 9353 5618 9382 5664
rect 9278 5558 9382 5618
rect 9278 5512 9307 5558
rect 9353 5512 9382 5558
rect 9278 5451 9382 5512
rect 9278 5405 9307 5451
rect 9353 5405 9382 5451
rect 9278 5344 9382 5405
rect 9278 5298 9307 5344
rect 9353 5298 9382 5344
rect 9278 5285 9382 5298
rect 9502 6406 9606 6419
rect 9502 6360 9531 6406
rect 9577 6360 9606 6406
rect 9502 6300 9606 6360
rect 9502 6254 9531 6300
rect 9577 6254 9606 6300
rect 9502 6194 9606 6254
rect 9502 6148 9531 6194
rect 9577 6148 9606 6194
rect 9502 6088 9606 6148
rect 9502 6042 9531 6088
rect 9577 6042 9606 6088
rect 9502 5982 9606 6042
rect 9502 5936 9531 5982
rect 9577 5936 9606 5982
rect 9502 5876 9606 5936
rect 9502 5830 9531 5876
rect 9577 5830 9606 5876
rect 9502 5770 9606 5830
rect 9502 5724 9531 5770
rect 9577 5724 9606 5770
rect 9502 5664 9606 5724
rect 9502 5618 9531 5664
rect 9577 5618 9606 5664
rect 9502 5558 9606 5618
rect 9502 5512 9531 5558
rect 9577 5512 9606 5558
rect 9502 5451 9606 5512
rect 9502 5405 9531 5451
rect 9577 5405 9606 5451
rect 9502 5344 9606 5405
rect 9502 5298 9531 5344
rect 9577 5298 9606 5344
rect 9502 5285 9606 5298
rect 9726 6406 9830 6419
rect 9726 6360 9755 6406
rect 9801 6360 9830 6406
rect 9726 6300 9830 6360
rect 9726 6254 9755 6300
rect 9801 6254 9830 6300
rect 9726 6194 9830 6254
rect 9726 6148 9755 6194
rect 9801 6148 9830 6194
rect 9726 6088 9830 6148
rect 9726 6042 9755 6088
rect 9801 6042 9830 6088
rect 9726 5982 9830 6042
rect 9726 5936 9755 5982
rect 9801 5936 9830 5982
rect 9726 5876 9830 5936
rect 9726 5830 9755 5876
rect 9801 5830 9830 5876
rect 9726 5770 9830 5830
rect 9726 5724 9755 5770
rect 9801 5724 9830 5770
rect 9726 5664 9830 5724
rect 9726 5618 9755 5664
rect 9801 5618 9830 5664
rect 9726 5558 9830 5618
rect 9726 5512 9755 5558
rect 9801 5512 9830 5558
rect 9726 5451 9830 5512
rect 9726 5405 9755 5451
rect 9801 5405 9830 5451
rect 9726 5344 9830 5405
rect 9726 5298 9755 5344
rect 9801 5298 9830 5344
rect 9726 5285 9830 5298
rect 9950 6406 10054 6419
rect 9950 6360 9979 6406
rect 10025 6360 10054 6406
rect 9950 6300 10054 6360
rect 9950 6254 9979 6300
rect 10025 6254 10054 6300
rect 9950 6194 10054 6254
rect 9950 6148 9979 6194
rect 10025 6148 10054 6194
rect 9950 6088 10054 6148
rect 9950 6042 9979 6088
rect 10025 6042 10054 6088
rect 9950 5982 10054 6042
rect 9950 5936 9979 5982
rect 10025 5936 10054 5982
rect 9950 5876 10054 5936
rect 9950 5830 9979 5876
rect 10025 5830 10054 5876
rect 9950 5770 10054 5830
rect 9950 5724 9979 5770
rect 10025 5724 10054 5770
rect 9950 5664 10054 5724
rect 9950 5618 9979 5664
rect 10025 5618 10054 5664
rect 9950 5558 10054 5618
rect 9950 5512 9979 5558
rect 10025 5512 10054 5558
rect 9950 5451 10054 5512
rect 9950 5405 9979 5451
rect 10025 5405 10054 5451
rect 9950 5344 10054 5405
rect 9950 5298 9979 5344
rect 10025 5298 10054 5344
rect 9950 5285 10054 5298
rect 10174 6406 10278 6419
rect 10174 6360 10203 6406
rect 10249 6360 10278 6406
rect 10174 6300 10278 6360
rect 10174 6254 10203 6300
rect 10249 6254 10278 6300
rect 10174 6194 10278 6254
rect 10174 6148 10203 6194
rect 10249 6148 10278 6194
rect 10174 6088 10278 6148
rect 10174 6042 10203 6088
rect 10249 6042 10278 6088
rect 10174 5982 10278 6042
rect 10174 5936 10203 5982
rect 10249 5936 10278 5982
rect 10174 5876 10278 5936
rect 10174 5830 10203 5876
rect 10249 5830 10278 5876
rect 10174 5770 10278 5830
rect 10174 5724 10203 5770
rect 10249 5724 10278 5770
rect 10174 5664 10278 5724
rect 10174 5618 10203 5664
rect 10249 5618 10278 5664
rect 10174 5558 10278 5618
rect 10174 5512 10203 5558
rect 10249 5512 10278 5558
rect 10174 5451 10278 5512
rect 10174 5405 10203 5451
rect 10249 5405 10278 5451
rect 10174 5344 10278 5405
rect 10174 5298 10203 5344
rect 10249 5298 10278 5344
rect 10174 5285 10278 5298
rect 10398 6406 10486 6419
rect 10398 6360 10427 6406
rect 10473 6360 10486 6406
rect 10398 6300 10486 6360
rect 10398 6254 10427 6300
rect 10473 6254 10486 6300
rect 10398 6194 10486 6254
rect 10398 6148 10427 6194
rect 10473 6148 10486 6194
rect 10398 6088 10486 6148
rect 10398 6042 10427 6088
rect 10473 6042 10486 6088
rect 10398 5982 10486 6042
rect 10398 5936 10427 5982
rect 10473 5936 10486 5982
rect 10398 5876 10486 5936
rect 10398 5830 10427 5876
rect 10473 5830 10486 5876
rect 10398 5770 10486 5830
rect 10398 5724 10427 5770
rect 10473 5724 10486 5770
rect 10398 5664 10486 5724
rect 10398 5618 10427 5664
rect 10473 5618 10486 5664
rect 10398 5558 10486 5618
rect 10398 5512 10427 5558
rect 10473 5512 10486 5558
rect 10398 5451 10486 5512
rect 10398 5405 10427 5451
rect 10473 5405 10486 5451
rect 10398 5344 10486 5405
rect 10398 5298 10427 5344
rect 10473 5298 10486 5344
rect 10398 5285 10486 5298
rect 10704 6406 10792 6419
rect 10704 6360 10717 6406
rect 10763 6360 10792 6406
rect 10704 6300 10792 6360
rect 10704 6254 10717 6300
rect 10763 6254 10792 6300
rect 10704 6194 10792 6254
rect 10704 6148 10717 6194
rect 10763 6148 10792 6194
rect 10704 6088 10792 6148
rect 10704 6042 10717 6088
rect 10763 6042 10792 6088
rect 10704 5982 10792 6042
rect 10704 5936 10717 5982
rect 10763 5936 10792 5982
rect 10704 5876 10792 5936
rect 10704 5830 10717 5876
rect 10763 5830 10792 5876
rect 10704 5770 10792 5830
rect 10704 5724 10717 5770
rect 10763 5724 10792 5770
rect 10704 5664 10792 5724
rect 10704 5618 10717 5664
rect 10763 5618 10792 5664
rect 10704 5558 10792 5618
rect 10704 5512 10717 5558
rect 10763 5512 10792 5558
rect 10704 5451 10792 5512
rect 10704 5405 10717 5451
rect 10763 5405 10792 5451
rect 10704 5344 10792 5405
rect 10704 5298 10717 5344
rect 10763 5298 10792 5344
rect 10704 5285 10792 5298
rect 10912 6406 11016 6419
rect 10912 6360 10941 6406
rect 10987 6360 11016 6406
rect 10912 6300 11016 6360
rect 10912 6254 10941 6300
rect 10987 6254 11016 6300
rect 10912 6194 11016 6254
rect 10912 6148 10941 6194
rect 10987 6148 11016 6194
rect 10912 6088 11016 6148
rect 10912 6042 10941 6088
rect 10987 6042 11016 6088
rect 10912 5982 11016 6042
rect 10912 5936 10941 5982
rect 10987 5936 11016 5982
rect 10912 5876 11016 5936
rect 10912 5830 10941 5876
rect 10987 5830 11016 5876
rect 10912 5770 11016 5830
rect 10912 5724 10941 5770
rect 10987 5724 11016 5770
rect 10912 5664 11016 5724
rect 10912 5618 10941 5664
rect 10987 5618 11016 5664
rect 10912 5558 11016 5618
rect 10912 5512 10941 5558
rect 10987 5512 11016 5558
rect 10912 5451 11016 5512
rect 10912 5405 10941 5451
rect 10987 5405 11016 5451
rect 10912 5344 11016 5405
rect 10912 5298 10941 5344
rect 10987 5298 11016 5344
rect 10912 5285 11016 5298
rect 11136 6406 11240 6419
rect 11136 6360 11165 6406
rect 11211 6360 11240 6406
rect 11136 6300 11240 6360
rect 11136 6254 11165 6300
rect 11211 6254 11240 6300
rect 11136 6194 11240 6254
rect 11136 6148 11165 6194
rect 11211 6148 11240 6194
rect 11136 6088 11240 6148
rect 11136 6042 11165 6088
rect 11211 6042 11240 6088
rect 11136 5982 11240 6042
rect 11136 5936 11165 5982
rect 11211 5936 11240 5982
rect 11136 5876 11240 5936
rect 11136 5830 11165 5876
rect 11211 5830 11240 5876
rect 11136 5770 11240 5830
rect 11136 5724 11165 5770
rect 11211 5724 11240 5770
rect 11136 5664 11240 5724
rect 11136 5618 11165 5664
rect 11211 5618 11240 5664
rect 11136 5558 11240 5618
rect 11136 5512 11165 5558
rect 11211 5512 11240 5558
rect 11136 5451 11240 5512
rect 11136 5405 11165 5451
rect 11211 5405 11240 5451
rect 11136 5344 11240 5405
rect 11136 5298 11165 5344
rect 11211 5298 11240 5344
rect 11136 5285 11240 5298
rect 11360 6406 11464 6419
rect 11360 6360 11389 6406
rect 11435 6360 11464 6406
rect 11360 6300 11464 6360
rect 11360 6254 11389 6300
rect 11435 6254 11464 6300
rect 11360 6194 11464 6254
rect 11360 6148 11389 6194
rect 11435 6148 11464 6194
rect 11360 6088 11464 6148
rect 11360 6042 11389 6088
rect 11435 6042 11464 6088
rect 11360 5982 11464 6042
rect 11360 5936 11389 5982
rect 11435 5936 11464 5982
rect 11360 5876 11464 5936
rect 11360 5830 11389 5876
rect 11435 5830 11464 5876
rect 11360 5770 11464 5830
rect 11360 5724 11389 5770
rect 11435 5724 11464 5770
rect 11360 5664 11464 5724
rect 11360 5618 11389 5664
rect 11435 5618 11464 5664
rect 11360 5558 11464 5618
rect 11360 5512 11389 5558
rect 11435 5512 11464 5558
rect 11360 5451 11464 5512
rect 11360 5405 11389 5451
rect 11435 5405 11464 5451
rect 11360 5344 11464 5405
rect 11360 5298 11389 5344
rect 11435 5298 11464 5344
rect 11360 5285 11464 5298
rect 11584 6406 11688 6419
rect 11584 6360 11613 6406
rect 11659 6360 11688 6406
rect 11584 6300 11688 6360
rect 11584 6254 11613 6300
rect 11659 6254 11688 6300
rect 11584 6194 11688 6254
rect 11584 6148 11613 6194
rect 11659 6148 11688 6194
rect 11584 6088 11688 6148
rect 11584 6042 11613 6088
rect 11659 6042 11688 6088
rect 11584 5982 11688 6042
rect 11584 5936 11613 5982
rect 11659 5936 11688 5982
rect 11584 5876 11688 5936
rect 11584 5830 11613 5876
rect 11659 5830 11688 5876
rect 11584 5770 11688 5830
rect 11584 5724 11613 5770
rect 11659 5724 11688 5770
rect 11584 5664 11688 5724
rect 11584 5618 11613 5664
rect 11659 5618 11688 5664
rect 11584 5558 11688 5618
rect 11584 5512 11613 5558
rect 11659 5512 11688 5558
rect 11584 5451 11688 5512
rect 11584 5405 11613 5451
rect 11659 5405 11688 5451
rect 11584 5344 11688 5405
rect 11584 5298 11613 5344
rect 11659 5298 11688 5344
rect 11584 5285 11688 5298
rect 11808 6406 11912 6419
rect 11808 6360 11837 6406
rect 11883 6360 11912 6406
rect 11808 6300 11912 6360
rect 11808 6254 11837 6300
rect 11883 6254 11912 6300
rect 11808 6194 11912 6254
rect 11808 6148 11837 6194
rect 11883 6148 11912 6194
rect 11808 6088 11912 6148
rect 11808 6042 11837 6088
rect 11883 6042 11912 6088
rect 11808 5982 11912 6042
rect 11808 5936 11837 5982
rect 11883 5936 11912 5982
rect 11808 5876 11912 5936
rect 11808 5830 11837 5876
rect 11883 5830 11912 5876
rect 11808 5770 11912 5830
rect 11808 5724 11837 5770
rect 11883 5724 11912 5770
rect 11808 5664 11912 5724
rect 11808 5618 11837 5664
rect 11883 5618 11912 5664
rect 11808 5558 11912 5618
rect 11808 5512 11837 5558
rect 11883 5512 11912 5558
rect 11808 5451 11912 5512
rect 11808 5405 11837 5451
rect 11883 5405 11912 5451
rect 11808 5344 11912 5405
rect 11808 5298 11837 5344
rect 11883 5298 11912 5344
rect 11808 5285 11912 5298
rect 12032 6406 12120 6419
rect 12032 6360 12061 6406
rect 12107 6360 12120 6406
rect 12032 6300 12120 6360
rect 12032 6254 12061 6300
rect 12107 6254 12120 6300
rect 12032 6194 12120 6254
rect 12032 6148 12061 6194
rect 12107 6148 12120 6194
rect 12032 6088 12120 6148
rect 12032 6042 12061 6088
rect 12107 6042 12120 6088
rect 12032 5982 12120 6042
rect 12032 5936 12061 5982
rect 12107 5936 12120 5982
rect 12032 5876 12120 5936
rect 12032 5830 12061 5876
rect 12107 5830 12120 5876
rect 12032 5770 12120 5830
rect 12032 5724 12061 5770
rect 12107 5724 12120 5770
rect 12032 5664 12120 5724
rect 12032 5618 12061 5664
rect 12107 5618 12120 5664
rect 12032 5558 12120 5618
rect 12032 5512 12061 5558
rect 12107 5512 12120 5558
rect 12032 5451 12120 5512
rect 12032 5405 12061 5451
rect 12107 5405 12120 5451
rect 12032 5344 12120 5405
rect 12032 5298 12061 5344
rect 12107 5298 12120 5344
rect 12032 5285 12120 5298
rect 12338 6406 12426 6419
rect 12338 6360 12351 6406
rect 12397 6360 12426 6406
rect 12338 6300 12426 6360
rect 12338 6254 12351 6300
rect 12397 6254 12426 6300
rect 12338 6194 12426 6254
rect 12338 6148 12351 6194
rect 12397 6148 12426 6194
rect 12338 6088 12426 6148
rect 12338 6042 12351 6088
rect 12397 6042 12426 6088
rect 12338 5982 12426 6042
rect 12338 5936 12351 5982
rect 12397 5936 12426 5982
rect 12338 5876 12426 5936
rect 12338 5830 12351 5876
rect 12397 5830 12426 5876
rect 12338 5770 12426 5830
rect 12338 5724 12351 5770
rect 12397 5724 12426 5770
rect 12338 5664 12426 5724
rect 12338 5618 12351 5664
rect 12397 5618 12426 5664
rect 12338 5558 12426 5618
rect 12338 5512 12351 5558
rect 12397 5512 12426 5558
rect 12338 5451 12426 5512
rect 12338 5405 12351 5451
rect 12397 5405 12426 5451
rect 12338 5344 12426 5405
rect 12338 5298 12351 5344
rect 12397 5298 12426 5344
rect 12338 5285 12426 5298
rect 12546 6406 12650 6419
rect 12546 6360 12575 6406
rect 12621 6360 12650 6406
rect 12546 6300 12650 6360
rect 12546 6254 12575 6300
rect 12621 6254 12650 6300
rect 12546 6194 12650 6254
rect 12546 6148 12575 6194
rect 12621 6148 12650 6194
rect 12546 6088 12650 6148
rect 12546 6042 12575 6088
rect 12621 6042 12650 6088
rect 12546 5982 12650 6042
rect 12546 5936 12575 5982
rect 12621 5936 12650 5982
rect 12546 5876 12650 5936
rect 12546 5830 12575 5876
rect 12621 5830 12650 5876
rect 12546 5770 12650 5830
rect 12546 5724 12575 5770
rect 12621 5724 12650 5770
rect 12546 5664 12650 5724
rect 12546 5618 12575 5664
rect 12621 5618 12650 5664
rect 12546 5558 12650 5618
rect 12546 5512 12575 5558
rect 12621 5512 12650 5558
rect 12546 5451 12650 5512
rect 12546 5405 12575 5451
rect 12621 5405 12650 5451
rect 12546 5344 12650 5405
rect 12546 5298 12575 5344
rect 12621 5298 12650 5344
rect 12546 5285 12650 5298
rect 12770 6406 12874 6419
rect 12770 6360 12799 6406
rect 12845 6360 12874 6406
rect 12770 6300 12874 6360
rect 12770 6254 12799 6300
rect 12845 6254 12874 6300
rect 12770 6194 12874 6254
rect 12770 6148 12799 6194
rect 12845 6148 12874 6194
rect 12770 6088 12874 6148
rect 12770 6042 12799 6088
rect 12845 6042 12874 6088
rect 12770 5982 12874 6042
rect 12770 5936 12799 5982
rect 12845 5936 12874 5982
rect 12770 5876 12874 5936
rect 12770 5830 12799 5876
rect 12845 5830 12874 5876
rect 12770 5770 12874 5830
rect 12770 5724 12799 5770
rect 12845 5724 12874 5770
rect 12770 5664 12874 5724
rect 12770 5618 12799 5664
rect 12845 5618 12874 5664
rect 12770 5558 12874 5618
rect 12770 5512 12799 5558
rect 12845 5512 12874 5558
rect 12770 5451 12874 5512
rect 12770 5405 12799 5451
rect 12845 5405 12874 5451
rect 12770 5344 12874 5405
rect 12770 5298 12799 5344
rect 12845 5298 12874 5344
rect 12770 5285 12874 5298
rect 12994 6406 13098 6419
rect 12994 6360 13023 6406
rect 13069 6360 13098 6406
rect 12994 6300 13098 6360
rect 12994 6254 13023 6300
rect 13069 6254 13098 6300
rect 12994 6194 13098 6254
rect 12994 6148 13023 6194
rect 13069 6148 13098 6194
rect 12994 6088 13098 6148
rect 12994 6042 13023 6088
rect 13069 6042 13098 6088
rect 12994 5982 13098 6042
rect 12994 5936 13023 5982
rect 13069 5936 13098 5982
rect 12994 5876 13098 5936
rect 12994 5830 13023 5876
rect 13069 5830 13098 5876
rect 12994 5770 13098 5830
rect 12994 5724 13023 5770
rect 13069 5724 13098 5770
rect 12994 5664 13098 5724
rect 12994 5618 13023 5664
rect 13069 5618 13098 5664
rect 12994 5558 13098 5618
rect 12994 5512 13023 5558
rect 13069 5512 13098 5558
rect 12994 5451 13098 5512
rect 12994 5405 13023 5451
rect 13069 5405 13098 5451
rect 12994 5344 13098 5405
rect 12994 5298 13023 5344
rect 13069 5298 13098 5344
rect 12994 5285 13098 5298
rect 13218 6406 13322 6419
rect 13218 6360 13247 6406
rect 13293 6360 13322 6406
rect 13218 6300 13322 6360
rect 13218 6254 13247 6300
rect 13293 6254 13322 6300
rect 13218 6194 13322 6254
rect 13218 6148 13247 6194
rect 13293 6148 13322 6194
rect 13218 6088 13322 6148
rect 13218 6042 13247 6088
rect 13293 6042 13322 6088
rect 13218 5982 13322 6042
rect 13218 5936 13247 5982
rect 13293 5936 13322 5982
rect 13218 5876 13322 5936
rect 13218 5830 13247 5876
rect 13293 5830 13322 5876
rect 13218 5770 13322 5830
rect 13218 5724 13247 5770
rect 13293 5724 13322 5770
rect 13218 5664 13322 5724
rect 13218 5618 13247 5664
rect 13293 5618 13322 5664
rect 13218 5558 13322 5618
rect 13218 5512 13247 5558
rect 13293 5512 13322 5558
rect 13218 5451 13322 5512
rect 13218 5405 13247 5451
rect 13293 5405 13322 5451
rect 13218 5344 13322 5405
rect 13218 5298 13247 5344
rect 13293 5298 13322 5344
rect 13218 5285 13322 5298
rect 13442 6406 13546 6419
rect 13442 6360 13471 6406
rect 13517 6360 13546 6406
rect 13442 6300 13546 6360
rect 13442 6254 13471 6300
rect 13517 6254 13546 6300
rect 13442 6194 13546 6254
rect 13442 6148 13471 6194
rect 13517 6148 13546 6194
rect 13442 6088 13546 6148
rect 13442 6042 13471 6088
rect 13517 6042 13546 6088
rect 13442 5982 13546 6042
rect 13442 5936 13471 5982
rect 13517 5936 13546 5982
rect 13442 5876 13546 5936
rect 13442 5830 13471 5876
rect 13517 5830 13546 5876
rect 13442 5770 13546 5830
rect 13442 5724 13471 5770
rect 13517 5724 13546 5770
rect 13442 5664 13546 5724
rect 13442 5618 13471 5664
rect 13517 5618 13546 5664
rect 13442 5558 13546 5618
rect 13442 5512 13471 5558
rect 13517 5512 13546 5558
rect 13442 5451 13546 5512
rect 13442 5405 13471 5451
rect 13517 5405 13546 5451
rect 13442 5344 13546 5405
rect 13442 5298 13471 5344
rect 13517 5298 13546 5344
rect 13442 5285 13546 5298
rect 13666 6406 13754 6419
rect 13666 6360 13695 6406
rect 13741 6360 13754 6406
rect 13666 6300 13754 6360
rect 13666 6254 13695 6300
rect 13741 6254 13754 6300
rect 13666 6194 13754 6254
rect 13666 6148 13695 6194
rect 13741 6148 13754 6194
rect 13666 6088 13754 6148
rect 13666 6042 13695 6088
rect 13741 6042 13754 6088
rect 13666 5982 13754 6042
rect 13666 5936 13695 5982
rect 13741 5936 13754 5982
rect 13666 5876 13754 5936
rect 13666 5830 13695 5876
rect 13741 5830 13754 5876
rect 13666 5770 13754 5830
rect 13666 5724 13695 5770
rect 13741 5724 13754 5770
rect 13666 5664 13754 5724
rect 13666 5618 13695 5664
rect 13741 5618 13754 5664
rect 13666 5558 13754 5618
rect 13666 5512 13695 5558
rect 13741 5512 13754 5558
rect 13666 5451 13754 5512
rect 13666 5405 13695 5451
rect 13741 5405 13754 5451
rect 13666 5344 13754 5405
rect 13666 5298 13695 5344
rect 13741 5298 13754 5344
rect 13666 5285 13754 5298
rect 6712 5255 6800 5268
rect 7719 1170 7807 1183
rect 7719 1124 7732 1170
rect 7778 1124 7807 1170
rect 7719 1035 7807 1124
rect 7719 989 7732 1035
rect 7778 989 7807 1035
rect 7719 900 7807 989
rect 7719 854 7732 900
rect 7778 854 7807 900
rect 7719 841 7807 854
rect 7927 1170 8031 1183
rect 7927 1124 7956 1170
rect 8002 1124 8031 1170
rect 7927 1035 8031 1124
rect 7927 989 7956 1035
rect 8002 989 8031 1035
rect 7927 900 8031 989
rect 7927 854 7956 900
rect 8002 854 8031 900
rect 7927 841 8031 854
rect 8151 1170 8239 1183
rect 8151 1124 8180 1170
rect 8226 1124 8239 1170
rect 8151 1035 8239 1124
rect 8151 989 8180 1035
rect 8226 989 8239 1035
rect 8151 900 8239 989
rect 8151 854 8180 900
rect 8226 854 8239 900
rect 8151 841 8239 854
rect 8717 1123 8836 1282
rect 8717 1077 8761 1123
rect 8807 1077 8836 1123
rect 8717 919 8836 1077
rect 8717 873 8761 919
rect 8807 873 8836 919
rect 8717 827 8836 873
rect 8956 827 9060 1282
rect 9180 1123 9284 1282
rect 9180 1077 9209 1123
rect 9255 1077 9284 1123
rect 9180 919 9284 1077
rect 9180 873 9209 919
rect 9255 873 9284 919
rect 9180 827 9284 873
rect 9404 827 9508 1282
rect 9628 1123 9746 1282
rect 9628 1077 9657 1123
rect 9703 1077 9746 1123
rect 9628 919 9746 1077
rect 9628 873 9657 919
rect 9703 873 9746 919
rect 9628 827 9746 873
<< mvndiffc >>
rect 1659 28594 1705 28640
rect 1659 28489 1705 28535
rect 1659 28384 1705 28430
rect 1659 28279 1705 28325
rect 1659 28174 1705 28220
rect 1659 28070 1705 28116
rect 1659 27966 1705 28012
rect 1659 27862 1705 27908
rect 1659 27758 1705 27804
rect 1883 28594 1929 28640
rect 1883 28489 1929 28535
rect 1883 28384 1929 28430
rect 1883 28279 1929 28325
rect 1883 28174 1929 28220
rect 1883 28070 1929 28116
rect 1883 27966 1929 28012
rect 1883 27862 1929 27908
rect 1883 27758 1929 27804
rect 2107 28594 2153 28640
rect 2107 28489 2153 28535
rect 2107 28384 2153 28430
rect 2107 28279 2153 28325
rect 2107 28174 2153 28220
rect 2107 28070 2153 28116
rect 2107 27966 2153 28012
rect 2107 27862 2153 27908
rect 2107 27758 2153 27804
rect 2331 28594 2377 28640
rect 2331 28489 2377 28535
rect 2331 28384 2377 28430
rect 2331 28279 2377 28325
rect 2331 28174 2377 28220
rect 2331 28070 2377 28116
rect 2331 27966 2377 28012
rect 2331 27862 2377 27908
rect 2331 27758 2377 27804
rect 2555 28594 2601 28640
rect 2555 28489 2601 28535
rect 2555 28384 2601 28430
rect 2555 28279 2601 28325
rect 2555 28174 2601 28220
rect 2555 28070 2601 28116
rect 2555 27966 2601 28012
rect 2555 27862 2601 27908
rect 2555 27758 2601 27804
rect 2779 28594 2825 28640
rect 2779 28489 2825 28535
rect 2779 28384 2825 28430
rect 2779 28279 2825 28325
rect 2779 28174 2825 28220
rect 2779 28070 2825 28116
rect 2779 27966 2825 28012
rect 2779 27862 2825 27908
rect 2779 27758 2825 27804
rect 3003 28594 3049 28640
rect 3003 28489 3049 28535
rect 3003 28384 3049 28430
rect 3003 28279 3049 28325
rect 3003 28174 3049 28220
rect 3003 28070 3049 28116
rect 3003 27966 3049 28012
rect 3003 27862 3049 27908
rect 3003 27758 3049 27804
rect 3227 28594 3273 28640
rect 3227 28489 3273 28535
rect 3227 28384 3273 28430
rect 3227 28279 3273 28325
rect 3227 28174 3273 28220
rect 3227 28070 3273 28116
rect 3227 27966 3273 28012
rect 3227 27862 3273 27908
rect 3227 27758 3273 27804
rect 3451 28594 3497 28640
rect 3451 28489 3497 28535
rect 3451 28384 3497 28430
rect 3451 28279 3497 28325
rect 3451 28174 3497 28220
rect 3451 28070 3497 28116
rect 3451 27966 3497 28012
rect 3451 27862 3497 27908
rect 3451 27758 3497 27804
rect 3675 28594 3721 28640
rect 3675 28489 3721 28535
rect 3675 28384 3721 28430
rect 3675 28279 3721 28325
rect 3675 28174 3721 28220
rect 3675 28070 3721 28116
rect 3675 27966 3721 28012
rect 3675 27862 3721 27908
rect 3675 27758 3721 27804
rect 3899 28594 3945 28640
rect 3899 28489 3945 28535
rect 3899 28384 3945 28430
rect 3899 28279 3945 28325
rect 3899 28174 3945 28220
rect 3899 28070 3945 28116
rect 3899 27966 3945 28012
rect 3899 27862 3945 27908
rect 3899 27758 3945 27804
rect 4123 28594 4169 28640
rect 4123 28489 4169 28535
rect 4123 28384 4169 28430
rect 4123 28279 4169 28325
rect 4123 28174 4169 28220
rect 4123 28070 4169 28116
rect 4123 27966 4169 28012
rect 4123 27862 4169 27908
rect 4123 27758 4169 27804
rect 4347 28594 4393 28640
rect 4347 28489 4393 28535
rect 4347 28384 4393 28430
rect 4347 28279 4393 28325
rect 4347 28174 4393 28220
rect 4347 28070 4393 28116
rect 4347 27966 4393 28012
rect 4347 27862 4393 27908
rect 4347 27758 4393 27804
rect 4571 28594 4617 28640
rect 4571 28489 4617 28535
rect 4571 28384 4617 28430
rect 4571 28279 4617 28325
rect 4571 28174 4617 28220
rect 4571 28070 4617 28116
rect 4571 27966 4617 28012
rect 4571 27862 4617 27908
rect 4571 27758 4617 27804
rect 4795 28594 4841 28640
rect 4795 28489 4841 28535
rect 4795 28384 4841 28430
rect 4795 28279 4841 28325
rect 4795 28174 4841 28220
rect 4795 28070 4841 28116
rect 4795 27966 4841 28012
rect 4795 27862 4841 27908
rect 4795 27758 4841 27804
rect 5019 28594 5065 28640
rect 5019 28489 5065 28535
rect 5019 28384 5065 28430
rect 5019 28279 5065 28325
rect 5019 28174 5065 28220
rect 5019 28070 5065 28116
rect 5019 27966 5065 28012
rect 5019 27862 5065 27908
rect 5019 27758 5065 27804
rect 5243 28594 5289 28640
rect 5243 28489 5289 28535
rect 5243 28384 5289 28430
rect 5243 28279 5289 28325
rect 5243 28174 5289 28220
rect 9038 28594 9084 28640
rect 9038 28489 9084 28535
rect 9038 28384 9084 28430
rect 9038 28279 9084 28325
rect 9038 28174 9084 28220
rect 5243 28070 5289 28116
rect 5243 27966 5289 28012
rect 5243 27862 5289 27908
rect 5933 27834 5979 28082
rect 6157 27834 6203 28082
rect 6381 27834 6427 28082
rect 9038 28070 9084 28116
rect 5243 27758 5289 27804
rect 7527 27950 7573 27996
rect 7527 27830 7573 27876
rect 7751 27950 7797 27996
rect 7751 27830 7797 27876
rect 9038 27966 9084 28012
rect 9038 27862 9084 27908
rect 9038 27758 9084 27804
rect 9262 28594 9308 28640
rect 9262 28489 9308 28535
rect 9262 28384 9308 28430
rect 9262 28279 9308 28325
rect 9262 28174 9308 28220
rect 9262 28070 9308 28116
rect 9262 27966 9308 28012
rect 9262 27862 9308 27908
rect 9262 27758 9308 27804
rect 9486 28594 9532 28640
rect 9486 28489 9532 28535
rect 9486 28384 9532 28430
rect 9486 28279 9532 28325
rect 9486 28174 9532 28220
rect 9486 28070 9532 28116
rect 9486 27966 9532 28012
rect 9486 27862 9532 27908
rect 9486 27758 9532 27804
rect 9710 28594 9756 28640
rect 9710 28489 9756 28535
rect 9710 28384 9756 28430
rect 9710 28279 9756 28325
rect 9710 28174 9756 28220
rect 9710 28070 9756 28116
rect 9710 27966 9756 28012
rect 9710 27862 9756 27908
rect 9710 27758 9756 27804
rect 9934 28594 9980 28640
rect 9934 28489 9980 28535
rect 9934 28384 9980 28430
rect 9934 28279 9980 28325
rect 9934 28174 9980 28220
rect 9934 28070 9980 28116
rect 9934 27966 9980 28012
rect 9934 27862 9980 27908
rect 9934 27758 9980 27804
rect 10158 28594 10204 28640
rect 10158 28489 10204 28535
rect 10158 28384 10204 28430
rect 10158 28279 10204 28325
rect 10158 28174 10204 28220
rect 10158 28070 10204 28116
rect 10158 27966 10204 28012
rect 10158 27862 10204 27908
rect 10158 27758 10204 27804
rect 10382 28594 10428 28640
rect 10382 28489 10428 28535
rect 10382 28384 10428 28430
rect 10382 28279 10428 28325
rect 10382 28174 10428 28220
rect 10382 28070 10428 28116
rect 10382 27966 10428 28012
rect 10382 27862 10428 27908
rect 10382 27758 10428 27804
rect 10606 28594 10652 28640
rect 10606 28489 10652 28535
rect 10606 28384 10652 28430
rect 10606 28279 10652 28325
rect 10606 28174 10652 28220
rect 10606 28070 10652 28116
rect 10606 27966 10652 28012
rect 10606 27862 10652 27908
rect 10606 27758 10652 27804
rect 10830 28594 10876 28640
rect 10830 28489 10876 28535
rect 10830 28384 10876 28430
rect 10830 28279 10876 28325
rect 10830 28174 10876 28220
rect 10830 28070 10876 28116
rect 10830 27966 10876 28012
rect 10830 27862 10876 27908
rect 10830 27758 10876 27804
rect 11054 28594 11100 28640
rect 11054 28489 11100 28535
rect 11054 28384 11100 28430
rect 11054 28279 11100 28325
rect 11054 28174 11100 28220
rect 11054 28070 11100 28116
rect 11054 27966 11100 28012
rect 11054 27862 11100 27908
rect 11054 27758 11100 27804
rect 11278 28594 11324 28640
rect 11278 28489 11324 28535
rect 11278 28384 11324 28430
rect 11278 28279 11324 28325
rect 11278 28174 11324 28220
rect 11278 28070 11324 28116
rect 11278 27966 11324 28012
rect 11278 27862 11324 27908
rect 11278 27758 11324 27804
rect 11502 28594 11548 28640
rect 11502 28489 11548 28535
rect 11502 28384 11548 28430
rect 11502 28279 11548 28325
rect 11502 28174 11548 28220
rect 11502 28070 11548 28116
rect 11502 27966 11548 28012
rect 11502 27862 11548 27908
rect 11502 27758 11548 27804
rect 11726 28594 11772 28640
rect 11726 28489 11772 28535
rect 11726 28384 11772 28430
rect 11726 28279 11772 28325
rect 11726 28174 11772 28220
rect 11726 28070 11772 28116
rect 11726 27966 11772 28012
rect 11726 27862 11772 27908
rect 11726 27758 11772 27804
rect 11950 28594 11996 28640
rect 11950 28489 11996 28535
rect 11950 28384 11996 28430
rect 11950 28279 11996 28325
rect 11950 28174 11996 28220
rect 11950 28070 11996 28116
rect 11950 27966 11996 28012
rect 11950 27862 11996 27908
rect 11950 27758 11996 27804
rect 12174 28594 12220 28640
rect 12174 28489 12220 28535
rect 12174 28384 12220 28430
rect 12174 28279 12220 28325
rect 12174 28174 12220 28220
rect 12174 28070 12220 28116
rect 12174 27966 12220 28012
rect 12174 27862 12220 27908
rect 12174 27758 12220 27804
rect 12398 28594 12444 28640
rect 12398 28489 12444 28535
rect 12398 28384 12444 28430
rect 12398 28279 12444 28325
rect 12398 28174 12444 28220
rect 12398 28070 12444 28116
rect 12398 27966 12444 28012
rect 12398 27862 12444 27908
rect 12398 27758 12444 27804
rect 12622 28594 12668 28640
rect 12622 28489 12668 28535
rect 12622 28384 12668 28430
rect 12622 28279 12668 28325
rect 12622 28174 12668 28220
rect 12622 28070 12668 28116
rect 23797 28144 23843 28190
rect 12622 27966 12668 28012
rect 12622 27862 12668 27908
rect 13312 27834 13358 28082
rect 13536 27834 13582 28082
rect 13760 27834 13806 28082
rect 16704 28030 16750 28076
rect 12622 27758 12668 27804
rect 14906 27950 14952 27996
rect 14906 27830 14952 27876
rect 15130 27950 15176 27996
rect 15130 27830 15176 27876
rect 16704 27925 16750 27971
rect 16704 27820 16750 27866
rect 6091 26379 6137 26731
rect 6091 26276 6137 26322
rect 6091 26173 6137 26219
rect 6091 26070 6137 26116
rect 6091 25967 6137 26013
rect 6091 25864 6137 25910
rect 6091 25761 6137 25807
rect 6091 25658 6137 25704
rect 6091 25555 6137 25601
rect 6091 25452 6137 25498
rect 6091 25349 6137 25395
rect 6315 26379 6361 26731
rect 6315 26276 6361 26322
rect 6315 26173 6361 26219
rect 6315 26070 6361 26116
rect 6315 25967 6361 26013
rect 6315 25864 6361 25910
rect 6315 25761 6361 25807
rect 6315 25658 6361 25704
rect 6315 25555 6361 25601
rect 6315 25452 6361 25498
rect 6605 26400 6651 26446
rect 6605 26292 6651 26338
rect 6605 26184 6651 26230
rect 6605 26076 6651 26122
rect 6605 25968 6651 26014
rect 6605 25860 6651 25906
rect 6605 25752 6651 25798
rect 6605 25644 6651 25690
rect 6605 25536 6651 25582
rect 6605 25428 6651 25474
rect 6829 26400 6875 26446
rect 6829 26292 6875 26338
rect 6829 26184 6875 26230
rect 6829 26076 6875 26122
rect 6829 25968 6875 26014
rect 6829 25860 6875 25906
rect 6829 25752 6875 25798
rect 6829 25644 6875 25690
rect 6829 25536 6875 25582
rect 6829 25428 6875 25474
rect 7782 26379 7828 26731
rect 7782 26276 7828 26322
rect 7782 26173 7828 26219
rect 7782 26070 7828 26116
rect 7782 25967 7828 26013
rect 7782 25864 7828 25910
rect 7782 25761 7828 25807
rect 7782 25658 7828 25704
rect 7782 25555 7828 25601
rect 7782 25452 7828 25498
rect 6315 25349 6361 25395
rect 7782 25349 7828 25395
rect 8006 26379 8052 26731
rect 8006 26276 8052 26322
rect 8006 26173 8052 26219
rect 8006 26070 8052 26116
rect 8006 25967 8052 26013
rect 8006 25864 8052 25910
rect 8006 25761 8052 25807
rect 8006 25658 8052 25704
rect 8006 25555 8052 25601
rect 8006 25452 8052 25498
rect 8296 26400 8342 26446
rect 8296 26292 8342 26338
rect 8296 26184 8342 26230
rect 8296 26076 8342 26122
rect 8296 25968 8342 26014
rect 8296 25860 8342 25906
rect 8296 25752 8342 25798
rect 8296 25644 8342 25690
rect 8296 25536 8342 25582
rect 8296 25428 8342 25474
rect 8520 26400 8566 26446
rect 8520 26292 8566 26338
rect 8520 26184 8566 26230
rect 8520 26076 8566 26122
rect 8520 25968 8566 26014
rect 8520 25860 8566 25906
rect 8520 25752 8566 25798
rect 8520 25644 8566 25690
rect 8520 25536 8566 25582
rect 8520 25428 8566 25474
rect 8006 25349 8052 25395
rect 16704 27715 16750 27761
rect 16704 27610 16750 27656
rect 16704 27506 16750 27552
rect 16704 27402 16750 27448
rect 16704 27298 16750 27344
rect 16704 27194 16750 27240
rect 16928 28030 16974 28076
rect 16928 27925 16974 27971
rect 16928 27820 16974 27866
rect 16928 27715 16974 27761
rect 16928 27610 16974 27656
rect 16928 27506 16974 27552
rect 16928 27402 16974 27448
rect 16928 27298 16974 27344
rect 16928 27194 16974 27240
rect 17152 28030 17198 28076
rect 17152 27925 17198 27971
rect 17152 27820 17198 27866
rect 17152 27715 17198 27761
rect 17152 27610 17198 27656
rect 17152 27506 17198 27552
rect 17152 27402 17198 27448
rect 17152 27298 17198 27344
rect 17152 27194 17198 27240
rect 17376 28030 17422 28076
rect 17376 27925 17422 27971
rect 17376 27820 17422 27866
rect 17376 27715 17422 27761
rect 17376 27610 17422 27656
rect 17376 27506 17422 27552
rect 17376 27402 17422 27448
rect 17376 27298 17422 27344
rect 17376 27194 17422 27240
rect 17600 28030 17646 28076
rect 17600 27925 17646 27971
rect 17600 27820 17646 27866
rect 17600 27715 17646 27761
rect 17600 27610 17646 27656
rect 17600 27506 17646 27552
rect 17600 27402 17646 27448
rect 17600 27298 17646 27344
rect 17600 27194 17646 27240
rect 17824 28030 17870 28076
rect 17824 27925 17870 27971
rect 17824 27820 17870 27866
rect 17824 27715 17870 27761
rect 17824 27610 17870 27656
rect 17824 27506 17870 27552
rect 17824 27402 17870 27448
rect 17824 27298 17870 27344
rect 17824 27194 17870 27240
rect 18048 28030 18094 28076
rect 18048 27925 18094 27971
rect 18048 27820 18094 27866
rect 18048 27715 18094 27761
rect 18048 27610 18094 27656
rect 18048 27506 18094 27552
rect 18048 27402 18094 27448
rect 18048 27298 18094 27344
rect 18048 27194 18094 27240
rect 18338 28030 18384 28076
rect 18338 27925 18384 27971
rect 18338 27820 18384 27866
rect 18338 27715 18384 27761
rect 18338 27610 18384 27656
rect 18338 27506 18384 27552
rect 18338 27402 18384 27448
rect 18338 27298 18384 27344
rect 18338 27194 18384 27240
rect 18562 28030 18608 28076
rect 18562 27925 18608 27971
rect 18562 27820 18608 27866
rect 18562 27715 18608 27761
rect 18562 27610 18608 27656
rect 18562 27506 18608 27552
rect 18562 27402 18608 27448
rect 18562 27298 18608 27344
rect 18562 27194 18608 27240
rect 18786 28030 18832 28076
rect 18786 27925 18832 27971
rect 18786 27820 18832 27866
rect 18786 27715 18832 27761
rect 18786 27610 18832 27656
rect 18786 27506 18832 27552
rect 18786 27402 18832 27448
rect 18786 27298 18832 27344
rect 18786 27194 18832 27240
rect 19010 28030 19056 28076
rect 19010 27925 19056 27971
rect 19010 27820 19056 27866
rect 19010 27715 19056 27761
rect 19010 27610 19056 27656
rect 19010 27506 19056 27552
rect 19010 27402 19056 27448
rect 19010 27298 19056 27344
rect 19010 27194 19056 27240
rect 19234 28030 19280 28076
rect 19234 27925 19280 27971
rect 19234 27820 19280 27866
rect 19234 27715 19280 27761
rect 19234 27610 19280 27656
rect 19234 27506 19280 27552
rect 19234 27402 19280 27448
rect 19234 27298 19280 27344
rect 19234 27194 19280 27240
rect 19458 28030 19504 28076
rect 19458 27925 19504 27971
rect 19458 27820 19504 27866
rect 19458 27715 19504 27761
rect 19458 27610 19504 27656
rect 19458 27506 19504 27552
rect 19458 27402 19504 27448
rect 19458 27298 19504 27344
rect 19458 27194 19504 27240
rect 19682 28030 19728 28076
rect 19682 27925 19728 27971
rect 19682 27820 19728 27866
rect 19682 27715 19728 27761
rect 19682 27610 19728 27656
rect 19682 27506 19728 27552
rect 19682 27402 19728 27448
rect 19682 27298 19728 27344
rect 19682 27194 19728 27240
rect 19971 28030 20017 28076
rect 19971 27925 20017 27971
rect 19971 27820 20017 27866
rect 19971 27715 20017 27761
rect 19971 27610 20017 27656
rect 19971 27506 20017 27552
rect 19971 27402 20017 27448
rect 19971 27298 20017 27344
rect 19971 27194 20017 27240
rect 20195 28030 20241 28076
rect 20195 27925 20241 27971
rect 20195 27820 20241 27866
rect 20195 27715 20241 27761
rect 20195 27610 20241 27656
rect 20195 27506 20241 27552
rect 20195 27402 20241 27448
rect 20195 27298 20241 27344
rect 20195 27194 20241 27240
rect 20419 28030 20465 28076
rect 20419 27925 20465 27971
rect 20419 27820 20465 27866
rect 20419 27715 20465 27761
rect 20419 27610 20465 27656
rect 20419 27506 20465 27552
rect 20419 27402 20465 27448
rect 20419 27298 20465 27344
rect 20419 27194 20465 27240
rect 20643 28030 20689 28076
rect 20643 27925 20689 27971
rect 20643 27820 20689 27866
rect 20643 27715 20689 27761
rect 20643 27610 20689 27656
rect 20643 27506 20689 27552
rect 20643 27402 20689 27448
rect 20643 27298 20689 27344
rect 20643 27194 20689 27240
rect 20867 28030 20913 28076
rect 20867 27925 20913 27971
rect 20867 27820 20913 27866
rect 20867 27715 20913 27761
rect 20867 27610 20913 27656
rect 20867 27506 20913 27552
rect 20867 27402 20913 27448
rect 20867 27298 20913 27344
rect 20867 27194 20913 27240
rect 21091 28030 21137 28076
rect 21091 27925 21137 27971
rect 21091 27820 21137 27866
rect 21091 27715 21137 27761
rect 21091 27610 21137 27656
rect 21091 27506 21137 27552
rect 21091 27402 21137 27448
rect 21091 27298 21137 27344
rect 21091 27194 21137 27240
rect 21315 28030 21361 28076
rect 21315 27925 21361 27971
rect 21315 27820 21361 27866
rect 21315 27715 21361 27761
rect 21315 27610 21361 27656
rect 21315 27506 21361 27552
rect 21315 27402 21361 27448
rect 21315 27298 21361 27344
rect 21315 27194 21361 27240
rect 21605 28030 21651 28076
rect 21605 27925 21651 27971
rect 21605 27820 21651 27866
rect 21605 27715 21651 27761
rect 21605 27610 21651 27656
rect 21605 27506 21651 27552
rect 21605 27402 21651 27448
rect 21605 27298 21651 27344
rect 21605 27194 21651 27240
rect 21829 28030 21875 28076
rect 21829 27925 21875 27971
rect 21829 27820 21875 27866
rect 21829 27715 21875 27761
rect 21829 27610 21875 27656
rect 21829 27506 21875 27552
rect 21829 27402 21875 27448
rect 21829 27298 21875 27344
rect 21829 27194 21875 27240
rect 22053 28030 22099 28076
rect 22053 27925 22099 27971
rect 22053 27820 22099 27866
rect 22053 27715 22099 27761
rect 22053 27610 22099 27656
rect 22053 27506 22099 27552
rect 22053 27402 22099 27448
rect 22053 27298 22099 27344
rect 22053 27194 22099 27240
rect 22277 28030 22323 28076
rect 22277 27925 22323 27971
rect 22277 27820 22323 27866
rect 22277 27715 22323 27761
rect 22277 27610 22323 27656
rect 22277 27506 22323 27552
rect 22277 27402 22323 27448
rect 22277 27298 22323 27344
rect 22277 27194 22323 27240
rect 22501 28030 22547 28076
rect 22501 27925 22547 27971
rect 22501 27820 22547 27866
rect 22501 27715 22547 27761
rect 22501 27610 22547 27656
rect 22501 27506 22547 27552
rect 22501 27402 22547 27448
rect 22501 27298 22547 27344
rect 22501 27194 22547 27240
rect 22725 28030 22771 28076
rect 22725 27925 22771 27971
rect 22725 27820 22771 27866
rect 22725 27715 22771 27761
rect 22725 27610 22771 27656
rect 22725 27506 22771 27552
rect 22725 27402 22771 27448
rect 22725 27298 22771 27344
rect 22725 27194 22771 27240
rect 22949 28030 22995 28076
rect 22949 27925 22995 27971
rect 22949 27820 22995 27866
rect 23797 28041 23843 28087
rect 23797 27938 23843 27984
rect 23797 27834 23843 27880
rect 24021 28144 24067 28190
rect 24021 28041 24067 28087
rect 24021 27938 24067 27984
rect 24021 27834 24067 27880
rect 24245 28144 24291 28190
rect 24245 28041 24291 28087
rect 24245 27938 24291 27984
rect 24245 27834 24291 27880
rect 22949 27715 22995 27761
rect 22949 27610 22995 27656
rect 22949 27506 22995 27552
rect 25392 27830 25438 28076
rect 25616 27830 25662 28076
rect 22949 27402 22995 27448
rect 22949 27298 22995 27344
rect 22949 27194 22995 27240
rect 13470 26379 13516 26731
rect 13470 26276 13516 26322
rect 13470 26173 13516 26219
rect 13470 26070 13516 26116
rect 13470 25967 13516 26013
rect 13470 25864 13516 25910
rect 13470 25761 13516 25807
rect 13470 25658 13516 25704
rect 13470 25555 13516 25601
rect 13470 25452 13516 25498
rect 13470 25349 13516 25395
rect 13694 26379 13740 26731
rect 13694 26276 13740 26322
rect 13694 26173 13740 26219
rect 13694 26070 13740 26116
rect 13694 25967 13740 26013
rect 13694 25864 13740 25910
rect 13694 25761 13740 25807
rect 13694 25658 13740 25704
rect 13694 25555 13740 25601
rect 13694 25452 13740 25498
rect 13984 26400 14030 26446
rect 13984 26292 14030 26338
rect 13984 26184 14030 26230
rect 13984 26076 14030 26122
rect 13984 25968 14030 26014
rect 13984 25860 14030 25906
rect 13984 25752 14030 25798
rect 13984 25644 14030 25690
rect 13984 25536 14030 25582
rect 13984 25428 14030 25474
rect 14208 26400 14254 26446
rect 14208 26292 14254 26338
rect 14208 26184 14254 26230
rect 14208 26076 14254 26122
rect 14208 25968 14254 26014
rect 14208 25860 14254 25906
rect 14208 25752 14254 25798
rect 14208 25644 14254 25690
rect 14208 25536 14254 25582
rect 14208 25428 14254 25474
rect 15161 26379 15207 26731
rect 15161 26276 15207 26322
rect 15161 26173 15207 26219
rect 15161 26070 15207 26116
rect 15161 25967 15207 26013
rect 15161 25864 15207 25910
rect 15161 25761 15207 25807
rect 15161 25658 15207 25704
rect 15161 25555 15207 25601
rect 15161 25452 15207 25498
rect 13694 25349 13740 25395
rect 15161 25349 15207 25395
rect 15385 26379 15431 26731
rect 15385 26276 15431 26322
rect 15385 26173 15431 26219
rect 15385 26070 15431 26116
rect 15385 25967 15431 26013
rect 15385 25864 15431 25910
rect 15385 25761 15431 25807
rect 15385 25658 15431 25704
rect 15385 25555 15431 25601
rect 15385 25452 15431 25498
rect 15675 26400 15721 26446
rect 15675 26292 15721 26338
rect 15675 26184 15721 26230
rect 15675 26076 15721 26122
rect 15675 25968 15721 26014
rect 15675 25860 15721 25906
rect 15675 25752 15721 25798
rect 15675 25644 15721 25690
rect 15675 25536 15721 25582
rect 15675 25428 15721 25474
rect 15899 26400 15945 26446
rect 15899 26292 15945 26338
rect 15899 26184 15945 26230
rect 15899 26076 15945 26122
rect 15899 25968 15945 26014
rect 15899 25860 15945 25906
rect 15899 25752 15945 25798
rect 15899 25644 15945 25690
rect 15899 25536 15945 25582
rect 15899 25428 15945 25474
rect 15385 25349 15431 25395
rect 23956 26684 24002 26730
rect 23956 26581 24002 26627
rect 23956 26478 24002 26524
rect 23956 26375 24002 26421
rect 23956 26272 24002 26318
rect 23956 26168 24002 26214
rect 23956 26064 24002 26110
rect 23956 25960 24002 26006
rect 23956 25856 24002 25902
rect 23956 25752 24002 25798
rect 23956 25648 24002 25694
rect 23956 25544 24002 25590
rect 23956 25440 24002 25486
rect 24180 26684 24226 26730
rect 24180 26581 24226 26627
rect 24180 26478 24226 26524
rect 24180 26375 24226 26421
rect 24180 26272 24226 26318
rect 24180 26168 24226 26214
rect 24180 26064 24226 26110
rect 24180 25960 24226 26006
rect 24180 25856 24226 25902
rect 24180 25752 24226 25798
rect 24180 25648 24226 25694
rect 24180 25544 24226 25590
rect 24180 25440 24226 25486
rect 24470 26684 24516 26730
rect 24470 26581 24516 26627
rect 24470 26478 24516 26524
rect 24470 26375 24516 26421
rect 24470 26272 24516 26318
rect 24470 26168 24516 26214
rect 24470 26064 24516 26110
rect 24470 25960 24516 26006
rect 24470 25856 24516 25902
rect 24470 25752 24516 25798
rect 24470 25648 24516 25694
rect 24470 25544 24516 25590
rect 24470 25440 24516 25486
rect 24694 26684 24740 26730
rect 24694 26581 24740 26627
rect 24694 26478 24740 26524
rect 24694 26375 24740 26421
rect 24694 26272 24740 26318
rect 24694 26168 24740 26214
rect 24694 26064 24740 26110
rect 24694 25960 24740 26006
rect 24694 25856 24740 25902
rect 24694 25752 24740 25798
rect 24694 25648 24740 25694
rect 24694 25544 24740 25590
rect 25646 26684 25692 26730
rect 25646 26581 25692 26627
rect 25646 26478 25692 26524
rect 25646 26375 25692 26421
rect 25646 26272 25692 26318
rect 25646 26168 25692 26214
rect 25646 26064 25692 26110
rect 25646 25960 25692 26006
rect 25646 25856 25692 25902
rect 25646 25752 25692 25798
rect 25646 25648 25692 25694
rect 24694 25440 24740 25486
rect 25646 25544 25692 25590
rect 25646 25440 25692 25486
rect 25870 26684 25916 26730
rect 25870 26581 25916 26627
rect 25870 26478 25916 26524
rect 25870 26375 25916 26421
rect 25870 26272 25916 26318
rect 25870 26168 25916 26214
rect 25870 26064 25916 26110
rect 25870 25960 25916 26006
rect 25870 25856 25916 25902
rect 25870 25752 25916 25798
rect 25870 25648 25916 25694
rect 25870 25544 25916 25590
rect 25870 25440 25916 25486
rect 26160 26684 26206 26730
rect 26160 26581 26206 26627
rect 26160 26478 26206 26524
rect 26160 26375 26206 26421
rect 26160 26272 26206 26318
rect 26160 26168 26206 26214
rect 26160 26064 26206 26110
rect 26160 25960 26206 26006
rect 26160 25856 26206 25902
rect 26160 25752 26206 25798
rect 26160 25648 26206 25694
rect 26160 25544 26206 25590
rect 26160 25440 26206 25486
rect 26384 26684 26430 26730
rect 26384 26581 26430 26627
rect 26384 26478 26430 26524
rect 26384 26375 26430 26421
rect 26384 26272 26430 26318
rect 26384 26168 26430 26214
rect 26384 26064 26430 26110
rect 26384 25960 26430 26006
rect 26384 25856 26430 25902
rect 26384 25752 26430 25798
rect 26384 25648 26430 25694
rect 26384 25544 26430 25590
rect 27337 26684 27383 26730
rect 27337 26581 27383 26627
rect 27337 26478 27383 26524
rect 27337 26375 27383 26421
rect 27337 26272 27383 26318
rect 27337 26168 27383 26214
rect 27337 26064 27383 26110
rect 27337 25960 27383 26006
rect 27337 25856 27383 25902
rect 27337 25752 27383 25798
rect 27337 25648 27383 25694
rect 26384 25440 26430 25486
rect 27337 25544 27383 25590
rect 27337 25440 27383 25486
rect 27561 26684 27607 26730
rect 27561 26581 27607 26627
rect 27561 26478 27607 26524
rect 27561 26375 27607 26421
rect 27561 26272 27607 26318
rect 27561 26168 27607 26214
rect 27561 26064 27607 26110
rect 27561 25960 27607 26006
rect 27561 25856 27607 25902
rect 27561 25752 27607 25798
rect 27561 25648 27607 25694
rect 27561 25544 27607 25590
rect 27561 25440 27607 25486
rect 27851 26684 27897 26730
rect 27851 26581 27897 26627
rect 27851 26478 27897 26524
rect 27851 26375 27897 26421
rect 27851 26272 27897 26318
rect 27851 26168 27897 26214
rect 27851 26064 27897 26110
rect 27851 25960 27897 26006
rect 27851 25856 27897 25902
rect 27851 25752 27897 25798
rect 27851 25648 27897 25694
rect 27851 25544 27897 25590
rect 27851 25440 27897 25486
rect 28075 26684 28121 26730
rect 28075 26581 28121 26627
rect 28075 26478 28121 26524
rect 28075 26375 28121 26421
rect 28075 26272 28121 26318
rect 28075 26168 28121 26214
rect 28075 26064 28121 26110
rect 28075 25960 28121 26006
rect 28075 25856 28121 25902
rect 28075 25752 28121 25798
rect 28075 25648 28121 25694
rect 28075 25544 28121 25590
rect 28075 25440 28121 25486
rect 1817 20460 1863 20506
rect 1817 20292 1863 20338
rect 1817 20125 1863 20171
rect 1817 19957 1863 20003
rect 1817 19789 1863 19835
rect 1817 19621 1863 19667
rect 1817 19453 1863 19499
rect 1817 19286 1863 19332
rect 1817 19118 1863 19164
rect 1817 18950 1863 18996
rect 1817 18782 1863 18828
rect 1817 18612 1863 18658
rect 1817 18442 1863 18488
rect 1817 18272 1863 18318
rect 2266 20460 2312 20506
rect 2266 20292 2312 20338
rect 2266 20125 2312 20171
rect 2266 19957 2312 20003
rect 2266 19789 2312 19835
rect 2266 19621 2312 19667
rect 2266 19453 2312 19499
rect 2266 19286 2312 19332
rect 2266 19118 2312 19164
rect 2266 18950 2312 18996
rect 2266 18782 2312 18828
rect 2266 18612 2312 18658
rect 2266 18442 2312 18488
rect 2266 18272 2312 18318
rect 2844 20460 2890 20506
rect 2844 20292 2890 20338
rect 2844 20125 2890 20171
rect 2844 19957 2890 20003
rect 2844 19789 2890 19835
rect 2844 19621 2890 19667
rect 2844 19453 2890 19499
rect 2844 19286 2890 19332
rect 2844 19118 2890 19164
rect 2844 18950 2890 18996
rect 2844 18782 2890 18828
rect 2844 18612 2890 18658
rect 2844 18442 2890 18488
rect 2844 18272 2890 18318
rect 3293 20460 3339 20506
rect 3293 20292 3339 20338
rect 3293 20125 3339 20171
rect 3293 19957 3339 20003
rect 3293 19789 3339 19835
rect 3293 19621 3339 19667
rect 3293 19453 3339 19499
rect 3293 19286 3339 19332
rect 3293 19118 3339 19164
rect 3293 18950 3339 18996
rect 3293 18782 3339 18828
rect 3293 18612 3339 18658
rect 3293 18442 3339 18488
rect 3293 18272 3339 18318
rect 3609 20460 3655 20506
rect 3609 20292 3655 20338
rect 3609 20125 3655 20171
rect 3609 19957 3655 20003
rect 3609 19789 3655 19835
rect 3609 19621 3655 19667
rect 3609 19453 3655 19499
rect 3609 19286 3655 19332
rect 3609 19118 3655 19164
rect 3609 18950 3655 18996
rect 3609 18782 3655 18828
rect 3609 18612 3655 18658
rect 3609 18442 3655 18488
rect 3609 18272 3655 18318
rect 4058 20460 4104 20506
rect 4058 20292 4104 20338
rect 4058 20125 4104 20171
rect 4058 19957 4104 20003
rect 4058 19789 4104 19835
rect 4058 19621 4104 19667
rect 4058 19453 4104 19499
rect 4058 19286 4104 19332
rect 4058 19118 4104 19164
rect 4058 18950 4104 18996
rect 4058 18782 4104 18828
rect 4058 18612 4104 18658
rect 4058 18442 4104 18488
rect 4058 18272 4104 18318
rect 4636 20460 4682 20506
rect 4636 20292 4682 20338
rect 4636 20125 4682 20171
rect 4636 19957 4682 20003
rect 4636 19789 4682 19835
rect 4636 19621 4682 19667
rect 4636 19453 4682 19499
rect 4636 19286 4682 19332
rect 4636 19118 4682 19164
rect 4636 18950 4682 18996
rect 4636 18782 4682 18828
rect 4636 18612 4682 18658
rect 4636 18442 4682 18488
rect 4636 18272 4682 18318
rect 5085 20460 5131 20506
rect 5085 20292 5131 20338
rect 5085 20125 5131 20171
rect 5085 19957 5131 20003
rect 5085 19789 5131 19835
rect 5085 19621 5131 19667
rect 5085 19453 5131 19499
rect 5085 19286 5131 19332
rect 5085 19118 5131 19164
rect 5085 18950 5131 18996
rect 5085 18782 5131 18828
rect 5085 18612 5131 18658
rect 5085 18442 5131 18488
rect 5085 18272 5131 18318
rect 9196 20460 9242 20506
rect 9196 20292 9242 20338
rect 9196 20125 9242 20171
rect 9196 19957 9242 20003
rect 9196 19789 9242 19835
rect 9196 19621 9242 19667
rect 9196 19453 9242 19499
rect 9196 19286 9242 19332
rect 9196 19118 9242 19164
rect 9196 18950 9242 18996
rect 9196 18782 9242 18828
rect 9196 18612 9242 18658
rect 9196 18442 9242 18488
rect 9196 18272 9242 18318
rect 9645 20460 9691 20506
rect 9645 20292 9691 20338
rect 9645 20125 9691 20171
rect 9645 19957 9691 20003
rect 9645 19789 9691 19835
rect 9645 19621 9691 19667
rect 9645 19453 9691 19499
rect 9645 19286 9691 19332
rect 9645 19118 9691 19164
rect 9645 18950 9691 18996
rect 9645 18782 9691 18828
rect 9645 18612 9691 18658
rect 9645 18442 9691 18488
rect 9645 18272 9691 18318
rect 10223 20460 10269 20506
rect 10223 20292 10269 20338
rect 10223 20125 10269 20171
rect 10223 19957 10269 20003
rect 10223 19789 10269 19835
rect 10223 19621 10269 19667
rect 10223 19453 10269 19499
rect 10223 19286 10269 19332
rect 10223 19118 10269 19164
rect 10223 18950 10269 18996
rect 10223 18782 10269 18828
rect 10223 18612 10269 18658
rect 10223 18442 10269 18488
rect 10223 18272 10269 18318
rect 10672 20460 10718 20506
rect 10672 20292 10718 20338
rect 10672 20125 10718 20171
rect 10672 19957 10718 20003
rect 10672 19789 10718 19835
rect 10672 19621 10718 19667
rect 10672 19453 10718 19499
rect 10672 19286 10718 19332
rect 10672 19118 10718 19164
rect 10672 18950 10718 18996
rect 10672 18782 10718 18828
rect 10672 18612 10718 18658
rect 10672 18442 10718 18488
rect 10672 18272 10718 18318
rect 10988 20460 11034 20506
rect 10988 20292 11034 20338
rect 10988 20125 11034 20171
rect 10988 19957 11034 20003
rect 10988 19789 11034 19835
rect 10988 19621 11034 19667
rect 10988 19453 11034 19499
rect 10988 19286 11034 19332
rect 10988 19118 11034 19164
rect 10988 18950 11034 18996
rect 10988 18782 11034 18828
rect 10988 18612 11034 18658
rect 10988 18442 11034 18488
rect 10988 18272 11034 18318
rect 11437 20460 11483 20506
rect 11437 20292 11483 20338
rect 11437 20125 11483 20171
rect 11437 19957 11483 20003
rect 11437 19789 11483 19835
rect 11437 19621 11483 19667
rect 11437 19453 11483 19499
rect 11437 19286 11483 19332
rect 11437 19118 11483 19164
rect 11437 18950 11483 18996
rect 11437 18782 11483 18828
rect 11437 18612 11483 18658
rect 11437 18442 11483 18488
rect 11437 18272 11483 18318
rect 12015 20460 12061 20506
rect 12015 20292 12061 20338
rect 12015 20125 12061 20171
rect 12015 19957 12061 20003
rect 12015 19789 12061 19835
rect 12015 19621 12061 19667
rect 12015 19453 12061 19499
rect 12015 19286 12061 19332
rect 12015 19118 12061 19164
rect 12015 18950 12061 18996
rect 12015 18782 12061 18828
rect 12015 18612 12061 18658
rect 12015 18442 12061 18488
rect 12015 18272 12061 18318
rect 12464 20460 12510 20506
rect 12464 20292 12510 20338
rect 12464 20125 12510 20171
rect 12464 19957 12510 20003
rect 12464 19789 12510 19835
rect 12464 19621 12510 19667
rect 12464 19453 12510 19499
rect 12464 19286 12510 19332
rect 12464 19118 12510 19164
rect 12464 18950 12510 18996
rect 12464 18782 12510 18828
rect 12464 18612 12510 18658
rect 12464 18442 12510 18488
rect 12464 18272 12510 18318
rect 16704 20446 16750 20492
rect 16704 20279 16750 20325
rect 16704 20111 16750 20157
rect 16704 19943 16750 19989
rect 16704 19775 16750 19821
rect 16704 19608 16750 19654
rect 16704 19440 16750 19486
rect 16704 19272 16750 19318
rect 16704 19104 16750 19150
rect 16704 18936 16750 18982
rect 16704 18769 16750 18815
rect 16704 18599 16750 18645
rect 16704 18429 16750 18475
rect 16704 18259 16750 18305
rect 16704 18089 16750 18135
rect 17376 20446 17422 20492
rect 17376 20279 17422 20325
rect 17376 20111 17422 20157
rect 17376 19943 17422 19989
rect 17376 19775 17422 19821
rect 17376 19608 17422 19654
rect 17376 19440 17422 19486
rect 17376 19272 17422 19318
rect 17376 19104 17422 19150
rect 17376 18936 17422 18982
rect 17376 18769 17422 18815
rect 17376 18599 17422 18645
rect 17376 18429 17422 18475
rect 17376 18259 17422 18305
rect 17376 18089 17422 18135
rect 18048 20446 18094 20492
rect 18048 20279 18094 20325
rect 18048 20111 18094 20157
rect 18048 19943 18094 19989
rect 18048 19775 18094 19821
rect 18048 19608 18094 19654
rect 18048 19440 18094 19486
rect 18048 19272 18094 19318
rect 18048 19104 18094 19150
rect 18048 18936 18094 18982
rect 18048 18769 18094 18815
rect 18048 18599 18094 18645
rect 18048 18429 18094 18475
rect 18048 18259 18094 18305
rect 18048 18089 18094 18135
rect 18338 20446 18384 20492
rect 18338 20279 18384 20325
rect 18338 20111 18384 20157
rect 18338 19943 18384 19989
rect 18338 19775 18384 19821
rect 18338 19608 18384 19654
rect 18338 19440 18384 19486
rect 18338 19272 18384 19318
rect 18338 19104 18384 19150
rect 18338 18936 18384 18982
rect 18338 18769 18384 18815
rect 18338 18599 18384 18645
rect 18338 18429 18384 18475
rect 18338 18259 18384 18305
rect 18338 18089 18384 18135
rect 19010 20446 19056 20492
rect 19010 20279 19056 20325
rect 19010 20111 19056 20157
rect 19010 19943 19056 19989
rect 19010 19775 19056 19821
rect 19010 19608 19056 19654
rect 19010 19440 19056 19486
rect 19010 19272 19056 19318
rect 19010 19104 19056 19150
rect 19010 18936 19056 18982
rect 19010 18769 19056 18815
rect 19010 18599 19056 18645
rect 19010 18429 19056 18475
rect 19010 18259 19056 18305
rect 19010 18089 19056 18135
rect 19682 20446 19728 20492
rect 19682 20279 19728 20325
rect 19682 20111 19728 20157
rect 19682 19943 19728 19989
rect 19682 19775 19728 19821
rect 19682 19608 19728 19654
rect 19682 19440 19728 19486
rect 19682 19272 19728 19318
rect 19682 19104 19728 19150
rect 19682 18936 19728 18982
rect 19682 18769 19728 18815
rect 19682 18599 19728 18645
rect 19682 18429 19728 18475
rect 19682 18259 19728 18305
rect 19682 18089 19728 18135
rect 19971 20446 20017 20492
rect 19971 20279 20017 20325
rect 19971 20111 20017 20157
rect 19971 19943 20017 19989
rect 19971 19775 20017 19821
rect 19971 19608 20017 19654
rect 19971 19440 20017 19486
rect 19971 19272 20017 19318
rect 19971 19104 20017 19150
rect 19971 18936 20017 18982
rect 19971 18769 20017 18815
rect 19971 18599 20017 18645
rect 19971 18429 20017 18475
rect 19971 18259 20017 18305
rect 19971 18089 20017 18135
rect 20643 20446 20689 20492
rect 20643 20279 20689 20325
rect 20643 20111 20689 20157
rect 20643 19943 20689 19989
rect 20643 19775 20689 19821
rect 20643 19608 20689 19654
rect 20643 19440 20689 19486
rect 20643 19272 20689 19318
rect 20643 19104 20689 19150
rect 20643 18936 20689 18982
rect 20643 18769 20689 18815
rect 20643 18599 20689 18645
rect 20643 18429 20689 18475
rect 20643 18259 20689 18305
rect 20643 18089 20689 18135
rect 21315 20446 21361 20492
rect 21315 20279 21361 20325
rect 21315 20111 21361 20157
rect 21315 19943 21361 19989
rect 21315 19775 21361 19821
rect 21315 19608 21361 19654
rect 21315 19440 21361 19486
rect 21315 19272 21361 19318
rect 21315 19104 21361 19150
rect 21315 18936 21361 18982
rect 21315 18769 21361 18815
rect 21315 18599 21361 18645
rect 21315 18429 21361 18475
rect 21315 18259 21361 18305
rect 21315 18089 21361 18135
rect 21605 20446 21651 20492
rect 21605 20279 21651 20325
rect 21605 20111 21651 20157
rect 21605 19943 21651 19989
rect 21605 19775 21651 19821
rect 21605 19608 21651 19654
rect 21605 19440 21651 19486
rect 21605 19272 21651 19318
rect 21605 19104 21651 19150
rect 21605 18936 21651 18982
rect 21605 18769 21651 18815
rect 21605 18599 21651 18645
rect 21605 18429 21651 18475
rect 21605 18259 21651 18305
rect 21605 18089 21651 18135
rect 22277 20446 22323 20492
rect 22277 20279 22323 20325
rect 22277 20111 22323 20157
rect 22277 19943 22323 19989
rect 22277 19775 22323 19821
rect 22277 19608 22323 19654
rect 22277 19440 22323 19486
rect 22277 19272 22323 19318
rect 22277 19104 22323 19150
rect 22277 18936 22323 18982
rect 22277 18769 22323 18815
rect 22277 18599 22323 18645
rect 22277 18429 22323 18475
rect 22277 18259 22323 18305
rect 22277 18089 22323 18135
rect 22949 20446 22995 20492
rect 22949 20279 22995 20325
rect 22949 20111 22995 20157
rect 22949 19943 22995 19989
rect 22949 19775 22995 19821
rect 22949 19608 22995 19654
rect 22949 19440 22995 19486
rect 22949 19272 22995 19318
rect 22949 19104 22995 19150
rect 22949 18936 22995 18982
rect 22949 18769 22995 18815
rect 22949 18599 22995 18645
rect 22949 18429 22995 18475
rect 22949 18259 22995 18305
rect 22949 18089 22995 18135
rect 1995 10997 2041 11757
rect 1995 10894 2041 10940
rect 1995 10791 2041 10837
rect 1995 10688 2041 10734
rect 1995 10585 2041 10631
rect 1995 10482 2041 10528
rect 1995 10379 2041 10425
rect 1995 10276 2041 10322
rect 1995 10173 2041 10219
rect 1995 10070 2041 10116
rect 1995 9967 2041 10013
rect 2219 10997 2265 11757
rect 2219 10894 2265 10940
rect 2219 10791 2265 10837
rect 2219 10688 2265 10734
rect 2219 10585 2265 10631
rect 2219 10482 2265 10528
rect 2219 10379 2265 10425
rect 2219 10276 2265 10322
rect 2219 10173 2265 10219
rect 2219 10070 2265 10116
rect 2219 9967 2265 10013
rect 2443 10997 2489 11757
rect 2443 10894 2489 10940
rect 2443 10791 2489 10837
rect 2443 10688 2489 10734
rect 2443 10585 2489 10631
rect 2443 10482 2489 10528
rect 2443 10379 2489 10425
rect 2443 10276 2489 10322
rect 2443 10173 2489 10219
rect 2443 10070 2489 10116
rect 2443 9967 2489 10013
rect 2667 10997 2713 11757
rect 2667 10894 2713 10940
rect 2667 10791 2713 10837
rect 2667 10688 2713 10734
rect 2667 10585 2713 10631
rect 2667 10482 2713 10528
rect 2667 10379 2713 10425
rect 2667 10276 2713 10322
rect 2667 10173 2713 10219
rect 2667 10070 2713 10116
rect 2667 9967 2713 10013
rect 2891 10997 2937 11757
rect 2891 10894 2937 10940
rect 2891 10791 2937 10837
rect 2891 10688 2937 10734
rect 2891 10585 2937 10631
rect 2891 10482 2937 10528
rect 2891 10379 2937 10425
rect 2891 10276 2937 10322
rect 2891 10173 2937 10219
rect 2891 10070 2937 10116
rect 2891 9967 2937 10013
rect 3115 10997 3161 11757
rect 3115 10894 3161 10940
rect 3115 10791 3161 10837
rect 3115 10688 3161 10734
rect 3115 10585 3161 10631
rect 3115 10482 3161 10528
rect 3115 10379 3161 10425
rect 3115 10276 3161 10322
rect 3115 10173 3161 10219
rect 3115 10070 3161 10116
rect 3115 9967 3161 10013
rect 3339 10997 3385 11757
rect 3339 10894 3385 10940
rect 3339 10791 3385 10837
rect 3339 10688 3385 10734
rect 3339 10585 3385 10631
rect 3339 10482 3385 10528
rect 3339 10379 3385 10425
rect 3339 10276 3385 10322
rect 3339 10173 3385 10219
rect 3339 10070 3385 10116
rect 3339 9967 3385 10013
rect 3563 10997 3609 11757
rect 3563 10894 3609 10940
rect 3563 10791 3609 10837
rect 3563 10688 3609 10734
rect 3563 10585 3609 10631
rect 3563 10482 3609 10528
rect 3563 10379 3609 10425
rect 3563 10276 3609 10322
rect 3563 10173 3609 10219
rect 3563 10070 3609 10116
rect 3563 9967 3609 10013
rect 3787 10997 3833 11757
rect 3787 10894 3833 10940
rect 3787 10791 3833 10837
rect 3787 10688 3833 10734
rect 3787 10585 3833 10631
rect 3787 10482 3833 10528
rect 3787 10379 3833 10425
rect 3787 10276 3833 10322
rect 3787 10173 3833 10219
rect 3787 10070 3833 10116
rect 3787 9967 3833 10013
rect 4011 10997 4057 11757
rect 4011 10894 4057 10940
rect 4011 10791 4057 10837
rect 4011 10688 4057 10734
rect 4011 10585 4057 10631
rect 4011 10482 4057 10528
rect 4011 10379 4057 10425
rect 4011 10276 4057 10322
rect 4011 10173 4057 10219
rect 4011 10070 4057 10116
rect 4011 9967 4057 10013
rect 4235 10997 4281 11757
rect 4235 10894 4281 10940
rect 4235 10791 4281 10837
rect 4235 10688 4281 10734
rect 4235 10585 4281 10631
rect 4235 10482 4281 10528
rect 4235 10379 4281 10425
rect 4235 10276 4281 10322
rect 4235 10173 4281 10219
rect 4235 10070 4281 10116
rect 4235 9967 4281 10013
rect 4459 10997 4505 11757
rect 4459 10894 4505 10940
rect 4459 10791 4505 10837
rect 4459 10688 4505 10734
rect 4459 10585 4505 10631
rect 4459 10482 4505 10528
rect 4459 10379 4505 10425
rect 4459 10276 4505 10322
rect 4459 10173 4505 10219
rect 4459 10070 4505 10116
rect 4459 9967 4505 10013
rect 4683 10997 4729 11757
rect 4683 10894 4729 10940
rect 4683 10791 4729 10837
rect 4683 10688 4729 10734
rect 4683 10585 4729 10631
rect 4683 10482 4729 10528
rect 4683 10379 4729 10425
rect 4683 10276 4729 10322
rect 4683 10173 4729 10219
rect 4683 10070 4729 10116
rect 4683 9967 4729 10013
rect 4907 10997 4953 11757
rect 4907 10894 4953 10940
rect 4907 10791 4953 10837
rect 4907 10688 4953 10734
rect 4907 10585 4953 10631
rect 4907 10482 4953 10528
rect 4907 10379 4953 10425
rect 4907 10276 4953 10322
rect 4907 10173 4953 10219
rect 4907 10070 4953 10116
rect 4907 9967 4953 10013
rect 5131 10997 5177 11757
rect 5131 10894 5177 10940
rect 5131 10791 5177 10837
rect 5131 10688 5177 10734
rect 5131 10585 5177 10631
rect 5131 10482 5177 10528
rect 5131 10379 5177 10425
rect 5131 10276 5177 10322
rect 5131 10173 5177 10219
rect 5131 10070 5177 10116
rect 5131 9967 5177 10013
rect 5355 10997 5401 11757
rect 5355 10894 5401 10940
rect 5355 10791 5401 10837
rect 5355 10688 5401 10734
rect 5355 10585 5401 10631
rect 5355 10482 5401 10528
rect 5355 10379 5401 10425
rect 5355 10276 5401 10322
rect 5355 10173 5401 10219
rect 5355 10070 5401 10116
rect 5355 9967 5401 10013
rect 5579 10997 5625 11757
rect 5579 10894 5625 10940
rect 5579 10791 5625 10837
rect 5579 10688 5625 10734
rect 5579 10585 5625 10631
rect 5579 10482 5625 10528
rect 5579 10379 5625 10425
rect 5579 10276 5625 10322
rect 5579 10173 5625 10219
rect 5579 10070 5625 10116
rect 5579 9967 5625 10013
rect 5803 10997 5849 11757
rect 5803 10894 5849 10940
rect 5803 10791 5849 10837
rect 5803 10688 5849 10734
rect 5803 10585 5849 10631
rect 5803 10482 5849 10528
rect 5803 10379 5849 10425
rect 5803 10276 5849 10322
rect 5803 10173 5849 10219
rect 5803 10070 5849 10116
rect 5803 9967 5849 10013
rect 6027 10997 6073 11757
rect 6027 10894 6073 10940
rect 6027 10791 6073 10837
rect 6027 10688 6073 10734
rect 6027 10585 6073 10631
rect 6027 10482 6073 10528
rect 6027 10379 6073 10425
rect 6027 10276 6073 10322
rect 6027 10173 6073 10219
rect 6027 10070 6073 10116
rect 6027 9967 6073 10013
rect 6251 10997 6297 11757
rect 6251 10894 6297 10940
rect 6251 10791 6297 10837
rect 6251 10688 6297 10734
rect 6251 10585 6297 10631
rect 6251 10482 6297 10528
rect 6251 10379 6297 10425
rect 6251 10276 6297 10322
rect 6251 10173 6297 10219
rect 6251 10070 6297 10116
rect 6251 9967 6297 10013
rect 6475 10997 6521 11757
rect 6475 10894 6521 10940
rect 6475 10791 6521 10837
rect 6475 10688 6521 10734
rect 6475 10585 6521 10631
rect 6475 10482 6521 10528
rect 6475 10379 6521 10425
rect 6475 10276 6521 10322
rect 6475 10173 6521 10219
rect 6475 10070 6521 10116
rect 6475 9967 6521 10013
rect 6699 10997 6745 11757
rect 6699 10894 6745 10940
rect 6699 10791 6745 10837
rect 6699 10688 6745 10734
rect 6699 10585 6745 10631
rect 6699 10482 6745 10528
rect 6699 10379 6745 10425
rect 6699 10276 6745 10322
rect 6699 10173 6745 10219
rect 6699 10070 6745 10116
rect 6699 9967 6745 10013
rect 6923 10997 6969 11757
rect 6923 10894 6969 10940
rect 6923 10791 6969 10837
rect 6923 10688 6969 10734
rect 6923 10585 6969 10631
rect 6923 10482 6969 10528
rect 6923 10379 6969 10425
rect 6923 10276 6969 10322
rect 6923 10173 6969 10219
rect 6923 10070 6969 10116
rect 6923 9967 6969 10013
rect 7147 10997 7193 11757
rect 7147 10894 7193 10940
rect 7147 10791 7193 10837
rect 7147 10688 7193 10734
rect 7147 10585 7193 10631
rect 7147 10482 7193 10528
rect 7147 10379 7193 10425
rect 7147 10276 7193 10322
rect 7147 10173 7193 10219
rect 7147 10070 7193 10116
rect 7147 9967 7193 10013
rect 7371 10997 7417 11757
rect 7371 10894 7417 10940
rect 7371 10791 7417 10837
rect 7371 10688 7417 10734
rect 7371 10585 7417 10631
rect 7371 10482 7417 10528
rect 7371 10379 7417 10425
rect 7371 10276 7417 10322
rect 7371 10173 7417 10219
rect 7371 10070 7417 10116
rect 7371 9967 7417 10013
rect 7595 10997 7641 11757
rect 7595 10894 7641 10940
rect 7595 10791 7641 10837
rect 7595 10688 7641 10734
rect 7595 10585 7641 10631
rect 7595 10482 7641 10528
rect 7595 10379 7641 10425
rect 7595 10276 7641 10322
rect 7595 10173 7641 10219
rect 7595 10070 7641 10116
rect 7595 9967 7641 10013
rect 7819 10997 7865 11757
rect 7819 10894 7865 10940
rect 7819 10791 7865 10837
rect 7819 10688 7865 10734
rect 7819 10585 7865 10631
rect 7819 10482 7865 10528
rect 7819 10379 7865 10425
rect 7819 10276 7865 10322
rect 7819 10173 7865 10219
rect 7819 10070 7865 10116
rect 7819 9967 7865 10013
rect 8043 10997 8089 11757
rect 8043 10894 8089 10940
rect 8043 10791 8089 10837
rect 8043 10688 8089 10734
rect 8043 10585 8089 10631
rect 8043 10482 8089 10528
rect 8043 10379 8089 10425
rect 8043 10276 8089 10322
rect 8043 10173 8089 10219
rect 8043 10070 8089 10116
rect 8043 9967 8089 10013
rect 8267 10997 8313 11757
rect 8267 10894 8313 10940
rect 8267 10791 8313 10837
rect 8267 10688 8313 10734
rect 8267 10585 8313 10631
rect 8267 10482 8313 10528
rect 8267 10379 8313 10425
rect 8267 10276 8313 10322
rect 8267 10173 8313 10219
rect 8267 10070 8313 10116
rect 8267 9967 8313 10013
rect 8491 10997 8537 11757
rect 8491 10894 8537 10940
rect 8491 10791 8537 10837
rect 8491 10688 8537 10734
rect 8491 10585 8537 10631
rect 8491 10482 8537 10528
rect 8491 10379 8537 10425
rect 8491 10276 8537 10322
rect 8491 10173 8537 10219
rect 8491 10070 8537 10116
rect 8491 9967 8537 10013
rect 8715 10997 8761 11757
rect 8715 10894 8761 10940
rect 8715 10791 8761 10837
rect 8715 10688 8761 10734
rect 8715 10585 8761 10631
rect 8715 10482 8761 10528
rect 8715 10379 8761 10425
rect 8715 10276 8761 10322
rect 8715 10173 8761 10219
rect 8715 10070 8761 10116
rect 8715 9967 8761 10013
rect 8939 10997 8985 11757
rect 8939 10894 8985 10940
rect 8939 10791 8985 10837
rect 8939 10688 8985 10734
rect 8939 10585 8985 10631
rect 8939 10482 8985 10528
rect 8939 10379 8985 10425
rect 8939 10276 8985 10322
rect 8939 10173 8985 10219
rect 8939 10070 8985 10116
rect 8939 9967 8985 10013
rect 9163 10997 9209 11757
rect 9163 10894 9209 10940
rect 9163 10791 9209 10837
rect 9163 10688 9209 10734
rect 9163 10585 9209 10631
rect 9163 10482 9209 10528
rect 9163 10379 9209 10425
rect 9163 10276 9209 10322
rect 9163 10173 9209 10219
rect 9163 10070 9209 10116
rect 9163 9967 9209 10013
rect 9387 10997 9433 11757
rect 9387 10894 9433 10940
rect 9387 10791 9433 10837
rect 9387 10688 9433 10734
rect 9387 10585 9433 10631
rect 9387 10482 9433 10528
rect 9387 10379 9433 10425
rect 9387 10276 9433 10322
rect 9387 10173 9433 10219
rect 9387 10070 9433 10116
rect 9387 9967 9433 10013
rect 9611 10997 9657 11757
rect 9611 10894 9657 10940
rect 9611 10791 9657 10837
rect 9611 10688 9657 10734
rect 9611 10585 9657 10631
rect 9611 10482 9657 10528
rect 9611 10379 9657 10425
rect 9611 10276 9657 10322
rect 9611 10173 9657 10219
rect 9611 10070 9657 10116
rect 9611 9967 9657 10013
rect 9835 10997 9881 11757
rect 9835 10894 9881 10940
rect 9835 10791 9881 10837
rect 9835 10688 9881 10734
rect 9835 10585 9881 10631
rect 9835 10482 9881 10528
rect 9835 10379 9881 10425
rect 9835 10276 9881 10322
rect 9835 10173 9881 10219
rect 9835 10070 9881 10116
rect 9835 9967 9881 10013
rect 10059 10997 10105 11757
rect 10059 10894 10105 10940
rect 10059 10791 10105 10837
rect 10059 10688 10105 10734
rect 10059 10585 10105 10631
rect 10059 10482 10105 10528
rect 10059 10379 10105 10425
rect 10059 10276 10105 10322
rect 10059 10173 10105 10219
rect 10059 10070 10105 10116
rect 10059 9967 10105 10013
rect 10283 10997 10329 11757
rect 10283 10894 10329 10940
rect 10283 10791 10329 10837
rect 10283 10688 10329 10734
rect 10283 10585 10329 10631
rect 10283 10482 10329 10528
rect 10283 10379 10329 10425
rect 10283 10276 10329 10322
rect 10283 10173 10329 10219
rect 10283 10070 10329 10116
rect 10283 9967 10329 10013
rect 10507 10997 10553 11757
rect 10507 10894 10553 10940
rect 10507 10791 10553 10837
rect 10507 10688 10553 10734
rect 10507 10585 10553 10631
rect 10507 10482 10553 10528
rect 10507 10379 10553 10425
rect 10507 10276 10553 10322
rect 10507 10173 10553 10219
rect 10507 10070 10553 10116
rect 10507 9967 10553 10013
rect 10731 10997 10777 11757
rect 10731 10894 10777 10940
rect 10731 10791 10777 10837
rect 10731 10688 10777 10734
rect 10731 10585 10777 10631
rect 10731 10482 10777 10528
rect 10731 10379 10777 10425
rect 10731 10276 10777 10322
rect 10731 10173 10777 10219
rect 10731 10070 10777 10116
rect 10731 9967 10777 10013
rect 10955 10997 11001 11757
rect 10955 10894 11001 10940
rect 10955 10791 11001 10837
rect 10955 10688 11001 10734
rect 10955 10585 11001 10631
rect 10955 10482 11001 10528
rect 10955 10379 11001 10425
rect 10955 10276 11001 10322
rect 10955 10173 11001 10219
rect 10955 10070 11001 10116
rect 10955 9967 11001 10013
rect 11179 10997 11225 11757
rect 11179 10894 11225 10940
rect 11179 10791 11225 10837
rect 11179 10688 11225 10734
rect 11179 10585 11225 10631
rect 11179 10482 11225 10528
rect 11179 10379 11225 10425
rect 11179 10276 11225 10322
rect 11179 10173 11225 10219
rect 11179 10070 11225 10116
rect 11179 9967 11225 10013
rect 11403 10997 11449 11757
rect 11403 10894 11449 10940
rect 11403 10791 11449 10837
rect 11403 10688 11449 10734
rect 11403 10585 11449 10631
rect 11403 10482 11449 10528
rect 11403 10379 11449 10425
rect 11403 10276 11449 10322
rect 11403 10173 11449 10219
rect 11403 10070 11449 10116
rect 11403 9967 11449 10013
rect 11627 10997 11673 11757
rect 11627 10894 11673 10940
rect 11627 10791 11673 10837
rect 11627 10688 11673 10734
rect 11627 10585 11673 10631
rect 11627 10482 11673 10528
rect 11627 10379 11673 10425
rect 11627 10276 11673 10322
rect 11627 10173 11673 10219
rect 11627 10070 11673 10116
rect 11627 9967 11673 10013
rect 11851 10997 11897 11757
rect 11851 10894 11897 10940
rect 11851 10791 11897 10837
rect 11851 10688 11897 10734
rect 11851 10585 11897 10631
rect 11851 10482 11897 10528
rect 11851 10379 11897 10425
rect 11851 10276 11897 10322
rect 11851 10173 11897 10219
rect 11851 10070 11897 10116
rect 11851 9967 11897 10013
rect 12075 10997 12121 11757
rect 12075 10894 12121 10940
rect 12075 10791 12121 10837
rect 12075 10688 12121 10734
rect 12075 10585 12121 10631
rect 12075 10482 12121 10528
rect 12075 10379 12121 10425
rect 12075 10276 12121 10322
rect 12075 10173 12121 10219
rect 12075 10070 12121 10116
rect 12075 9967 12121 10013
rect 12299 10997 12345 11757
rect 12299 10894 12345 10940
rect 12299 10791 12345 10837
rect 12299 10688 12345 10734
rect 12299 10585 12345 10631
rect 12299 10482 12345 10528
rect 12299 10379 12345 10425
rect 12299 10276 12345 10322
rect 12299 10173 12345 10219
rect 12299 10070 12345 10116
rect 12299 9967 12345 10013
rect 12523 10997 12569 11757
rect 12523 10894 12569 10940
rect 12523 10791 12569 10837
rect 12523 10688 12569 10734
rect 12523 10585 12569 10631
rect 12523 10482 12569 10528
rect 12523 10379 12569 10425
rect 12523 10276 12569 10322
rect 12523 10173 12569 10219
rect 12523 10070 12569 10116
rect 12523 9967 12569 10013
rect 12747 10997 12793 11757
rect 12747 10894 12793 10940
rect 12747 10791 12793 10837
rect 12747 10688 12793 10734
rect 12747 10585 12793 10631
rect 12747 10482 12793 10528
rect 12747 10379 12793 10425
rect 12747 10276 12793 10322
rect 12747 10173 12793 10219
rect 12747 10070 12793 10116
rect 12747 9967 12793 10013
rect 12971 10997 13017 11757
rect 12971 10894 13017 10940
rect 12971 10791 13017 10837
rect 12971 10688 13017 10734
rect 12971 10585 13017 10631
rect 12971 10482 13017 10528
rect 12971 10379 13017 10425
rect 12971 10276 13017 10322
rect 12971 10173 13017 10219
rect 12971 10070 13017 10116
rect 12971 9967 13017 10013
rect 13195 10997 13241 11757
rect 13195 10894 13241 10940
rect 13195 10791 13241 10837
rect 13195 10688 13241 10734
rect 13195 10585 13241 10631
rect 13195 10482 13241 10528
rect 13195 10379 13241 10425
rect 13195 10276 13241 10322
rect 13195 10173 13241 10219
rect 13195 10070 13241 10116
rect 13195 9967 13241 10013
rect 13419 10997 13465 11757
rect 13419 10894 13465 10940
rect 13419 10791 13465 10837
rect 13419 10688 13465 10734
rect 13419 10585 13465 10631
rect 13419 10482 13465 10528
rect 13419 10379 13465 10425
rect 13419 10276 13465 10322
rect 13419 10173 13465 10219
rect 13419 10070 13465 10116
rect 13419 9967 13465 10013
rect 13643 10997 13689 11757
rect 13643 10894 13689 10940
rect 13643 10791 13689 10837
rect 13643 10688 13689 10734
rect 13643 10585 13689 10631
rect 13643 10482 13689 10528
rect 13643 10379 13689 10425
rect 13643 10276 13689 10322
rect 13643 10173 13689 10219
rect 13643 10070 13689 10116
rect 13643 9967 13689 10013
rect 13867 10997 13913 11757
rect 13867 10894 13913 10940
rect 13867 10791 13913 10837
rect 13867 10688 13913 10734
rect 13867 10585 13913 10631
rect 13867 10482 13913 10528
rect 13867 10379 13913 10425
rect 13867 10276 13913 10322
rect 13867 10173 13913 10219
rect 13867 10070 13913 10116
rect 13867 9967 13913 10013
rect 14091 10997 14137 11757
rect 14091 10894 14137 10940
rect 14091 10791 14137 10837
rect 14091 10688 14137 10734
rect 14091 10585 14137 10631
rect 14091 10482 14137 10528
rect 14091 10379 14137 10425
rect 14091 10276 14137 10322
rect 14091 10173 14137 10219
rect 14091 10070 14137 10116
rect 14091 9967 14137 10013
rect 14315 10997 14361 11757
rect 14315 10894 14361 10940
rect 14315 10791 14361 10837
rect 14315 10688 14361 10734
rect 14315 10585 14361 10631
rect 14315 10482 14361 10528
rect 14315 10379 14361 10425
rect 14315 10276 14361 10322
rect 14315 10173 14361 10219
rect 14315 10070 14361 10116
rect 14315 9967 14361 10013
rect 14539 10997 14585 11757
rect 14539 10894 14585 10940
rect 14539 10791 14585 10837
rect 14539 10688 14585 10734
rect 14539 10585 14585 10631
rect 14539 10482 14585 10528
rect 14539 10379 14585 10425
rect 14539 10276 14585 10322
rect 14539 10173 14585 10219
rect 14539 10070 14585 10116
rect 14539 9967 14585 10013
rect 14763 10997 14809 11757
rect 14763 10894 14809 10940
rect 14763 10791 14809 10837
rect 14763 10688 14809 10734
rect 14763 10585 14809 10631
rect 14763 10482 14809 10528
rect 14763 10379 14809 10425
rect 14763 10276 14809 10322
rect 14763 10173 14809 10219
rect 14763 10070 14809 10116
rect 14763 9967 14809 10013
rect 14987 10997 15033 11757
rect 14987 10894 15033 10940
rect 14987 10791 15033 10837
rect 14987 10688 15033 10734
rect 14987 10585 15033 10631
rect 14987 10482 15033 10528
rect 14987 10379 15033 10425
rect 14987 10276 15033 10322
rect 14987 10173 15033 10219
rect 14987 10070 15033 10116
rect 14987 9967 15033 10013
rect 15211 10997 15257 11757
rect 15211 10894 15257 10940
rect 15211 10791 15257 10837
rect 15211 10688 15257 10734
rect 15211 10585 15257 10631
rect 15211 10482 15257 10528
rect 15211 10379 15257 10425
rect 15211 10276 15257 10322
rect 15211 10173 15257 10219
rect 15211 10070 15257 10116
rect 15211 9967 15257 10013
rect 15435 10997 15481 11757
rect 15435 10894 15481 10940
rect 15435 10791 15481 10837
rect 15435 10688 15481 10734
rect 15435 10585 15481 10631
rect 15435 10482 15481 10528
rect 15435 10379 15481 10425
rect 15435 10276 15481 10322
rect 15435 10173 15481 10219
rect 15435 10070 15481 10116
rect 15435 9967 15481 10013
rect 15659 10997 15705 11757
rect 15659 10894 15705 10940
rect 15659 10791 15705 10837
rect 15659 10688 15705 10734
rect 15659 10585 15705 10631
rect 15659 10482 15705 10528
rect 15659 10379 15705 10425
rect 15659 10276 15705 10322
rect 15659 10173 15705 10219
rect 15659 10070 15705 10116
rect 15659 9967 15705 10013
rect 15883 10997 15929 11757
rect 15883 10894 15929 10940
rect 15883 10791 15929 10837
rect 15883 10688 15929 10734
rect 15883 10585 15929 10631
rect 15883 10482 15929 10528
rect 15883 10379 15929 10425
rect 15883 10276 15929 10322
rect 15883 10173 15929 10219
rect 15883 10070 15929 10116
rect 15883 9967 15929 10013
rect 16107 10997 16153 11757
rect 16107 10894 16153 10940
rect 16107 10791 16153 10837
rect 16107 10688 16153 10734
rect 16107 10585 16153 10631
rect 16107 10482 16153 10528
rect 16107 10379 16153 10425
rect 16107 10276 16153 10322
rect 16107 10173 16153 10219
rect 16107 10070 16153 10116
rect 16107 9967 16153 10013
rect 16331 10997 16377 11757
rect 16331 10894 16377 10940
rect 16331 10791 16377 10837
rect 16331 10688 16377 10734
rect 16331 10585 16377 10631
rect 16331 10482 16377 10528
rect 16331 10379 16377 10425
rect 16331 10276 16377 10322
rect 16331 10173 16377 10219
rect 16331 10070 16377 10116
rect 16331 9967 16377 10013
rect 16555 10997 16601 11757
rect 16555 10894 16601 10940
rect 16555 10791 16601 10837
rect 16555 10688 16601 10734
rect 16555 10585 16601 10631
rect 16555 10482 16601 10528
rect 16555 10379 16601 10425
rect 16555 10276 16601 10322
rect 16555 10173 16601 10219
rect 16555 10070 16601 10116
rect 16555 9967 16601 10013
rect 16779 10997 16825 11757
rect 16779 10894 16825 10940
rect 16779 10791 16825 10837
rect 16779 10688 16825 10734
rect 16779 10585 16825 10631
rect 16779 10482 16825 10528
rect 16779 10379 16825 10425
rect 16779 10276 16825 10322
rect 16779 10173 16825 10219
rect 16779 10070 16825 10116
rect 16779 9967 16825 10013
rect 17003 10997 17049 11757
rect 17003 10894 17049 10940
rect 17003 10791 17049 10837
rect 17003 10688 17049 10734
rect 17003 10585 17049 10631
rect 17003 10482 17049 10528
rect 17003 10379 17049 10425
rect 17003 10276 17049 10322
rect 17003 10173 17049 10219
rect 17003 10070 17049 10116
rect 17003 9967 17049 10013
rect 17227 10997 17273 11757
rect 17227 10894 17273 10940
rect 17227 10791 17273 10837
rect 17227 10688 17273 10734
rect 17227 10585 17273 10631
rect 17227 10482 17273 10528
rect 17227 10379 17273 10425
rect 17227 10276 17273 10322
rect 17227 10173 17273 10219
rect 17227 10070 17273 10116
rect 17227 9967 17273 10013
rect 17451 10997 17497 11757
rect 17451 10894 17497 10940
rect 17451 10791 17497 10837
rect 17451 10688 17497 10734
rect 17451 10585 17497 10631
rect 17451 10482 17497 10528
rect 17451 10379 17497 10425
rect 17451 10276 17497 10322
rect 17451 10173 17497 10219
rect 17451 10070 17497 10116
rect 17451 9967 17497 10013
rect 17675 10997 17721 11757
rect 17675 10894 17721 10940
rect 17675 10791 17721 10837
rect 17675 10688 17721 10734
rect 17675 10585 17721 10631
rect 17675 10482 17721 10528
rect 17675 10379 17721 10425
rect 17675 10276 17721 10322
rect 17675 10173 17721 10219
rect 17675 10070 17721 10116
rect 17675 9967 17721 10013
rect 17899 10997 17945 11757
rect 17899 10894 17945 10940
rect 17899 10791 17945 10837
rect 17899 10688 17945 10734
rect 17899 10585 17945 10631
rect 17899 10482 17945 10528
rect 17899 10379 17945 10425
rect 17899 10276 17945 10322
rect 17899 10173 17945 10219
rect 17899 10070 17945 10116
rect 17899 9967 17945 10013
rect 18123 10997 18169 11757
rect 18123 10894 18169 10940
rect 18123 10791 18169 10837
rect 18123 10688 18169 10734
rect 18123 10585 18169 10631
rect 18123 10482 18169 10528
rect 18123 10379 18169 10425
rect 18123 10276 18169 10322
rect 18123 10173 18169 10219
rect 18123 10070 18169 10116
rect 18123 9967 18169 10013
rect 18347 10997 18393 11757
rect 18347 10894 18393 10940
rect 18347 10791 18393 10837
rect 18347 10688 18393 10734
rect 18347 10585 18393 10631
rect 18347 10482 18393 10528
rect 18347 10379 18393 10425
rect 18347 10276 18393 10322
rect 18347 10173 18393 10219
rect 18347 10070 18393 10116
rect 18347 9967 18393 10013
rect 18571 10997 18617 11757
rect 18571 10894 18617 10940
rect 18571 10791 18617 10837
rect 18571 10688 18617 10734
rect 18571 10585 18617 10631
rect 18571 10482 18617 10528
rect 18571 10379 18617 10425
rect 18571 10276 18617 10322
rect 18571 10173 18617 10219
rect 18571 10070 18617 10116
rect 18571 9967 18617 10013
rect 18795 10997 18841 11757
rect 18795 10894 18841 10940
rect 18795 10791 18841 10837
rect 18795 10688 18841 10734
rect 18795 10585 18841 10631
rect 18795 10482 18841 10528
rect 18795 10379 18841 10425
rect 18795 10276 18841 10322
rect 18795 10173 18841 10219
rect 18795 10070 18841 10116
rect 18795 9967 18841 10013
rect 19019 10997 19065 11757
rect 19019 10894 19065 10940
rect 19019 10791 19065 10837
rect 19019 10688 19065 10734
rect 19019 10585 19065 10631
rect 19019 10482 19065 10528
rect 19019 10379 19065 10425
rect 19019 10276 19065 10322
rect 19019 10173 19065 10219
rect 19019 10070 19065 10116
rect 19019 9967 19065 10013
rect 19243 10997 19289 11757
rect 19243 10894 19289 10940
rect 19243 10791 19289 10837
rect 19243 10688 19289 10734
rect 19243 10585 19289 10631
rect 19243 10482 19289 10528
rect 19243 10379 19289 10425
rect 19243 10276 19289 10322
rect 19243 10173 19289 10219
rect 19243 10070 19289 10116
rect 19243 9967 19289 10013
rect 19467 10997 19513 11757
rect 19467 10894 19513 10940
rect 19467 10791 19513 10837
rect 19467 10688 19513 10734
rect 19467 10585 19513 10631
rect 19467 10482 19513 10528
rect 19467 10379 19513 10425
rect 19467 10276 19513 10322
rect 19467 10173 19513 10219
rect 19467 10070 19513 10116
rect 19467 9967 19513 10013
rect 19691 10997 19737 11757
rect 19691 10894 19737 10940
rect 19691 10791 19737 10837
rect 19691 10688 19737 10734
rect 19691 10585 19737 10631
rect 19691 10482 19737 10528
rect 19691 10379 19737 10425
rect 19691 10276 19737 10322
rect 19691 10173 19737 10219
rect 19691 10070 19737 10116
rect 19691 9967 19737 10013
rect 19915 10997 19961 11757
rect 19915 10894 19961 10940
rect 19915 10791 19961 10837
rect 19915 10688 19961 10734
rect 19915 10585 19961 10631
rect 19915 10482 19961 10528
rect 19915 10379 19961 10425
rect 19915 10276 19961 10322
rect 19915 10173 19961 10219
rect 19915 10070 19961 10116
rect 19915 9967 19961 10013
rect 2621 9106 2667 9152
rect 2621 9002 2667 9048
rect 2621 8898 2667 8944
rect 2621 8794 2667 8840
rect 2621 8690 2667 8736
rect 2621 8585 2667 8631
rect 2621 8480 2667 8526
rect 2621 8375 2667 8421
rect 2621 8270 2667 8316
rect 2845 9106 2891 9152
rect 2845 9002 2891 9048
rect 2845 8898 2891 8944
rect 2845 8794 2891 8840
rect 2845 8690 2891 8736
rect 2845 8585 2891 8631
rect 2845 8480 2891 8526
rect 2845 8375 2891 8421
rect 2845 8270 2891 8316
rect 3135 9106 3181 9152
rect 3135 9002 3181 9048
rect 3135 8898 3181 8944
rect 3135 8794 3181 8840
rect 3135 8690 3181 8736
rect 3135 8585 3181 8631
rect 3135 8480 3181 8526
rect 3135 8375 3181 8421
rect 3135 8270 3181 8316
rect 3359 9106 3405 9152
rect 3359 9002 3405 9048
rect 3359 8898 3405 8944
rect 3359 8794 3405 8840
rect 3359 8690 3405 8736
rect 3359 8585 3405 8631
rect 3359 8480 3405 8526
rect 4312 9106 4358 9152
rect 4312 9002 4358 9048
rect 4312 8898 4358 8944
rect 4312 8794 4358 8840
rect 4312 8690 4358 8736
rect 4312 8585 4358 8631
rect 3359 8375 3405 8421
rect 3359 8270 3405 8316
rect 4312 8480 4358 8526
rect 4312 8375 4358 8421
rect 4312 8270 4358 8316
rect 4536 9106 4582 9152
rect 4536 9002 4582 9048
rect 4536 8898 4582 8944
rect 4536 8794 4582 8840
rect 4536 8690 4582 8736
rect 4536 8585 4582 8631
rect 4536 8480 4582 8526
rect 4536 8375 4582 8421
rect 4536 8270 4582 8316
rect 4826 9106 4872 9152
rect 4826 9002 4872 9048
rect 4826 8898 4872 8944
rect 4826 8794 4872 8840
rect 4826 8690 4872 8736
rect 4826 8585 4872 8631
rect 4826 8480 4872 8526
rect 4826 8375 4872 8421
rect 4826 8270 4872 8316
rect 5050 9106 5096 9152
rect 5050 9002 5096 9048
rect 5050 8898 5096 8944
rect 5050 8794 5096 8840
rect 5050 8690 5096 8736
rect 5050 8585 5096 8631
rect 5050 8480 5096 8526
rect 6003 9106 6049 9152
rect 6003 9002 6049 9048
rect 6003 8898 6049 8944
rect 6003 8794 6049 8840
rect 6003 8690 6049 8736
rect 6003 8585 6049 8631
rect 5050 8375 5096 8421
rect 5050 8270 5096 8316
rect 6003 8480 6049 8526
rect 6003 8375 6049 8421
rect 6003 8270 6049 8316
rect 6227 9106 6273 9152
rect 6227 9002 6273 9048
rect 6227 8898 6273 8944
rect 6227 8794 6273 8840
rect 6227 8690 6273 8736
rect 6227 8585 6273 8631
rect 6227 8480 6273 8526
rect 6227 8375 6273 8421
rect 6227 8270 6273 8316
rect 6517 9106 6563 9152
rect 6517 9002 6563 9048
rect 6517 8898 6563 8944
rect 6517 8794 6563 8840
rect 6517 8690 6563 8736
rect 6517 8585 6563 8631
rect 6517 8480 6563 8526
rect 6517 8375 6563 8421
rect 6517 8270 6563 8316
rect 6741 9106 6787 9152
rect 6741 9002 6787 9048
rect 6741 8898 6787 8944
rect 6741 8794 6787 8840
rect 6741 8690 6787 8736
rect 6741 8585 6787 8631
rect 7450 8962 7496 9008
rect 7450 8834 7496 8880
rect 7450 8707 7496 8753
rect 7450 8580 7496 8626
rect 7674 8962 7720 9008
rect 7674 8834 7720 8880
rect 7674 8707 7720 8753
rect 7674 8580 7720 8626
rect 7898 8962 7944 9008
rect 7898 8834 7944 8880
rect 7898 8707 7944 8753
rect 7898 8580 7944 8626
rect 8122 8962 8168 9008
rect 8122 8834 8168 8880
rect 8122 8707 8168 8753
rect 8122 8580 8168 8626
rect 8346 8962 8392 9008
rect 8346 8834 8392 8880
rect 8346 8707 8392 8753
rect 8346 8580 8392 8626
rect 8570 8962 8616 9008
rect 8570 8834 8616 8880
rect 8570 8707 8616 8753
rect 8570 8580 8616 8626
rect 8794 8962 8840 9008
rect 8794 8834 8840 8880
rect 8794 8707 8840 8753
rect 8794 8580 8840 8626
rect 9083 8962 9129 9008
rect 9083 8834 9129 8880
rect 9083 8707 9129 8753
rect 9083 8580 9129 8626
rect 9307 8962 9353 9008
rect 9307 8834 9353 8880
rect 9307 8707 9353 8753
rect 9307 8580 9353 8626
rect 9531 8962 9577 9008
rect 9531 8834 9577 8880
rect 9531 8707 9577 8753
rect 9531 8580 9577 8626
rect 9755 8962 9801 9008
rect 9755 8834 9801 8880
rect 9755 8707 9801 8753
rect 9755 8580 9801 8626
rect 9979 8962 10025 9008
rect 9979 8834 10025 8880
rect 9979 8707 10025 8753
rect 9979 8580 10025 8626
rect 10203 8962 10249 9008
rect 10203 8834 10249 8880
rect 10203 8707 10249 8753
rect 10203 8580 10249 8626
rect 10427 8962 10473 9008
rect 10427 8834 10473 8880
rect 10427 8707 10473 8753
rect 10427 8580 10473 8626
rect 10717 8962 10763 9008
rect 10717 8834 10763 8880
rect 10717 8707 10763 8753
rect 10717 8580 10763 8626
rect 10941 8962 10987 9008
rect 10941 8834 10987 8880
rect 10941 8707 10987 8753
rect 10941 8580 10987 8626
rect 11165 8962 11211 9008
rect 11165 8834 11211 8880
rect 11165 8707 11211 8753
rect 11165 8580 11211 8626
rect 11389 8962 11435 9008
rect 11389 8834 11435 8880
rect 11389 8707 11435 8753
rect 11389 8580 11435 8626
rect 11613 8962 11659 9008
rect 11613 8834 11659 8880
rect 11613 8707 11659 8753
rect 11613 8580 11659 8626
rect 11837 8962 11883 9008
rect 11837 8834 11883 8880
rect 11837 8707 11883 8753
rect 11837 8580 11883 8626
rect 12061 8962 12107 9008
rect 12061 8834 12107 8880
rect 12061 8707 12107 8753
rect 12061 8580 12107 8626
rect 12351 8962 12397 9008
rect 12351 8834 12397 8880
rect 12351 8707 12397 8753
rect 12351 8580 12397 8626
rect 12575 8962 12621 9008
rect 12575 8834 12621 8880
rect 12575 8707 12621 8753
rect 12575 8580 12621 8626
rect 12799 8962 12845 9008
rect 12799 8834 12845 8880
rect 12799 8707 12845 8753
rect 12799 8580 12845 8626
rect 13023 8962 13069 9008
rect 13023 8834 13069 8880
rect 13023 8707 13069 8753
rect 13023 8580 13069 8626
rect 13247 8962 13293 9008
rect 13247 8834 13293 8880
rect 13247 8707 13293 8753
rect 13247 8580 13293 8626
rect 13471 8962 13517 9008
rect 13471 8834 13517 8880
rect 13471 8707 13517 8753
rect 13471 8580 13517 8626
rect 13695 8962 13741 9008
rect 13695 8834 13741 8880
rect 13695 8707 13741 8753
rect 13695 8580 13741 8626
rect 6741 8480 6787 8526
rect 6741 8375 6787 8421
rect 6741 8270 6787 8316
rect 7450 3820 7496 3866
rect 7450 3652 7496 3698
rect 7450 3484 7496 3530
rect 7450 3317 7496 3363
rect 7450 3149 7496 3195
rect 7450 2981 7496 3027
rect 7450 2813 7496 2859
rect 7450 2646 7496 2692
rect 8122 3820 8168 3866
rect 8122 3652 8168 3698
rect 8122 3484 8168 3530
rect 8122 3317 8168 3363
rect 8122 3149 8168 3195
rect 8122 2981 8168 3027
rect 8122 2813 8168 2859
rect 8122 2646 8168 2692
rect 8794 3820 8840 3866
rect 8794 3652 8840 3698
rect 8794 3484 8840 3530
rect 8794 3317 8840 3363
rect 8794 3149 8840 3195
rect 8794 2981 8840 3027
rect 8794 2813 8840 2859
rect 8794 2646 8840 2692
rect 9083 3820 9129 3866
rect 9083 3652 9129 3698
rect 9083 3484 9129 3530
rect 9083 3317 9129 3363
rect 9083 3149 9129 3195
rect 9083 2981 9129 3027
rect 9083 2813 9129 2859
rect 9083 2646 9129 2692
rect 9755 3820 9801 3866
rect 9755 3652 9801 3698
rect 9755 3484 9801 3530
rect 9755 3317 9801 3363
rect 9755 3149 9801 3195
rect 9755 2981 9801 3027
rect 9755 2813 9801 2859
rect 9755 2646 9801 2692
rect 10427 3820 10473 3866
rect 10427 3652 10473 3698
rect 10427 3484 10473 3530
rect 10427 3317 10473 3363
rect 10427 3149 10473 3195
rect 10427 2981 10473 3027
rect 10427 2813 10473 2859
rect 10427 2646 10473 2692
rect 10717 3820 10763 3866
rect 10717 3652 10763 3698
rect 10717 3484 10763 3530
rect 10717 3317 10763 3363
rect 10717 3149 10763 3195
rect 10717 2981 10763 3027
rect 10717 2813 10763 2859
rect 10717 2646 10763 2692
rect 11389 3820 11435 3866
rect 11389 3652 11435 3698
rect 11389 3484 11435 3530
rect 11389 3317 11435 3363
rect 11389 3149 11435 3195
rect 11389 2981 11435 3027
rect 11389 2813 11435 2859
rect 11389 2646 11435 2692
rect 12061 3820 12107 3866
rect 12061 3652 12107 3698
rect 12061 3484 12107 3530
rect 12061 3317 12107 3363
rect 12061 3149 12107 3195
rect 12061 2981 12107 3027
rect 12061 2813 12107 2859
rect 12061 2646 12107 2692
rect 12351 3820 12397 3866
rect 12351 3652 12397 3698
rect 12351 3484 12397 3530
rect 12351 3317 12397 3363
rect 12351 3149 12397 3195
rect 12351 2981 12397 3027
rect 12351 2813 12397 2859
rect 12351 2646 12397 2692
rect 13023 3820 13069 3866
rect 13023 3652 13069 3698
rect 13023 3484 13069 3530
rect 13023 3317 13069 3363
rect 13023 3149 13069 3195
rect 13023 2981 13069 3027
rect 13023 2813 13069 2859
rect 13023 2646 13069 2692
rect 13695 3820 13741 3866
rect 13695 3652 13741 3698
rect 13695 3484 13741 3530
rect 13695 3317 13741 3363
rect 13695 3149 13741 3195
rect 13695 2981 13741 3027
rect 13695 2813 13741 2859
rect 13695 2646 13741 2692
rect 9208 1885 9254 1931
rect 7838 1570 7884 1816
rect 8062 1570 8108 1816
rect 9208 1782 9254 1828
rect 9208 1679 9254 1725
rect 9208 1575 9254 1621
rect 9432 1885 9478 1931
rect 9432 1782 9478 1828
rect 9432 1679 9478 1725
rect 9432 1575 9478 1621
rect 9656 1885 9702 1931
rect 9656 1782 9702 1828
rect 9656 1679 9702 1725
rect 9656 1575 9702 1621
<< mvpdiffc >>
rect 1659 27406 1705 27452
rect 1659 27301 1705 27347
rect 1659 27196 1705 27242
rect 1659 27091 1705 27137
rect 1659 26986 1705 27032
rect 1659 26881 1705 26927
rect 1659 26776 1705 26822
rect 1659 26671 1705 26717
rect 1659 26566 1705 26612
rect 1659 26461 1705 26507
rect 1659 26356 1705 26402
rect 1659 26251 1705 26297
rect 1659 26146 1705 26192
rect 1659 26042 1705 26088
rect 1659 25938 1705 25984
rect 1659 25834 1705 25880
rect 1659 25730 1705 25776
rect 1659 25626 1705 25672
rect 1659 25522 1705 25568
rect 1659 25418 1705 25464
rect 1659 25314 1705 25360
rect 1659 25210 1705 25256
rect 1883 27406 1929 27452
rect 1883 27301 1929 27347
rect 1883 27196 1929 27242
rect 1883 27091 1929 27137
rect 1883 26986 1929 27032
rect 1883 26881 1929 26927
rect 1883 26776 1929 26822
rect 1883 26671 1929 26717
rect 1883 26566 1929 26612
rect 1883 26461 1929 26507
rect 1883 26356 1929 26402
rect 1883 26251 1929 26297
rect 1883 26146 1929 26192
rect 1883 26042 1929 26088
rect 1883 25938 1929 25984
rect 1883 25834 1929 25880
rect 1883 25730 1929 25776
rect 1883 25626 1929 25672
rect 1883 25522 1929 25568
rect 1883 25418 1929 25464
rect 1883 25314 1929 25360
rect 1883 25210 1929 25256
rect 2107 27406 2153 27452
rect 2107 27301 2153 27347
rect 2107 27196 2153 27242
rect 2107 27091 2153 27137
rect 2107 26986 2153 27032
rect 2107 26881 2153 26927
rect 2107 26776 2153 26822
rect 2107 26671 2153 26717
rect 2107 26566 2153 26612
rect 2107 26461 2153 26507
rect 2107 26356 2153 26402
rect 2107 26251 2153 26297
rect 2107 26146 2153 26192
rect 2107 26042 2153 26088
rect 2107 25938 2153 25984
rect 2107 25834 2153 25880
rect 2107 25730 2153 25776
rect 2107 25626 2153 25672
rect 2107 25522 2153 25568
rect 2107 25418 2153 25464
rect 2107 25314 2153 25360
rect 2107 25210 2153 25256
rect 2331 27406 2377 27452
rect 2331 27301 2377 27347
rect 2331 27196 2377 27242
rect 2331 27091 2377 27137
rect 2331 26986 2377 27032
rect 2331 26881 2377 26927
rect 2331 26776 2377 26822
rect 2331 26671 2377 26717
rect 2331 26566 2377 26612
rect 2331 26461 2377 26507
rect 2331 26356 2377 26402
rect 2331 26251 2377 26297
rect 2331 26146 2377 26192
rect 2331 26042 2377 26088
rect 2331 25938 2377 25984
rect 2331 25834 2377 25880
rect 2331 25730 2377 25776
rect 2331 25626 2377 25672
rect 2331 25522 2377 25568
rect 2331 25418 2377 25464
rect 2331 25314 2377 25360
rect 2331 25210 2377 25256
rect 2555 27406 2601 27452
rect 2555 27301 2601 27347
rect 2555 27196 2601 27242
rect 2555 27091 2601 27137
rect 2555 26986 2601 27032
rect 2555 26881 2601 26927
rect 2555 26776 2601 26822
rect 2555 26671 2601 26717
rect 2555 26566 2601 26612
rect 2555 26461 2601 26507
rect 2555 26356 2601 26402
rect 2555 26251 2601 26297
rect 2555 26146 2601 26192
rect 2555 26042 2601 26088
rect 2555 25938 2601 25984
rect 2555 25834 2601 25880
rect 2555 25730 2601 25776
rect 2555 25626 2601 25672
rect 2555 25522 2601 25568
rect 2555 25418 2601 25464
rect 2555 25314 2601 25360
rect 2555 25210 2601 25256
rect 2779 27406 2825 27452
rect 2779 27301 2825 27347
rect 2779 27196 2825 27242
rect 2779 27091 2825 27137
rect 2779 26986 2825 27032
rect 2779 26881 2825 26927
rect 2779 26776 2825 26822
rect 2779 26671 2825 26717
rect 2779 26566 2825 26612
rect 2779 26461 2825 26507
rect 2779 26356 2825 26402
rect 2779 26251 2825 26297
rect 2779 26146 2825 26192
rect 2779 26042 2825 26088
rect 2779 25938 2825 25984
rect 2779 25834 2825 25880
rect 2779 25730 2825 25776
rect 2779 25626 2825 25672
rect 2779 25522 2825 25568
rect 2779 25418 2825 25464
rect 2779 25314 2825 25360
rect 2779 25210 2825 25256
rect 3003 27406 3049 27452
rect 3003 27301 3049 27347
rect 3003 27196 3049 27242
rect 3003 27091 3049 27137
rect 3003 26986 3049 27032
rect 3003 26881 3049 26927
rect 3003 26776 3049 26822
rect 3003 26671 3049 26717
rect 3003 26566 3049 26612
rect 3003 26461 3049 26507
rect 3003 26356 3049 26402
rect 3003 26251 3049 26297
rect 3003 26146 3049 26192
rect 3003 26042 3049 26088
rect 3003 25938 3049 25984
rect 3003 25834 3049 25880
rect 3003 25730 3049 25776
rect 3003 25626 3049 25672
rect 3003 25522 3049 25568
rect 3003 25418 3049 25464
rect 3003 25314 3049 25360
rect 3003 25210 3049 25256
rect 3227 27406 3273 27452
rect 3227 27301 3273 27347
rect 3227 27196 3273 27242
rect 3227 27091 3273 27137
rect 3227 26986 3273 27032
rect 3227 26881 3273 26927
rect 3227 26776 3273 26822
rect 3227 26671 3273 26717
rect 3227 26566 3273 26612
rect 3227 26461 3273 26507
rect 3227 26356 3273 26402
rect 3227 26251 3273 26297
rect 3227 26146 3273 26192
rect 3227 26042 3273 26088
rect 3227 25938 3273 25984
rect 3227 25834 3273 25880
rect 3227 25730 3273 25776
rect 3227 25626 3273 25672
rect 3227 25522 3273 25568
rect 3227 25418 3273 25464
rect 3227 25314 3273 25360
rect 3227 25210 3273 25256
rect 3451 27406 3497 27452
rect 3451 27301 3497 27347
rect 3451 27196 3497 27242
rect 3451 27091 3497 27137
rect 3451 26986 3497 27032
rect 3451 26881 3497 26927
rect 3451 26776 3497 26822
rect 3451 26671 3497 26717
rect 3451 26566 3497 26612
rect 3451 26461 3497 26507
rect 3451 26356 3497 26402
rect 3451 26251 3497 26297
rect 3451 26146 3497 26192
rect 3451 26042 3497 26088
rect 3451 25938 3497 25984
rect 3451 25834 3497 25880
rect 3451 25730 3497 25776
rect 3451 25626 3497 25672
rect 3451 25522 3497 25568
rect 3451 25418 3497 25464
rect 3451 25314 3497 25360
rect 3451 25210 3497 25256
rect 3675 27406 3721 27452
rect 3675 27301 3721 27347
rect 3675 27196 3721 27242
rect 3675 27091 3721 27137
rect 3675 26986 3721 27032
rect 3675 26881 3721 26927
rect 3675 26776 3721 26822
rect 3675 26671 3721 26717
rect 3675 26566 3721 26612
rect 3675 26461 3721 26507
rect 3675 26356 3721 26402
rect 3675 26251 3721 26297
rect 3675 26146 3721 26192
rect 3675 26042 3721 26088
rect 3675 25938 3721 25984
rect 3675 25834 3721 25880
rect 3675 25730 3721 25776
rect 3675 25626 3721 25672
rect 3675 25522 3721 25568
rect 3675 25418 3721 25464
rect 3675 25314 3721 25360
rect 3675 25210 3721 25256
rect 3899 27406 3945 27452
rect 3899 27301 3945 27347
rect 3899 27196 3945 27242
rect 3899 27091 3945 27137
rect 3899 26986 3945 27032
rect 3899 26881 3945 26927
rect 3899 26776 3945 26822
rect 3899 26671 3945 26717
rect 3899 26566 3945 26612
rect 3899 26461 3945 26507
rect 3899 26356 3945 26402
rect 3899 26251 3945 26297
rect 3899 26146 3945 26192
rect 3899 26042 3945 26088
rect 3899 25938 3945 25984
rect 3899 25834 3945 25880
rect 3899 25730 3945 25776
rect 3899 25626 3945 25672
rect 3899 25522 3945 25568
rect 3899 25418 3945 25464
rect 3899 25314 3945 25360
rect 3899 25210 3945 25256
rect 4123 27406 4169 27452
rect 4123 27301 4169 27347
rect 4123 27196 4169 27242
rect 4123 27091 4169 27137
rect 4123 26986 4169 27032
rect 4123 26881 4169 26927
rect 4123 26776 4169 26822
rect 4123 26671 4169 26717
rect 4123 26566 4169 26612
rect 4123 26461 4169 26507
rect 4123 26356 4169 26402
rect 4123 26251 4169 26297
rect 4123 26146 4169 26192
rect 4123 26042 4169 26088
rect 4123 25938 4169 25984
rect 4123 25834 4169 25880
rect 4123 25730 4169 25776
rect 4123 25626 4169 25672
rect 4123 25522 4169 25568
rect 4123 25418 4169 25464
rect 4123 25314 4169 25360
rect 4123 25210 4169 25256
rect 4347 27406 4393 27452
rect 4347 27301 4393 27347
rect 4347 27196 4393 27242
rect 4347 27091 4393 27137
rect 4347 26986 4393 27032
rect 4347 26881 4393 26927
rect 4347 26776 4393 26822
rect 4347 26671 4393 26717
rect 4347 26566 4393 26612
rect 4347 26461 4393 26507
rect 4347 26356 4393 26402
rect 4347 26251 4393 26297
rect 4347 26146 4393 26192
rect 4347 26042 4393 26088
rect 4347 25938 4393 25984
rect 4347 25834 4393 25880
rect 4347 25730 4393 25776
rect 4347 25626 4393 25672
rect 4347 25522 4393 25568
rect 4347 25418 4393 25464
rect 4347 25314 4393 25360
rect 4347 25210 4393 25256
rect 4571 27406 4617 27452
rect 4571 27301 4617 27347
rect 4571 27196 4617 27242
rect 4571 27091 4617 27137
rect 4571 26986 4617 27032
rect 4571 26881 4617 26927
rect 4571 26776 4617 26822
rect 4571 26671 4617 26717
rect 4571 26566 4617 26612
rect 4571 26461 4617 26507
rect 4571 26356 4617 26402
rect 4571 26251 4617 26297
rect 4571 26146 4617 26192
rect 4571 26042 4617 26088
rect 4571 25938 4617 25984
rect 4571 25834 4617 25880
rect 4571 25730 4617 25776
rect 4571 25626 4617 25672
rect 4571 25522 4617 25568
rect 4571 25418 4617 25464
rect 4571 25314 4617 25360
rect 4571 25210 4617 25256
rect 4795 27406 4841 27452
rect 4795 27301 4841 27347
rect 4795 27196 4841 27242
rect 4795 27091 4841 27137
rect 4795 26986 4841 27032
rect 4795 26881 4841 26927
rect 4795 26776 4841 26822
rect 4795 26671 4841 26717
rect 4795 26566 4841 26612
rect 4795 26461 4841 26507
rect 4795 26356 4841 26402
rect 4795 26251 4841 26297
rect 4795 26146 4841 26192
rect 4795 26042 4841 26088
rect 4795 25938 4841 25984
rect 4795 25834 4841 25880
rect 4795 25730 4841 25776
rect 4795 25626 4841 25672
rect 4795 25522 4841 25568
rect 4795 25418 4841 25464
rect 4795 25314 4841 25360
rect 4795 25210 4841 25256
rect 5019 27406 5065 27452
rect 5019 27301 5065 27347
rect 5019 27196 5065 27242
rect 5019 27091 5065 27137
rect 5019 26986 5065 27032
rect 5019 26881 5065 26927
rect 5019 26776 5065 26822
rect 5019 26671 5065 26717
rect 5019 26566 5065 26612
rect 5019 26461 5065 26507
rect 5019 26356 5065 26402
rect 5019 26251 5065 26297
rect 5019 26146 5065 26192
rect 5019 26042 5065 26088
rect 5019 25938 5065 25984
rect 5019 25834 5065 25880
rect 5019 25730 5065 25776
rect 5019 25626 5065 25672
rect 5019 25522 5065 25568
rect 5019 25418 5065 25464
rect 5019 25314 5065 25360
rect 5019 25210 5065 25256
rect 5243 27406 5289 27452
rect 5243 27301 5289 27347
rect 5243 27196 5289 27242
rect 5243 27091 5289 27137
rect 5933 27336 5979 27382
rect 5933 27132 5979 27178
rect 6381 27336 6427 27382
rect 6381 27132 6427 27178
rect 6829 27336 6875 27382
rect 9038 27406 9084 27452
rect 6829 27132 6875 27178
rect 7409 27269 7455 27315
rect 7409 27113 7455 27159
rect 7633 27269 7679 27315
rect 7633 27113 7679 27159
rect 7857 27269 7903 27315
rect 7857 27113 7903 27159
rect 9038 27301 9084 27347
rect 9038 27196 9084 27242
rect 5243 26986 5289 27032
rect 9038 27091 9084 27137
rect 9038 26986 9084 27032
rect 5243 26881 5289 26927
rect 5243 26776 5289 26822
rect 9038 26881 9084 26927
rect 9038 26776 9084 26822
rect 5243 26671 5289 26717
rect 5243 26566 5289 26612
rect 5243 26461 5289 26507
rect 5243 26356 5289 26402
rect 5243 26251 5289 26297
rect 5243 26146 5289 26192
rect 5243 26042 5289 26088
rect 5243 25938 5289 25984
rect 5243 25834 5289 25880
rect 5243 25730 5289 25776
rect 5243 25626 5289 25672
rect 5243 25522 5289 25568
rect 5243 25418 5289 25464
rect 5243 25314 5289 25360
rect 9038 26671 9084 26717
rect 9038 26566 9084 26612
rect 9038 26461 9084 26507
rect 9038 26356 9084 26402
rect 9038 26251 9084 26297
rect 9038 26146 9084 26192
rect 9038 26042 9084 26088
rect 9038 25938 9084 25984
rect 9038 25834 9084 25880
rect 9038 25730 9084 25776
rect 9038 25626 9084 25672
rect 9038 25522 9084 25568
rect 9038 25418 9084 25464
rect 5243 25210 5289 25256
rect 9038 25314 9084 25360
rect 9038 25210 9084 25256
rect 9262 27406 9308 27452
rect 9262 27301 9308 27347
rect 9262 27196 9308 27242
rect 9262 27091 9308 27137
rect 9262 26986 9308 27032
rect 9262 26881 9308 26927
rect 9262 26776 9308 26822
rect 9262 26671 9308 26717
rect 9262 26566 9308 26612
rect 9262 26461 9308 26507
rect 9262 26356 9308 26402
rect 9262 26251 9308 26297
rect 9262 26146 9308 26192
rect 9262 26042 9308 26088
rect 9262 25938 9308 25984
rect 9262 25834 9308 25880
rect 9262 25730 9308 25776
rect 9262 25626 9308 25672
rect 9262 25522 9308 25568
rect 9262 25418 9308 25464
rect 9262 25314 9308 25360
rect 9262 25210 9308 25256
rect 9486 27406 9532 27452
rect 9486 27301 9532 27347
rect 9486 27196 9532 27242
rect 9486 27091 9532 27137
rect 9486 26986 9532 27032
rect 9486 26881 9532 26927
rect 9486 26776 9532 26822
rect 9486 26671 9532 26717
rect 9486 26566 9532 26612
rect 9486 26461 9532 26507
rect 9486 26356 9532 26402
rect 9486 26251 9532 26297
rect 9486 26146 9532 26192
rect 9486 26042 9532 26088
rect 9486 25938 9532 25984
rect 9486 25834 9532 25880
rect 9486 25730 9532 25776
rect 9486 25626 9532 25672
rect 9486 25522 9532 25568
rect 9486 25418 9532 25464
rect 9486 25314 9532 25360
rect 9486 25210 9532 25256
rect 9710 27406 9756 27452
rect 9710 27301 9756 27347
rect 9710 27196 9756 27242
rect 9710 27091 9756 27137
rect 9710 26986 9756 27032
rect 9710 26881 9756 26927
rect 9710 26776 9756 26822
rect 9710 26671 9756 26717
rect 9710 26566 9756 26612
rect 9710 26461 9756 26507
rect 9710 26356 9756 26402
rect 9710 26251 9756 26297
rect 9710 26146 9756 26192
rect 9710 26042 9756 26088
rect 9710 25938 9756 25984
rect 9710 25834 9756 25880
rect 9710 25730 9756 25776
rect 9710 25626 9756 25672
rect 9710 25522 9756 25568
rect 9710 25418 9756 25464
rect 9710 25314 9756 25360
rect 9710 25210 9756 25256
rect 9934 27406 9980 27452
rect 9934 27301 9980 27347
rect 9934 27196 9980 27242
rect 9934 27091 9980 27137
rect 9934 26986 9980 27032
rect 9934 26881 9980 26927
rect 9934 26776 9980 26822
rect 9934 26671 9980 26717
rect 9934 26566 9980 26612
rect 9934 26461 9980 26507
rect 9934 26356 9980 26402
rect 9934 26251 9980 26297
rect 9934 26146 9980 26192
rect 9934 26042 9980 26088
rect 9934 25938 9980 25984
rect 9934 25834 9980 25880
rect 9934 25730 9980 25776
rect 9934 25626 9980 25672
rect 9934 25522 9980 25568
rect 9934 25418 9980 25464
rect 9934 25314 9980 25360
rect 9934 25210 9980 25256
rect 10158 27406 10204 27452
rect 10158 27301 10204 27347
rect 10158 27196 10204 27242
rect 10158 27091 10204 27137
rect 10158 26986 10204 27032
rect 10158 26881 10204 26927
rect 10158 26776 10204 26822
rect 10158 26671 10204 26717
rect 10158 26566 10204 26612
rect 10158 26461 10204 26507
rect 10158 26356 10204 26402
rect 10158 26251 10204 26297
rect 10158 26146 10204 26192
rect 10158 26042 10204 26088
rect 10158 25938 10204 25984
rect 10158 25834 10204 25880
rect 10158 25730 10204 25776
rect 10158 25626 10204 25672
rect 10158 25522 10204 25568
rect 10158 25418 10204 25464
rect 10158 25314 10204 25360
rect 10158 25210 10204 25256
rect 10382 27406 10428 27452
rect 10382 27301 10428 27347
rect 10382 27196 10428 27242
rect 10382 27091 10428 27137
rect 10382 26986 10428 27032
rect 10382 26881 10428 26927
rect 10382 26776 10428 26822
rect 10382 26671 10428 26717
rect 10382 26566 10428 26612
rect 10382 26461 10428 26507
rect 10382 26356 10428 26402
rect 10382 26251 10428 26297
rect 10382 26146 10428 26192
rect 10382 26042 10428 26088
rect 10382 25938 10428 25984
rect 10382 25834 10428 25880
rect 10382 25730 10428 25776
rect 10382 25626 10428 25672
rect 10382 25522 10428 25568
rect 10382 25418 10428 25464
rect 10382 25314 10428 25360
rect 10382 25210 10428 25256
rect 10606 27406 10652 27452
rect 10606 27301 10652 27347
rect 10606 27196 10652 27242
rect 10606 27091 10652 27137
rect 10606 26986 10652 27032
rect 10606 26881 10652 26927
rect 10606 26776 10652 26822
rect 10606 26671 10652 26717
rect 10606 26566 10652 26612
rect 10606 26461 10652 26507
rect 10606 26356 10652 26402
rect 10606 26251 10652 26297
rect 10606 26146 10652 26192
rect 10606 26042 10652 26088
rect 10606 25938 10652 25984
rect 10606 25834 10652 25880
rect 10606 25730 10652 25776
rect 10606 25626 10652 25672
rect 10606 25522 10652 25568
rect 10606 25418 10652 25464
rect 10606 25314 10652 25360
rect 10606 25210 10652 25256
rect 10830 27406 10876 27452
rect 10830 27301 10876 27347
rect 10830 27196 10876 27242
rect 10830 27091 10876 27137
rect 10830 26986 10876 27032
rect 10830 26881 10876 26927
rect 10830 26776 10876 26822
rect 10830 26671 10876 26717
rect 10830 26566 10876 26612
rect 10830 26461 10876 26507
rect 10830 26356 10876 26402
rect 10830 26251 10876 26297
rect 10830 26146 10876 26192
rect 10830 26042 10876 26088
rect 10830 25938 10876 25984
rect 10830 25834 10876 25880
rect 10830 25730 10876 25776
rect 10830 25626 10876 25672
rect 10830 25522 10876 25568
rect 10830 25418 10876 25464
rect 10830 25314 10876 25360
rect 10830 25210 10876 25256
rect 11054 27406 11100 27452
rect 11054 27301 11100 27347
rect 11054 27196 11100 27242
rect 11054 27091 11100 27137
rect 11054 26986 11100 27032
rect 11054 26881 11100 26927
rect 11054 26776 11100 26822
rect 11054 26671 11100 26717
rect 11054 26566 11100 26612
rect 11054 26461 11100 26507
rect 11054 26356 11100 26402
rect 11054 26251 11100 26297
rect 11054 26146 11100 26192
rect 11054 26042 11100 26088
rect 11054 25938 11100 25984
rect 11054 25834 11100 25880
rect 11054 25730 11100 25776
rect 11054 25626 11100 25672
rect 11054 25522 11100 25568
rect 11054 25418 11100 25464
rect 11054 25314 11100 25360
rect 11054 25210 11100 25256
rect 11278 27406 11324 27452
rect 11278 27301 11324 27347
rect 11278 27196 11324 27242
rect 11278 27091 11324 27137
rect 11278 26986 11324 27032
rect 11278 26881 11324 26927
rect 11278 26776 11324 26822
rect 11278 26671 11324 26717
rect 11278 26566 11324 26612
rect 11278 26461 11324 26507
rect 11278 26356 11324 26402
rect 11278 26251 11324 26297
rect 11278 26146 11324 26192
rect 11278 26042 11324 26088
rect 11278 25938 11324 25984
rect 11278 25834 11324 25880
rect 11278 25730 11324 25776
rect 11278 25626 11324 25672
rect 11278 25522 11324 25568
rect 11278 25418 11324 25464
rect 11278 25314 11324 25360
rect 11278 25210 11324 25256
rect 11502 27406 11548 27452
rect 11502 27301 11548 27347
rect 11502 27196 11548 27242
rect 11502 27091 11548 27137
rect 11502 26986 11548 27032
rect 11502 26881 11548 26927
rect 11502 26776 11548 26822
rect 11502 26671 11548 26717
rect 11502 26566 11548 26612
rect 11502 26461 11548 26507
rect 11502 26356 11548 26402
rect 11502 26251 11548 26297
rect 11502 26146 11548 26192
rect 11502 26042 11548 26088
rect 11502 25938 11548 25984
rect 11502 25834 11548 25880
rect 11502 25730 11548 25776
rect 11502 25626 11548 25672
rect 11502 25522 11548 25568
rect 11502 25418 11548 25464
rect 11502 25314 11548 25360
rect 11502 25210 11548 25256
rect 11726 27406 11772 27452
rect 11726 27301 11772 27347
rect 11726 27196 11772 27242
rect 11726 27091 11772 27137
rect 11726 26986 11772 27032
rect 11726 26881 11772 26927
rect 11726 26776 11772 26822
rect 11726 26671 11772 26717
rect 11726 26566 11772 26612
rect 11726 26461 11772 26507
rect 11726 26356 11772 26402
rect 11726 26251 11772 26297
rect 11726 26146 11772 26192
rect 11726 26042 11772 26088
rect 11726 25938 11772 25984
rect 11726 25834 11772 25880
rect 11726 25730 11772 25776
rect 11726 25626 11772 25672
rect 11726 25522 11772 25568
rect 11726 25418 11772 25464
rect 11726 25314 11772 25360
rect 11726 25210 11772 25256
rect 11950 27406 11996 27452
rect 11950 27301 11996 27347
rect 11950 27196 11996 27242
rect 11950 27091 11996 27137
rect 11950 26986 11996 27032
rect 11950 26881 11996 26927
rect 11950 26776 11996 26822
rect 11950 26671 11996 26717
rect 11950 26566 11996 26612
rect 11950 26461 11996 26507
rect 11950 26356 11996 26402
rect 11950 26251 11996 26297
rect 11950 26146 11996 26192
rect 11950 26042 11996 26088
rect 11950 25938 11996 25984
rect 11950 25834 11996 25880
rect 11950 25730 11996 25776
rect 11950 25626 11996 25672
rect 11950 25522 11996 25568
rect 11950 25418 11996 25464
rect 11950 25314 11996 25360
rect 11950 25210 11996 25256
rect 12174 27406 12220 27452
rect 12174 27301 12220 27347
rect 12174 27196 12220 27242
rect 12174 27091 12220 27137
rect 12174 26986 12220 27032
rect 12174 26881 12220 26927
rect 12174 26776 12220 26822
rect 12174 26671 12220 26717
rect 12174 26566 12220 26612
rect 12174 26461 12220 26507
rect 12174 26356 12220 26402
rect 12174 26251 12220 26297
rect 12174 26146 12220 26192
rect 12174 26042 12220 26088
rect 12174 25938 12220 25984
rect 12174 25834 12220 25880
rect 12174 25730 12220 25776
rect 12174 25626 12220 25672
rect 12174 25522 12220 25568
rect 12174 25418 12220 25464
rect 12174 25314 12220 25360
rect 12174 25210 12220 25256
rect 12398 27406 12444 27452
rect 12398 27301 12444 27347
rect 12398 27196 12444 27242
rect 12398 27091 12444 27137
rect 12398 26986 12444 27032
rect 12398 26881 12444 26927
rect 12398 26776 12444 26822
rect 12398 26671 12444 26717
rect 12398 26566 12444 26612
rect 12398 26461 12444 26507
rect 12398 26356 12444 26402
rect 12398 26251 12444 26297
rect 12398 26146 12444 26192
rect 12398 26042 12444 26088
rect 12398 25938 12444 25984
rect 12398 25834 12444 25880
rect 12398 25730 12444 25776
rect 12398 25626 12444 25672
rect 12398 25522 12444 25568
rect 12398 25418 12444 25464
rect 12398 25314 12444 25360
rect 12398 25210 12444 25256
rect 12622 27406 12668 27452
rect 12622 27301 12668 27347
rect 12622 27196 12668 27242
rect 12622 27091 12668 27137
rect 13312 27336 13358 27382
rect 13312 27132 13358 27178
rect 13760 27336 13806 27382
rect 13760 27132 13806 27178
rect 14208 27336 14254 27382
rect 14208 27132 14254 27178
rect 14788 27269 14834 27315
rect 14788 27113 14834 27159
rect 15012 27269 15058 27315
rect 15012 27113 15058 27159
rect 15236 27269 15282 27315
rect 15236 27113 15282 27159
rect 23797 27336 23843 27382
rect 12622 26986 12668 27032
rect 12622 26881 12668 26927
rect 23797 27132 23843 27178
rect 24245 27336 24291 27382
rect 24245 27132 24291 27178
rect 24693 27336 24739 27382
rect 25273 27383 25319 27429
rect 25273 27248 25319 27294
rect 24693 27132 24739 27178
rect 25273 27113 25319 27159
rect 25497 27383 25543 27429
rect 25497 27248 25543 27294
rect 25497 27113 25543 27159
rect 25721 27383 25767 27429
rect 25721 27248 25767 27294
rect 25721 27113 25767 27159
rect 12622 26776 12668 26822
rect 16704 26842 16750 26888
rect 12622 26671 12668 26717
rect 12622 26566 12668 26612
rect 12622 26461 12668 26507
rect 12622 26356 12668 26402
rect 12622 26251 12668 26297
rect 12622 26146 12668 26192
rect 12622 26042 12668 26088
rect 12622 25938 12668 25984
rect 12622 25834 12668 25880
rect 12622 25730 12668 25776
rect 12622 25626 12668 25672
rect 12622 25522 12668 25568
rect 12622 25418 12668 25464
rect 12622 25314 12668 25360
rect 16704 26737 16750 26783
rect 16704 26632 16750 26678
rect 16704 26527 16750 26573
rect 16704 26422 16750 26468
rect 16704 26317 16750 26363
rect 16704 26212 16750 26258
rect 16704 26107 16750 26153
rect 16704 26002 16750 26048
rect 16704 25897 16750 25943
rect 16704 25792 16750 25838
rect 16704 25687 16750 25733
rect 16704 25582 16750 25628
rect 16704 25478 16750 25524
rect 12622 25210 12668 25256
rect 1817 22566 1863 24550
rect 1817 22463 1863 22509
rect 1817 22360 1863 22406
rect 1817 22257 1863 22303
rect 1817 22154 1863 22200
rect 1817 22051 1863 22097
rect 1817 21948 1863 21994
rect 1817 21845 1863 21891
rect 1817 21742 1863 21788
rect 1817 21639 1863 21685
rect 1817 21536 1863 21582
rect 2041 22566 2087 24550
rect 2041 22463 2087 22509
rect 2041 22360 2087 22406
rect 2041 22257 2087 22303
rect 2041 22154 2087 22200
rect 2041 22051 2087 22097
rect 2041 21948 2087 21994
rect 2041 21845 2087 21891
rect 2041 21742 2087 21788
rect 2041 21639 2087 21685
rect 2041 21536 2087 21582
rect 2265 22566 2311 24550
rect 2265 22463 2311 22509
rect 2265 22360 2311 22406
rect 2265 22257 2311 22303
rect 2265 22154 2311 22200
rect 2265 22051 2311 22097
rect 2845 22566 2891 24550
rect 2845 22463 2891 22509
rect 2845 22360 2891 22406
rect 2845 22257 2891 22303
rect 2845 22154 2891 22200
rect 2845 22051 2891 22097
rect 2265 21948 2311 21994
rect 2265 21845 2311 21891
rect 2265 21742 2311 21788
rect 2265 21639 2311 21685
rect 2845 21948 2891 21994
rect 2845 21845 2891 21891
rect 2845 21742 2891 21788
rect 2265 21536 2311 21582
rect 2845 21639 2891 21685
rect 2845 21536 2891 21582
rect 3069 22566 3115 24550
rect 3069 22463 3115 22509
rect 3069 22360 3115 22406
rect 3069 22257 3115 22303
rect 3069 22154 3115 22200
rect 3069 22051 3115 22097
rect 3069 21948 3115 21994
rect 3069 21845 3115 21891
rect 3069 21742 3115 21788
rect 3069 21639 3115 21685
rect 3069 21536 3115 21582
rect 3293 22566 3339 24550
rect 3293 22463 3339 22509
rect 3293 22360 3339 22406
rect 3293 22257 3339 22303
rect 3293 22154 3339 22200
rect 3293 22051 3339 22097
rect 3293 21948 3339 21994
rect 3293 21845 3339 21891
rect 3293 21742 3339 21788
rect 3293 21639 3339 21685
rect 3293 21536 3339 21582
rect 3609 22566 3655 24550
rect 3609 22463 3655 22509
rect 3609 22360 3655 22406
rect 3609 22257 3655 22303
rect 3609 22154 3655 22200
rect 3609 22051 3655 22097
rect 3609 21948 3655 21994
rect 3609 21845 3655 21891
rect 3609 21742 3655 21788
rect 3609 21639 3655 21685
rect 3609 21536 3655 21582
rect 3833 22566 3879 24550
rect 3833 22463 3879 22509
rect 3833 22360 3879 22406
rect 3833 22257 3879 22303
rect 3833 22154 3879 22200
rect 3833 22051 3879 22097
rect 3833 21948 3879 21994
rect 3833 21845 3879 21891
rect 3833 21742 3879 21788
rect 3833 21639 3879 21685
rect 3833 21536 3879 21582
rect 4057 22566 4103 24550
rect 4057 22463 4103 22509
rect 4057 22360 4103 22406
rect 4057 22257 4103 22303
rect 4057 22154 4103 22200
rect 4057 22051 4103 22097
rect 4637 22566 4683 24550
rect 4637 22463 4683 22509
rect 4637 22360 4683 22406
rect 4637 22257 4683 22303
rect 4637 22154 4683 22200
rect 4637 22051 4683 22097
rect 4057 21948 4103 21994
rect 4057 21845 4103 21891
rect 4057 21742 4103 21788
rect 4057 21639 4103 21685
rect 4637 21948 4683 21994
rect 4637 21845 4683 21891
rect 4637 21742 4683 21788
rect 4057 21536 4103 21582
rect 4637 21639 4683 21685
rect 4637 21536 4683 21582
rect 4861 22566 4907 24550
rect 4861 22463 4907 22509
rect 4861 22360 4907 22406
rect 4861 22257 4907 22303
rect 4861 22154 4907 22200
rect 4861 22051 4907 22097
rect 4861 21948 4907 21994
rect 4861 21845 4907 21891
rect 4861 21742 4907 21788
rect 4861 21639 4907 21685
rect 4861 21536 4907 21582
rect 5085 22566 5131 24550
rect 5085 22463 5131 22509
rect 5085 22360 5131 22406
rect 5085 22257 5131 22303
rect 5085 22154 5131 22200
rect 5085 22051 5131 22097
rect 5085 21948 5131 21994
rect 5085 21845 5131 21891
rect 5085 21742 5131 21788
rect 5085 21639 5131 21685
rect 5085 21536 5131 21582
rect 6091 21490 6137 25002
rect 6315 21490 6361 25002
rect 6605 23427 6651 25003
rect 6605 23324 6651 23370
rect 6605 23221 6651 23267
rect 6605 23118 6651 23164
rect 6605 23015 6651 23061
rect 6605 22912 6651 22958
rect 6605 22809 6651 22855
rect 6605 22706 6651 22752
rect 6605 22603 6651 22649
rect 6605 22500 6651 22546
rect 6605 22397 6651 22443
rect 6829 23427 6875 25003
rect 6829 23324 6875 23370
rect 6829 23221 6875 23267
rect 6829 23118 6875 23164
rect 6829 23015 6875 23061
rect 6829 22912 6875 22958
rect 6829 22809 6875 22855
rect 6829 22706 6875 22752
rect 6829 22603 6875 22649
rect 6829 22500 6875 22546
rect 6829 22397 6875 22443
rect 7782 21490 7828 25002
rect 8006 21490 8052 25002
rect 8296 23427 8342 25003
rect 8296 23324 8342 23370
rect 8296 23221 8342 23267
rect 8296 23118 8342 23164
rect 8296 23015 8342 23061
rect 8296 22912 8342 22958
rect 8296 22809 8342 22855
rect 8296 22706 8342 22752
rect 8296 22603 8342 22649
rect 8296 22500 8342 22546
rect 8296 22397 8342 22443
rect 8520 23427 8566 25003
rect 8520 23324 8566 23370
rect 8520 23221 8566 23267
rect 8520 23118 8566 23164
rect 8520 23015 8566 23061
rect 8520 22912 8566 22958
rect 8520 22809 8566 22855
rect 8520 22706 8566 22752
rect 8520 22603 8566 22649
rect 8520 22500 8566 22546
rect 8520 22397 8566 22443
rect 9196 22566 9242 24550
rect 9196 22463 9242 22509
rect 9196 22360 9242 22406
rect 9196 22257 9242 22303
rect 9196 22154 9242 22200
rect 9196 22051 9242 22097
rect 9196 21948 9242 21994
rect 9196 21845 9242 21891
rect 9196 21742 9242 21788
rect 9196 21639 9242 21685
rect 9196 21536 9242 21582
rect 9420 22566 9466 24550
rect 9420 22463 9466 22509
rect 9420 22360 9466 22406
rect 9420 22257 9466 22303
rect 9420 22154 9466 22200
rect 9420 22051 9466 22097
rect 9420 21948 9466 21994
rect 9420 21845 9466 21891
rect 9420 21742 9466 21788
rect 9420 21639 9466 21685
rect 9420 21536 9466 21582
rect 9644 22566 9690 24550
rect 9644 22463 9690 22509
rect 9644 22360 9690 22406
rect 9644 22257 9690 22303
rect 9644 22154 9690 22200
rect 9644 22051 9690 22097
rect 10224 22566 10270 24550
rect 10224 22463 10270 22509
rect 10224 22360 10270 22406
rect 10224 22257 10270 22303
rect 10224 22154 10270 22200
rect 10224 22051 10270 22097
rect 9644 21948 9690 21994
rect 9644 21845 9690 21891
rect 9644 21742 9690 21788
rect 9644 21639 9690 21685
rect 10224 21948 10270 21994
rect 10224 21845 10270 21891
rect 10224 21742 10270 21788
rect 9644 21536 9690 21582
rect 10224 21639 10270 21685
rect 10224 21536 10270 21582
rect 10448 22566 10494 24550
rect 10448 22463 10494 22509
rect 10448 22360 10494 22406
rect 10448 22257 10494 22303
rect 10448 22154 10494 22200
rect 10448 22051 10494 22097
rect 10448 21948 10494 21994
rect 10448 21845 10494 21891
rect 10448 21742 10494 21788
rect 10448 21639 10494 21685
rect 10448 21536 10494 21582
rect 10672 22566 10718 24550
rect 10672 22463 10718 22509
rect 10672 22360 10718 22406
rect 10672 22257 10718 22303
rect 10672 22154 10718 22200
rect 10672 22051 10718 22097
rect 10672 21948 10718 21994
rect 10672 21845 10718 21891
rect 10672 21742 10718 21788
rect 10672 21639 10718 21685
rect 10672 21536 10718 21582
rect 10988 22566 11034 24550
rect 10988 22463 11034 22509
rect 10988 22360 11034 22406
rect 10988 22257 11034 22303
rect 10988 22154 11034 22200
rect 10988 22051 11034 22097
rect 10988 21948 11034 21994
rect 10988 21845 11034 21891
rect 10988 21742 11034 21788
rect 10988 21639 11034 21685
rect 10988 21536 11034 21582
rect 11212 22566 11258 24550
rect 11212 22463 11258 22509
rect 11212 22360 11258 22406
rect 11212 22257 11258 22303
rect 11212 22154 11258 22200
rect 11212 22051 11258 22097
rect 11212 21948 11258 21994
rect 11212 21845 11258 21891
rect 11212 21742 11258 21788
rect 11212 21639 11258 21685
rect 11212 21536 11258 21582
rect 11436 22566 11482 24550
rect 11436 22463 11482 22509
rect 11436 22360 11482 22406
rect 11436 22257 11482 22303
rect 11436 22154 11482 22200
rect 11436 22051 11482 22097
rect 12016 22566 12062 24550
rect 12016 22463 12062 22509
rect 12016 22360 12062 22406
rect 12016 22257 12062 22303
rect 12016 22154 12062 22200
rect 12016 22051 12062 22097
rect 11436 21948 11482 21994
rect 11436 21845 11482 21891
rect 11436 21742 11482 21788
rect 11436 21639 11482 21685
rect 12016 21948 12062 21994
rect 12016 21845 12062 21891
rect 12016 21742 12062 21788
rect 11436 21536 11482 21582
rect 12016 21639 12062 21685
rect 12016 21536 12062 21582
rect 12240 22566 12286 24550
rect 12240 22463 12286 22509
rect 12240 22360 12286 22406
rect 12240 22257 12286 22303
rect 12240 22154 12286 22200
rect 12240 22051 12286 22097
rect 12240 21948 12286 21994
rect 12240 21845 12286 21891
rect 12240 21742 12286 21788
rect 12240 21639 12286 21685
rect 12240 21536 12286 21582
rect 12464 22566 12510 24550
rect 12464 22463 12510 22509
rect 12464 22360 12510 22406
rect 12464 22257 12510 22303
rect 12464 22154 12510 22200
rect 12464 22051 12510 22097
rect 12464 21948 12510 21994
rect 12464 21845 12510 21891
rect 12464 21742 12510 21788
rect 12464 21639 12510 21685
rect 12464 21536 12510 21582
rect 13470 21490 13516 25002
rect 13694 21490 13740 25002
rect 13984 23427 14030 25003
rect 13984 23324 14030 23370
rect 13984 23221 14030 23267
rect 13984 23118 14030 23164
rect 13984 23015 14030 23061
rect 13984 22912 14030 22958
rect 13984 22809 14030 22855
rect 13984 22706 14030 22752
rect 13984 22603 14030 22649
rect 13984 22500 14030 22546
rect 13984 22397 14030 22443
rect 16704 25374 16750 25420
rect 16704 25270 16750 25316
rect 16704 25166 16750 25212
rect 16704 25062 16750 25108
rect 14208 23427 14254 25003
rect 14208 23324 14254 23370
rect 14208 23221 14254 23267
rect 14208 23118 14254 23164
rect 14208 23015 14254 23061
rect 14208 22912 14254 22958
rect 14208 22809 14254 22855
rect 14208 22706 14254 22752
rect 14208 22603 14254 22649
rect 14208 22500 14254 22546
rect 14208 22397 14254 22443
rect 15161 21490 15207 25002
rect 15385 21490 15431 25002
rect 15675 23427 15721 25003
rect 15675 23324 15721 23370
rect 15675 23221 15721 23267
rect 15675 23118 15721 23164
rect 15675 23015 15721 23061
rect 15675 22912 15721 22958
rect 15675 22809 15721 22855
rect 15675 22706 15721 22752
rect 15675 22603 15721 22649
rect 15675 22500 15721 22546
rect 15675 22397 15721 22443
rect 15899 23427 15945 25003
rect 16704 24958 16750 25004
rect 16704 24854 16750 24900
rect 16704 24750 16750 24796
rect 16704 24646 16750 24692
rect 16928 26842 16974 26888
rect 16928 26737 16974 26783
rect 16928 26632 16974 26678
rect 16928 26527 16974 26573
rect 16928 26422 16974 26468
rect 16928 26317 16974 26363
rect 16928 26212 16974 26258
rect 16928 26107 16974 26153
rect 16928 26002 16974 26048
rect 16928 25897 16974 25943
rect 16928 25792 16974 25838
rect 16928 25687 16974 25733
rect 16928 25582 16974 25628
rect 16928 25478 16974 25524
rect 16928 25374 16974 25420
rect 16928 25270 16974 25316
rect 16928 25166 16974 25212
rect 16928 25062 16974 25108
rect 16928 24958 16974 25004
rect 16928 24854 16974 24900
rect 16928 24750 16974 24796
rect 16928 24646 16974 24692
rect 17152 26842 17198 26888
rect 17152 26737 17198 26783
rect 17152 26632 17198 26678
rect 17152 26527 17198 26573
rect 17152 26422 17198 26468
rect 17152 26317 17198 26363
rect 17152 26212 17198 26258
rect 17152 26107 17198 26153
rect 17152 26002 17198 26048
rect 17152 25897 17198 25943
rect 17152 25792 17198 25838
rect 17152 25687 17198 25733
rect 17152 25582 17198 25628
rect 17152 25478 17198 25524
rect 17152 25374 17198 25420
rect 17152 25270 17198 25316
rect 17152 25166 17198 25212
rect 17152 25062 17198 25108
rect 17152 24958 17198 25004
rect 17152 24854 17198 24900
rect 17152 24750 17198 24796
rect 17152 24646 17198 24692
rect 17376 26842 17422 26888
rect 17376 26737 17422 26783
rect 17376 26632 17422 26678
rect 17376 26527 17422 26573
rect 17376 26422 17422 26468
rect 17376 26317 17422 26363
rect 17376 26212 17422 26258
rect 17376 26107 17422 26153
rect 17376 26002 17422 26048
rect 17376 25897 17422 25943
rect 17376 25792 17422 25838
rect 17376 25687 17422 25733
rect 17376 25582 17422 25628
rect 17376 25478 17422 25524
rect 17376 25374 17422 25420
rect 17376 25270 17422 25316
rect 17376 25166 17422 25212
rect 17376 25062 17422 25108
rect 17376 24958 17422 25004
rect 17376 24854 17422 24900
rect 17376 24750 17422 24796
rect 17376 24646 17422 24692
rect 17600 26842 17646 26888
rect 17600 26737 17646 26783
rect 17600 26632 17646 26678
rect 17600 26527 17646 26573
rect 17600 26422 17646 26468
rect 17600 26317 17646 26363
rect 17600 26212 17646 26258
rect 17600 26107 17646 26153
rect 17600 26002 17646 26048
rect 17600 25897 17646 25943
rect 17600 25792 17646 25838
rect 17600 25687 17646 25733
rect 17600 25582 17646 25628
rect 17600 25478 17646 25524
rect 17600 25374 17646 25420
rect 17600 25270 17646 25316
rect 17600 25166 17646 25212
rect 17600 25062 17646 25108
rect 17600 24958 17646 25004
rect 17600 24854 17646 24900
rect 17600 24750 17646 24796
rect 17600 24646 17646 24692
rect 17824 26842 17870 26888
rect 17824 26737 17870 26783
rect 17824 26632 17870 26678
rect 17824 26527 17870 26573
rect 17824 26422 17870 26468
rect 17824 26317 17870 26363
rect 17824 26212 17870 26258
rect 17824 26107 17870 26153
rect 17824 26002 17870 26048
rect 17824 25897 17870 25943
rect 17824 25792 17870 25838
rect 17824 25687 17870 25733
rect 17824 25582 17870 25628
rect 17824 25478 17870 25524
rect 17824 25374 17870 25420
rect 17824 25270 17870 25316
rect 17824 25166 17870 25212
rect 17824 25062 17870 25108
rect 17824 24958 17870 25004
rect 17824 24854 17870 24900
rect 17824 24750 17870 24796
rect 17824 24646 17870 24692
rect 18048 26842 18094 26888
rect 18048 26737 18094 26783
rect 18048 26632 18094 26678
rect 18048 26527 18094 26573
rect 18048 26422 18094 26468
rect 18048 26317 18094 26363
rect 18048 26212 18094 26258
rect 18048 26107 18094 26153
rect 18048 26002 18094 26048
rect 18048 25897 18094 25943
rect 18048 25792 18094 25838
rect 18048 25687 18094 25733
rect 18048 25582 18094 25628
rect 18048 25478 18094 25524
rect 18048 25374 18094 25420
rect 18048 25270 18094 25316
rect 18048 25166 18094 25212
rect 18048 25062 18094 25108
rect 18048 24958 18094 25004
rect 18048 24854 18094 24900
rect 18048 24750 18094 24796
rect 18048 24646 18094 24692
rect 18338 26842 18384 26888
rect 18338 26737 18384 26783
rect 18338 26632 18384 26678
rect 18338 26527 18384 26573
rect 18338 26422 18384 26468
rect 18338 26317 18384 26363
rect 18338 26212 18384 26258
rect 18338 26107 18384 26153
rect 18338 26002 18384 26048
rect 18338 25897 18384 25943
rect 18338 25792 18384 25838
rect 18338 25687 18384 25733
rect 18338 25582 18384 25628
rect 18338 25478 18384 25524
rect 18338 25374 18384 25420
rect 18338 25270 18384 25316
rect 18338 25166 18384 25212
rect 18338 25062 18384 25108
rect 18338 24958 18384 25004
rect 18338 24854 18384 24900
rect 18338 24750 18384 24796
rect 18338 24646 18384 24692
rect 18562 26842 18608 26888
rect 18562 26737 18608 26783
rect 18562 26632 18608 26678
rect 18562 26527 18608 26573
rect 18562 26422 18608 26468
rect 18562 26317 18608 26363
rect 18562 26212 18608 26258
rect 18562 26107 18608 26153
rect 18562 26002 18608 26048
rect 18562 25897 18608 25943
rect 18562 25792 18608 25838
rect 18562 25687 18608 25733
rect 18562 25582 18608 25628
rect 18562 25478 18608 25524
rect 18562 25374 18608 25420
rect 18562 25270 18608 25316
rect 18562 25166 18608 25212
rect 18562 25062 18608 25108
rect 18562 24958 18608 25004
rect 18562 24854 18608 24900
rect 18562 24750 18608 24796
rect 18562 24646 18608 24692
rect 18786 26842 18832 26888
rect 18786 26737 18832 26783
rect 18786 26632 18832 26678
rect 18786 26527 18832 26573
rect 18786 26422 18832 26468
rect 18786 26317 18832 26363
rect 18786 26212 18832 26258
rect 18786 26107 18832 26153
rect 18786 26002 18832 26048
rect 18786 25897 18832 25943
rect 18786 25792 18832 25838
rect 18786 25687 18832 25733
rect 18786 25582 18832 25628
rect 18786 25478 18832 25524
rect 18786 25374 18832 25420
rect 18786 25270 18832 25316
rect 18786 25166 18832 25212
rect 18786 25062 18832 25108
rect 18786 24958 18832 25004
rect 18786 24854 18832 24900
rect 18786 24750 18832 24796
rect 18786 24646 18832 24692
rect 19010 26842 19056 26888
rect 19010 26737 19056 26783
rect 19010 26632 19056 26678
rect 19010 26527 19056 26573
rect 19010 26422 19056 26468
rect 19010 26317 19056 26363
rect 19010 26212 19056 26258
rect 19010 26107 19056 26153
rect 19010 26002 19056 26048
rect 19010 25897 19056 25943
rect 19010 25792 19056 25838
rect 19010 25687 19056 25733
rect 19010 25582 19056 25628
rect 19010 25478 19056 25524
rect 19010 25374 19056 25420
rect 19010 25270 19056 25316
rect 19010 25166 19056 25212
rect 19010 25062 19056 25108
rect 19010 24958 19056 25004
rect 19010 24854 19056 24900
rect 19010 24750 19056 24796
rect 19010 24646 19056 24692
rect 19234 26842 19280 26888
rect 19234 26737 19280 26783
rect 19234 26632 19280 26678
rect 19234 26527 19280 26573
rect 19234 26422 19280 26468
rect 19234 26317 19280 26363
rect 19234 26212 19280 26258
rect 19234 26107 19280 26153
rect 19234 26002 19280 26048
rect 19234 25897 19280 25943
rect 19234 25792 19280 25838
rect 19234 25687 19280 25733
rect 19234 25582 19280 25628
rect 19234 25478 19280 25524
rect 19234 25374 19280 25420
rect 19234 25270 19280 25316
rect 19234 25166 19280 25212
rect 19234 25062 19280 25108
rect 19234 24958 19280 25004
rect 19234 24854 19280 24900
rect 19234 24750 19280 24796
rect 19234 24646 19280 24692
rect 19458 26842 19504 26888
rect 19458 26737 19504 26783
rect 19458 26632 19504 26678
rect 19458 26527 19504 26573
rect 19458 26422 19504 26468
rect 19458 26317 19504 26363
rect 19458 26212 19504 26258
rect 19458 26107 19504 26153
rect 19458 26002 19504 26048
rect 19458 25897 19504 25943
rect 19458 25792 19504 25838
rect 19458 25687 19504 25733
rect 19458 25582 19504 25628
rect 19458 25478 19504 25524
rect 19458 25374 19504 25420
rect 19458 25270 19504 25316
rect 19458 25166 19504 25212
rect 19458 25062 19504 25108
rect 19458 24958 19504 25004
rect 19458 24854 19504 24900
rect 19458 24750 19504 24796
rect 19458 24646 19504 24692
rect 19682 26842 19728 26888
rect 19682 26737 19728 26783
rect 19682 26632 19728 26678
rect 19682 26527 19728 26573
rect 19682 26422 19728 26468
rect 19682 26317 19728 26363
rect 19682 26212 19728 26258
rect 19682 26107 19728 26153
rect 19682 26002 19728 26048
rect 19682 25897 19728 25943
rect 19682 25792 19728 25838
rect 19682 25687 19728 25733
rect 19682 25582 19728 25628
rect 19682 25478 19728 25524
rect 19682 25374 19728 25420
rect 19682 25270 19728 25316
rect 19682 25166 19728 25212
rect 19682 25062 19728 25108
rect 19682 24958 19728 25004
rect 19682 24854 19728 24900
rect 19682 24750 19728 24796
rect 19682 24646 19728 24692
rect 19971 26842 20017 26888
rect 19971 26737 20017 26783
rect 19971 26632 20017 26678
rect 19971 26527 20017 26573
rect 19971 26422 20017 26468
rect 19971 26317 20017 26363
rect 19971 26212 20017 26258
rect 19971 26107 20017 26153
rect 19971 26002 20017 26048
rect 19971 25897 20017 25943
rect 19971 25792 20017 25838
rect 19971 25687 20017 25733
rect 19971 25582 20017 25628
rect 19971 25478 20017 25524
rect 19971 25374 20017 25420
rect 19971 25270 20017 25316
rect 19971 25166 20017 25212
rect 19971 25062 20017 25108
rect 19971 24958 20017 25004
rect 19971 24854 20017 24900
rect 19971 24750 20017 24796
rect 19971 24646 20017 24692
rect 20195 26842 20241 26888
rect 20195 26737 20241 26783
rect 20195 26632 20241 26678
rect 20195 26527 20241 26573
rect 20195 26422 20241 26468
rect 20195 26317 20241 26363
rect 20195 26212 20241 26258
rect 20195 26107 20241 26153
rect 20195 26002 20241 26048
rect 20195 25897 20241 25943
rect 20195 25792 20241 25838
rect 20195 25687 20241 25733
rect 20195 25582 20241 25628
rect 20195 25478 20241 25524
rect 20195 25374 20241 25420
rect 20195 25270 20241 25316
rect 20195 25166 20241 25212
rect 20195 25062 20241 25108
rect 20195 24958 20241 25004
rect 20195 24854 20241 24900
rect 20195 24750 20241 24796
rect 20195 24646 20241 24692
rect 20419 26842 20465 26888
rect 20419 26737 20465 26783
rect 20419 26632 20465 26678
rect 20419 26527 20465 26573
rect 20419 26422 20465 26468
rect 20419 26317 20465 26363
rect 20419 26212 20465 26258
rect 20419 26107 20465 26153
rect 20419 26002 20465 26048
rect 20419 25897 20465 25943
rect 20419 25792 20465 25838
rect 20419 25687 20465 25733
rect 20419 25582 20465 25628
rect 20419 25478 20465 25524
rect 20419 25374 20465 25420
rect 20419 25270 20465 25316
rect 20419 25166 20465 25212
rect 20419 25062 20465 25108
rect 20419 24958 20465 25004
rect 20419 24854 20465 24900
rect 20419 24750 20465 24796
rect 20419 24646 20465 24692
rect 20643 26842 20689 26888
rect 20643 26737 20689 26783
rect 20643 26632 20689 26678
rect 20643 26527 20689 26573
rect 20643 26422 20689 26468
rect 20643 26317 20689 26363
rect 20643 26212 20689 26258
rect 20643 26107 20689 26153
rect 20643 26002 20689 26048
rect 20643 25897 20689 25943
rect 20643 25792 20689 25838
rect 20643 25687 20689 25733
rect 20643 25582 20689 25628
rect 20643 25478 20689 25524
rect 20643 25374 20689 25420
rect 20643 25270 20689 25316
rect 20643 25166 20689 25212
rect 20643 25062 20689 25108
rect 20643 24958 20689 25004
rect 20643 24854 20689 24900
rect 20643 24750 20689 24796
rect 20643 24646 20689 24692
rect 20867 26842 20913 26888
rect 20867 26737 20913 26783
rect 20867 26632 20913 26678
rect 20867 26527 20913 26573
rect 20867 26422 20913 26468
rect 20867 26317 20913 26363
rect 20867 26212 20913 26258
rect 20867 26107 20913 26153
rect 20867 26002 20913 26048
rect 20867 25897 20913 25943
rect 20867 25792 20913 25838
rect 20867 25687 20913 25733
rect 20867 25582 20913 25628
rect 20867 25478 20913 25524
rect 20867 25374 20913 25420
rect 20867 25270 20913 25316
rect 20867 25166 20913 25212
rect 20867 25062 20913 25108
rect 20867 24958 20913 25004
rect 20867 24854 20913 24900
rect 20867 24750 20913 24796
rect 20867 24646 20913 24692
rect 21091 26842 21137 26888
rect 21091 26737 21137 26783
rect 21091 26632 21137 26678
rect 21091 26527 21137 26573
rect 21091 26422 21137 26468
rect 21091 26317 21137 26363
rect 21091 26212 21137 26258
rect 21091 26107 21137 26153
rect 21091 26002 21137 26048
rect 21091 25897 21137 25943
rect 21091 25792 21137 25838
rect 21091 25687 21137 25733
rect 21091 25582 21137 25628
rect 21091 25478 21137 25524
rect 21091 25374 21137 25420
rect 21091 25270 21137 25316
rect 21091 25166 21137 25212
rect 21091 25062 21137 25108
rect 21091 24958 21137 25004
rect 21091 24854 21137 24900
rect 21091 24750 21137 24796
rect 21091 24646 21137 24692
rect 21315 26842 21361 26888
rect 21315 26737 21361 26783
rect 21315 26632 21361 26678
rect 21315 26527 21361 26573
rect 21315 26422 21361 26468
rect 21315 26317 21361 26363
rect 21315 26212 21361 26258
rect 21315 26107 21361 26153
rect 21315 26002 21361 26048
rect 21315 25897 21361 25943
rect 21315 25792 21361 25838
rect 21315 25687 21361 25733
rect 21315 25582 21361 25628
rect 21315 25478 21361 25524
rect 21315 25374 21361 25420
rect 21315 25270 21361 25316
rect 21315 25166 21361 25212
rect 21315 25062 21361 25108
rect 21315 24958 21361 25004
rect 21315 24854 21361 24900
rect 21315 24750 21361 24796
rect 21315 24646 21361 24692
rect 21605 26842 21651 26888
rect 21605 26737 21651 26783
rect 21605 26632 21651 26678
rect 21605 26527 21651 26573
rect 21605 26422 21651 26468
rect 21605 26317 21651 26363
rect 21605 26212 21651 26258
rect 21605 26107 21651 26153
rect 21605 26002 21651 26048
rect 21605 25897 21651 25943
rect 21605 25792 21651 25838
rect 21605 25687 21651 25733
rect 21605 25582 21651 25628
rect 21605 25478 21651 25524
rect 21605 25374 21651 25420
rect 21605 25270 21651 25316
rect 21605 25166 21651 25212
rect 21605 25062 21651 25108
rect 21605 24958 21651 25004
rect 21605 24854 21651 24900
rect 21605 24750 21651 24796
rect 21605 24646 21651 24692
rect 21829 26842 21875 26888
rect 21829 26737 21875 26783
rect 21829 26632 21875 26678
rect 21829 26527 21875 26573
rect 21829 26422 21875 26468
rect 21829 26317 21875 26363
rect 21829 26212 21875 26258
rect 21829 26107 21875 26153
rect 21829 26002 21875 26048
rect 21829 25897 21875 25943
rect 21829 25792 21875 25838
rect 21829 25687 21875 25733
rect 21829 25582 21875 25628
rect 21829 25478 21875 25524
rect 21829 25374 21875 25420
rect 21829 25270 21875 25316
rect 21829 25166 21875 25212
rect 21829 25062 21875 25108
rect 21829 24958 21875 25004
rect 21829 24854 21875 24900
rect 21829 24750 21875 24796
rect 21829 24646 21875 24692
rect 22053 26842 22099 26888
rect 22053 26737 22099 26783
rect 22053 26632 22099 26678
rect 22053 26527 22099 26573
rect 22053 26422 22099 26468
rect 22053 26317 22099 26363
rect 22053 26212 22099 26258
rect 22053 26107 22099 26153
rect 22053 26002 22099 26048
rect 22053 25897 22099 25943
rect 22053 25792 22099 25838
rect 22053 25687 22099 25733
rect 22053 25582 22099 25628
rect 22053 25478 22099 25524
rect 22053 25374 22099 25420
rect 22053 25270 22099 25316
rect 22053 25166 22099 25212
rect 22053 25062 22099 25108
rect 22053 24958 22099 25004
rect 22053 24854 22099 24900
rect 22053 24750 22099 24796
rect 22053 24646 22099 24692
rect 22277 26842 22323 26888
rect 22277 26737 22323 26783
rect 22277 26632 22323 26678
rect 22277 26527 22323 26573
rect 22277 26422 22323 26468
rect 22277 26317 22323 26363
rect 22277 26212 22323 26258
rect 22277 26107 22323 26153
rect 22277 26002 22323 26048
rect 22277 25897 22323 25943
rect 22277 25792 22323 25838
rect 22277 25687 22323 25733
rect 22277 25582 22323 25628
rect 22277 25478 22323 25524
rect 22277 25374 22323 25420
rect 22277 25270 22323 25316
rect 22277 25166 22323 25212
rect 22277 25062 22323 25108
rect 22277 24958 22323 25004
rect 22277 24854 22323 24900
rect 22277 24750 22323 24796
rect 22277 24646 22323 24692
rect 22501 26842 22547 26888
rect 22501 26737 22547 26783
rect 22501 26632 22547 26678
rect 22501 26527 22547 26573
rect 22501 26422 22547 26468
rect 22501 26317 22547 26363
rect 22501 26212 22547 26258
rect 22501 26107 22547 26153
rect 22501 26002 22547 26048
rect 22501 25897 22547 25943
rect 22501 25792 22547 25838
rect 22501 25687 22547 25733
rect 22501 25582 22547 25628
rect 22501 25478 22547 25524
rect 22501 25374 22547 25420
rect 22501 25270 22547 25316
rect 22501 25166 22547 25212
rect 22501 25062 22547 25108
rect 22501 24958 22547 25004
rect 22501 24854 22547 24900
rect 22501 24750 22547 24796
rect 22501 24646 22547 24692
rect 22725 26842 22771 26888
rect 22725 26737 22771 26783
rect 22725 26632 22771 26678
rect 22725 26527 22771 26573
rect 22725 26422 22771 26468
rect 22725 26317 22771 26363
rect 22725 26212 22771 26258
rect 22725 26107 22771 26153
rect 22725 26002 22771 26048
rect 22725 25897 22771 25943
rect 22725 25792 22771 25838
rect 22725 25687 22771 25733
rect 22725 25582 22771 25628
rect 22725 25478 22771 25524
rect 22725 25374 22771 25420
rect 22725 25270 22771 25316
rect 22725 25166 22771 25212
rect 22725 25062 22771 25108
rect 22725 24958 22771 25004
rect 22725 24854 22771 24900
rect 22725 24750 22771 24796
rect 22725 24646 22771 24692
rect 22949 26842 22995 26888
rect 22949 26737 22995 26783
rect 22949 26632 22995 26678
rect 22949 26527 22995 26573
rect 22949 26422 22995 26468
rect 22949 26317 22995 26363
rect 22949 26212 22995 26258
rect 22949 26107 22995 26153
rect 22949 26002 22995 26048
rect 22949 25897 22995 25943
rect 22949 25792 22995 25838
rect 22949 25687 22995 25733
rect 22949 25582 22995 25628
rect 22949 25478 22995 25524
rect 22949 25374 22995 25420
rect 22949 25270 22995 25316
rect 22949 25166 22995 25212
rect 22949 25062 22995 25108
rect 22949 24958 22995 25004
rect 22949 24854 22995 24900
rect 23956 25088 24002 25134
rect 23956 24985 24002 25031
rect 23956 24882 24002 24928
rect 22949 24750 22995 24796
rect 22949 24646 22995 24692
rect 15899 23324 15945 23370
rect 15899 23221 15945 23267
rect 15899 23118 15945 23164
rect 15899 23015 15945 23061
rect 15899 22912 15945 22958
rect 15899 22809 15945 22855
rect 15899 22706 15945 22752
rect 15899 22603 15945 22649
rect 15899 22500 15945 22546
rect 15899 22397 15945 22443
rect 16704 21924 16750 23984
rect 16928 21924 16974 23984
rect 17152 21924 17198 23984
rect 17376 21924 17422 23984
rect 17600 21924 17646 23984
rect 17824 21924 17870 23984
rect 18048 21924 18094 23984
rect 18338 21924 18384 23984
rect 18562 21924 18608 23984
rect 18786 21924 18832 23984
rect 19010 21924 19056 23984
rect 19234 21924 19280 23984
rect 19458 21924 19504 23984
rect 19682 21924 19728 23984
rect 19971 21924 20017 23984
rect 20195 21924 20241 23984
rect 20419 21924 20465 23984
rect 20643 21924 20689 23984
rect 20867 21924 20913 23984
rect 21091 21924 21137 23984
rect 21315 21924 21361 23984
rect 21605 21924 21651 23984
rect 21829 21924 21875 23984
rect 22053 21924 22099 23984
rect 22277 21924 22323 23984
rect 22501 21924 22547 23984
rect 22725 21924 22771 23984
rect 22949 21924 22995 23984
rect 23956 24779 24002 24825
rect 23956 24676 24002 24722
rect 23956 24573 24002 24619
rect 23956 24470 24002 24516
rect 23956 24367 24002 24413
rect 23956 24264 24002 24310
rect 23956 24161 24002 24207
rect 23956 24058 24002 24104
rect 23956 23955 24002 24001
rect 23956 23852 24002 23898
rect 23956 23749 24002 23795
rect 23956 23646 24002 23692
rect 23956 23543 24002 23589
rect 23956 23440 24002 23486
rect 23956 23337 24002 23383
rect 23956 23234 24002 23280
rect 23956 23131 24002 23177
rect 23956 23028 24002 23074
rect 23956 22925 24002 22971
rect 23956 22822 24002 22868
rect 23956 22719 24002 22765
rect 23956 22616 24002 22662
rect 23956 22513 24002 22559
rect 23956 22410 24002 22456
rect 23956 22307 24002 22353
rect 23956 22204 24002 22250
rect 23956 22101 24002 22147
rect 23956 21998 24002 22044
rect 23956 21894 24002 21940
rect 24180 25088 24226 25134
rect 24180 24985 24226 25031
rect 24180 24882 24226 24928
rect 24180 24779 24226 24825
rect 24180 24676 24226 24722
rect 24180 24573 24226 24619
rect 24180 24470 24226 24516
rect 24180 24367 24226 24413
rect 24180 24264 24226 24310
rect 24180 24161 24226 24207
rect 24180 24058 24226 24104
rect 24180 23955 24226 24001
rect 24180 23852 24226 23898
rect 24180 23749 24226 23795
rect 24180 23646 24226 23692
rect 24180 23543 24226 23589
rect 24180 23440 24226 23486
rect 24180 23337 24226 23383
rect 24180 23234 24226 23280
rect 24180 23131 24226 23177
rect 24180 23028 24226 23074
rect 24180 22925 24226 22971
rect 24180 22822 24226 22868
rect 24180 22719 24226 22765
rect 24180 22616 24226 22662
rect 24180 22513 24226 22559
rect 24180 22410 24226 22456
rect 24180 22307 24226 22353
rect 24180 22204 24226 22250
rect 24180 22101 24226 22147
rect 24180 21998 24226 22044
rect 24180 21894 24226 21940
rect 24470 25088 24516 25134
rect 24470 24985 24516 25031
rect 24470 24882 24516 24928
rect 24470 24779 24516 24825
rect 24470 24676 24516 24722
rect 24470 24573 24516 24619
rect 24470 24470 24516 24516
rect 24470 24367 24516 24413
rect 24470 24264 24516 24310
rect 24470 24161 24516 24207
rect 24470 24058 24516 24104
rect 24470 23955 24516 24001
rect 24470 23852 24516 23898
rect 24470 23749 24516 23795
rect 24470 23646 24516 23692
rect 24470 23543 24516 23589
rect 24470 23440 24516 23486
rect 24470 23337 24516 23383
rect 24470 23234 24516 23280
rect 24470 23131 24516 23177
rect 24470 23028 24516 23074
rect 24470 22925 24516 22971
rect 24470 22822 24516 22868
rect 24470 22719 24516 22765
rect 24470 22616 24516 22662
rect 24470 22513 24516 22559
rect 24470 22410 24516 22456
rect 24470 22307 24516 22353
rect 24470 22204 24516 22250
rect 24470 22101 24516 22147
rect 24470 21998 24516 22044
rect 24470 21894 24516 21940
rect 24694 25088 24740 25134
rect 24694 24985 24740 25031
rect 24694 24882 24740 24928
rect 24694 24779 24740 24825
rect 25646 25088 25692 25134
rect 25646 24985 25692 25031
rect 25646 24882 25692 24928
rect 24694 24676 24740 24722
rect 24694 24573 24740 24619
rect 24694 24470 24740 24516
rect 24694 24367 24740 24413
rect 24694 24264 24740 24310
rect 24694 24161 24740 24207
rect 24694 24058 24740 24104
rect 24694 23955 24740 24001
rect 24694 23852 24740 23898
rect 24694 23749 24740 23795
rect 24694 23646 24740 23692
rect 24694 23543 24740 23589
rect 24694 23440 24740 23486
rect 24694 23337 24740 23383
rect 24694 23234 24740 23280
rect 24694 23131 24740 23177
rect 24694 23028 24740 23074
rect 24694 22925 24740 22971
rect 24694 22822 24740 22868
rect 24694 22719 24740 22765
rect 24694 22616 24740 22662
rect 24694 22513 24740 22559
rect 24694 22410 24740 22456
rect 24694 22307 24740 22353
rect 24694 22204 24740 22250
rect 24694 22101 24740 22147
rect 24694 21998 24740 22044
rect 24694 21894 24740 21940
rect 25646 24779 25692 24825
rect 25646 24676 25692 24722
rect 25646 24573 25692 24619
rect 25646 24470 25692 24516
rect 25646 24367 25692 24413
rect 25646 24264 25692 24310
rect 25646 24161 25692 24207
rect 25646 24058 25692 24104
rect 25646 23955 25692 24001
rect 25646 23852 25692 23898
rect 25646 23749 25692 23795
rect 25646 23646 25692 23692
rect 25646 23543 25692 23589
rect 25646 23440 25692 23486
rect 25646 23337 25692 23383
rect 25646 23234 25692 23280
rect 25646 23131 25692 23177
rect 25646 23028 25692 23074
rect 25646 22925 25692 22971
rect 25646 22822 25692 22868
rect 25646 22719 25692 22765
rect 25646 22616 25692 22662
rect 25646 22513 25692 22559
rect 25646 22410 25692 22456
rect 25646 22307 25692 22353
rect 25646 22204 25692 22250
rect 25646 22101 25692 22147
rect 25646 21998 25692 22044
rect 25646 21894 25692 21940
rect 25870 25088 25916 25134
rect 25870 24985 25916 25031
rect 25870 24882 25916 24928
rect 25870 24779 25916 24825
rect 25870 24676 25916 24722
rect 25870 24573 25916 24619
rect 25870 24470 25916 24516
rect 25870 24367 25916 24413
rect 25870 24264 25916 24310
rect 25870 24161 25916 24207
rect 25870 24058 25916 24104
rect 25870 23955 25916 24001
rect 25870 23852 25916 23898
rect 25870 23749 25916 23795
rect 25870 23646 25916 23692
rect 25870 23543 25916 23589
rect 25870 23440 25916 23486
rect 25870 23337 25916 23383
rect 25870 23234 25916 23280
rect 25870 23131 25916 23177
rect 25870 23028 25916 23074
rect 25870 22925 25916 22971
rect 25870 22822 25916 22868
rect 25870 22719 25916 22765
rect 25870 22616 25916 22662
rect 25870 22513 25916 22559
rect 25870 22410 25916 22456
rect 25870 22307 25916 22353
rect 25870 22204 25916 22250
rect 25870 22101 25916 22147
rect 25870 21998 25916 22044
rect 25870 21894 25916 21940
rect 26160 25088 26206 25134
rect 26160 24985 26206 25031
rect 26160 24882 26206 24928
rect 26160 24779 26206 24825
rect 26160 24676 26206 24722
rect 26160 24573 26206 24619
rect 26160 24470 26206 24516
rect 26160 24367 26206 24413
rect 26160 24264 26206 24310
rect 26160 24161 26206 24207
rect 26160 24058 26206 24104
rect 26160 23955 26206 24001
rect 26160 23852 26206 23898
rect 26160 23749 26206 23795
rect 26160 23646 26206 23692
rect 26160 23543 26206 23589
rect 26160 23440 26206 23486
rect 26160 23337 26206 23383
rect 26160 23234 26206 23280
rect 26160 23131 26206 23177
rect 26160 23028 26206 23074
rect 26160 22925 26206 22971
rect 26160 22822 26206 22868
rect 26160 22719 26206 22765
rect 26160 22616 26206 22662
rect 26160 22513 26206 22559
rect 26160 22410 26206 22456
rect 26160 22307 26206 22353
rect 26160 22204 26206 22250
rect 26160 22101 26206 22147
rect 26160 21998 26206 22044
rect 26160 21894 26206 21940
rect 26384 25088 26430 25134
rect 26384 24985 26430 25031
rect 26384 24882 26430 24928
rect 26384 24779 26430 24825
rect 27337 25088 27383 25134
rect 27337 24985 27383 25031
rect 27337 24882 27383 24928
rect 26384 24676 26430 24722
rect 26384 24573 26430 24619
rect 26384 24470 26430 24516
rect 26384 24367 26430 24413
rect 26384 24264 26430 24310
rect 26384 24161 26430 24207
rect 26384 24058 26430 24104
rect 26384 23955 26430 24001
rect 26384 23852 26430 23898
rect 26384 23749 26430 23795
rect 26384 23646 26430 23692
rect 26384 23543 26430 23589
rect 26384 23440 26430 23486
rect 26384 23337 26430 23383
rect 26384 23234 26430 23280
rect 26384 23131 26430 23177
rect 26384 23028 26430 23074
rect 26384 22925 26430 22971
rect 26384 22822 26430 22868
rect 26384 22719 26430 22765
rect 26384 22616 26430 22662
rect 26384 22513 26430 22559
rect 26384 22410 26430 22456
rect 26384 22307 26430 22353
rect 26384 22204 26430 22250
rect 26384 22101 26430 22147
rect 26384 21998 26430 22044
rect 26384 21894 26430 21940
rect 27337 24779 27383 24825
rect 27337 24676 27383 24722
rect 27337 24573 27383 24619
rect 27337 24470 27383 24516
rect 27337 24367 27383 24413
rect 27337 24264 27383 24310
rect 27337 24161 27383 24207
rect 27337 24058 27383 24104
rect 27337 23955 27383 24001
rect 27337 23852 27383 23898
rect 27337 23749 27383 23795
rect 27337 23646 27383 23692
rect 27337 23543 27383 23589
rect 27337 23440 27383 23486
rect 27337 23337 27383 23383
rect 27337 23234 27383 23280
rect 27337 23131 27383 23177
rect 27337 23028 27383 23074
rect 27337 22925 27383 22971
rect 27337 22822 27383 22868
rect 27337 22719 27383 22765
rect 27337 22616 27383 22662
rect 27337 22513 27383 22559
rect 27337 22410 27383 22456
rect 27337 22307 27383 22353
rect 27337 22204 27383 22250
rect 27337 22101 27383 22147
rect 27337 21998 27383 22044
rect 27337 21894 27383 21940
rect 27561 25088 27607 25134
rect 27561 24985 27607 25031
rect 27561 24882 27607 24928
rect 27561 24779 27607 24825
rect 27561 24676 27607 24722
rect 27561 24573 27607 24619
rect 27561 24470 27607 24516
rect 27561 24367 27607 24413
rect 27561 24264 27607 24310
rect 27561 24161 27607 24207
rect 27561 24058 27607 24104
rect 27561 23955 27607 24001
rect 27561 23852 27607 23898
rect 27561 23749 27607 23795
rect 27561 23646 27607 23692
rect 27561 23543 27607 23589
rect 27561 23440 27607 23486
rect 27561 23337 27607 23383
rect 27561 23234 27607 23280
rect 27561 23131 27607 23177
rect 27561 23028 27607 23074
rect 27561 22925 27607 22971
rect 27561 22822 27607 22868
rect 27561 22719 27607 22765
rect 27561 22616 27607 22662
rect 27561 22513 27607 22559
rect 27561 22410 27607 22456
rect 27561 22307 27607 22353
rect 27561 22204 27607 22250
rect 27561 22101 27607 22147
rect 27561 21998 27607 22044
rect 27561 21894 27607 21940
rect 27851 25088 27897 25134
rect 27851 24985 27897 25031
rect 27851 24882 27897 24928
rect 27851 24779 27897 24825
rect 27851 24676 27897 24722
rect 27851 24573 27897 24619
rect 27851 24470 27897 24516
rect 27851 24367 27897 24413
rect 27851 24264 27897 24310
rect 27851 24161 27897 24207
rect 27851 24058 27897 24104
rect 27851 23955 27897 24001
rect 27851 23852 27897 23898
rect 27851 23749 27897 23795
rect 27851 23646 27897 23692
rect 27851 23543 27897 23589
rect 27851 23440 27897 23486
rect 27851 23337 27897 23383
rect 27851 23234 27897 23280
rect 27851 23131 27897 23177
rect 27851 23028 27897 23074
rect 27851 22925 27897 22971
rect 27851 22822 27897 22868
rect 27851 22719 27897 22765
rect 27851 22616 27897 22662
rect 27851 22513 27897 22559
rect 27851 22410 27897 22456
rect 27851 22307 27897 22353
rect 27851 22204 27897 22250
rect 27851 22101 27897 22147
rect 27851 21998 27897 22044
rect 27851 21894 27897 21940
rect 28075 25088 28121 25134
rect 28075 24985 28121 25031
rect 28075 24882 28121 24928
rect 28075 24779 28121 24825
rect 28075 24676 28121 24722
rect 28075 24573 28121 24619
rect 28075 24470 28121 24516
rect 28075 24367 28121 24413
rect 28075 24264 28121 24310
rect 28075 24161 28121 24207
rect 28075 24058 28121 24104
rect 28075 23955 28121 24001
rect 28075 23852 28121 23898
rect 28075 23749 28121 23795
rect 28075 23646 28121 23692
rect 28075 23543 28121 23589
rect 28075 23440 28121 23486
rect 28075 23337 28121 23383
rect 28075 23234 28121 23280
rect 28075 23131 28121 23177
rect 28075 23028 28121 23074
rect 28075 22925 28121 22971
rect 28075 22822 28121 22868
rect 28075 22719 28121 22765
rect 28075 22616 28121 22662
rect 28075 22513 28121 22559
rect 28075 22410 28121 22456
rect 28075 22307 28121 22353
rect 28075 22204 28121 22250
rect 28075 22101 28121 22147
rect 28075 21998 28121 22044
rect 28075 21894 28121 21940
rect 1995 12598 2041 16572
rect 2219 12598 2265 16572
rect 2443 12598 2489 16572
rect 2667 12598 2713 16572
rect 2891 12598 2937 16572
rect 3115 12598 3161 16572
rect 3339 12598 3385 16572
rect 3563 12598 3609 16572
rect 3787 12598 3833 16572
rect 4011 12598 4057 16572
rect 4235 12598 4281 16572
rect 4459 12598 4505 16572
rect 4683 12598 4729 16572
rect 4907 12598 4953 16572
rect 5131 12598 5177 16572
rect 5355 12598 5401 16572
rect 5579 12598 5625 16572
rect 5803 12598 5849 16572
rect 6027 12598 6073 16572
rect 6251 12598 6297 16572
rect 6475 12598 6521 16572
rect 6699 12598 6745 16572
rect 6923 12598 6969 16572
rect 7147 12598 7193 16572
rect 7371 12598 7417 16572
rect 7595 12598 7641 16572
rect 7819 12598 7865 16572
rect 8043 12598 8089 16572
rect 8267 12598 8313 16572
rect 8491 12598 8537 16572
rect 8715 12598 8761 16572
rect 8939 12598 8985 16572
rect 9163 12598 9209 16572
rect 9387 12598 9433 16572
rect 9611 12598 9657 16572
rect 9835 12598 9881 16572
rect 10059 12598 10105 16572
rect 10283 12598 10329 16572
rect 10507 12598 10553 16572
rect 10731 12598 10777 16572
rect 10955 12598 11001 16572
rect 11179 12598 11225 16572
rect 11403 12598 11449 16572
rect 11627 12598 11673 16572
rect 11851 12598 11897 16572
rect 12075 12598 12121 16572
rect 12299 12598 12345 16572
rect 12523 12598 12569 16572
rect 12747 12598 12793 16572
rect 12971 12598 13017 16572
rect 13195 12598 13241 16572
rect 13419 12598 13465 16572
rect 13643 12598 13689 16572
rect 13867 12598 13913 16572
rect 14091 12598 14137 16572
rect 14315 12598 14361 16572
rect 14539 12598 14585 16572
rect 14763 12598 14809 16572
rect 14987 12598 15033 16572
rect 15211 12598 15257 16572
rect 15435 12598 15481 16572
rect 15659 12598 15705 16572
rect 15883 12598 15929 16572
rect 16107 12598 16153 16572
rect 16331 12598 16377 16572
rect 16555 12598 16601 16572
rect 16779 12598 16825 16572
rect 17003 12598 17049 16572
rect 17227 12598 17273 16572
rect 17451 12598 17497 16572
rect 17675 12598 17721 16572
rect 17899 12598 17945 16572
rect 18123 12598 18169 16572
rect 18347 12598 18393 16572
rect 18571 12598 18617 16572
rect 18795 12598 18841 16572
rect 19019 12598 19065 16572
rect 19243 12598 19289 16572
rect 19467 12598 19513 16572
rect 19691 12598 19737 16572
rect 19915 12598 19961 16572
rect 7450 8227 7496 8273
rect 7450 8118 7496 8164
rect 7450 8009 7496 8055
rect 2621 5268 2667 7964
rect 2845 5268 2891 7964
rect 3135 5268 3181 7964
rect 3359 5268 3405 7964
rect 4312 5268 4358 7964
rect 4536 5268 4582 7964
rect 4826 5268 4872 7964
rect 5050 5268 5096 7964
rect 6003 5268 6049 7964
rect 6227 5268 6273 7964
rect 6517 5268 6563 7964
rect 6741 5268 6787 7964
rect 7450 7901 7496 7947
rect 7450 7793 7496 7839
rect 7450 7685 7496 7731
rect 7450 7577 7496 7623
rect 7450 7469 7496 7515
rect 7450 7361 7496 7407
rect 7450 7253 7496 7299
rect 7450 7145 7496 7191
rect 7674 8227 7720 8273
rect 7674 8118 7720 8164
rect 7674 8009 7720 8055
rect 7674 7901 7720 7947
rect 7674 7793 7720 7839
rect 7674 7685 7720 7731
rect 7674 7577 7720 7623
rect 7674 7469 7720 7515
rect 7674 7361 7720 7407
rect 7674 7253 7720 7299
rect 7674 7145 7720 7191
rect 7898 8227 7944 8273
rect 7898 8118 7944 8164
rect 7898 8009 7944 8055
rect 7898 7901 7944 7947
rect 7898 7793 7944 7839
rect 7898 7685 7944 7731
rect 7898 7577 7944 7623
rect 7898 7469 7944 7515
rect 7898 7361 7944 7407
rect 7898 7253 7944 7299
rect 7898 7145 7944 7191
rect 8122 8227 8168 8273
rect 8122 8118 8168 8164
rect 8122 8009 8168 8055
rect 8122 7901 8168 7947
rect 8122 7793 8168 7839
rect 8122 7685 8168 7731
rect 8122 7577 8168 7623
rect 8122 7469 8168 7515
rect 8122 7361 8168 7407
rect 8122 7253 8168 7299
rect 8122 7145 8168 7191
rect 8346 8227 8392 8273
rect 8346 8118 8392 8164
rect 8346 8009 8392 8055
rect 8346 7901 8392 7947
rect 8346 7793 8392 7839
rect 8346 7685 8392 7731
rect 8346 7577 8392 7623
rect 8346 7469 8392 7515
rect 8346 7361 8392 7407
rect 8346 7253 8392 7299
rect 8346 7145 8392 7191
rect 8570 8227 8616 8273
rect 8570 8118 8616 8164
rect 8570 8009 8616 8055
rect 8570 7901 8616 7947
rect 8570 7793 8616 7839
rect 8570 7685 8616 7731
rect 8570 7577 8616 7623
rect 8570 7469 8616 7515
rect 8570 7361 8616 7407
rect 8570 7253 8616 7299
rect 8570 7145 8616 7191
rect 8794 8227 8840 8273
rect 8794 8118 8840 8164
rect 8794 8009 8840 8055
rect 8794 7901 8840 7947
rect 8794 7793 8840 7839
rect 8794 7685 8840 7731
rect 8794 7577 8840 7623
rect 8794 7469 8840 7515
rect 8794 7361 8840 7407
rect 8794 7253 8840 7299
rect 8794 7145 8840 7191
rect 9083 8227 9129 8273
rect 9083 8118 9129 8164
rect 9083 8009 9129 8055
rect 9083 7901 9129 7947
rect 9083 7793 9129 7839
rect 9083 7685 9129 7731
rect 9083 7577 9129 7623
rect 9083 7469 9129 7515
rect 9083 7361 9129 7407
rect 9083 7253 9129 7299
rect 9083 7145 9129 7191
rect 9307 8227 9353 8273
rect 9307 8118 9353 8164
rect 9307 8009 9353 8055
rect 9307 7901 9353 7947
rect 9307 7793 9353 7839
rect 9307 7685 9353 7731
rect 9307 7577 9353 7623
rect 9307 7469 9353 7515
rect 9307 7361 9353 7407
rect 9307 7253 9353 7299
rect 9307 7145 9353 7191
rect 9531 8227 9577 8273
rect 9531 8118 9577 8164
rect 9531 8009 9577 8055
rect 9531 7901 9577 7947
rect 9531 7793 9577 7839
rect 9531 7685 9577 7731
rect 9531 7577 9577 7623
rect 9531 7469 9577 7515
rect 9531 7361 9577 7407
rect 9531 7253 9577 7299
rect 9531 7145 9577 7191
rect 9755 8227 9801 8273
rect 9755 8118 9801 8164
rect 9755 8009 9801 8055
rect 9755 7901 9801 7947
rect 9755 7793 9801 7839
rect 9755 7685 9801 7731
rect 9755 7577 9801 7623
rect 9755 7469 9801 7515
rect 9755 7361 9801 7407
rect 9755 7253 9801 7299
rect 9755 7145 9801 7191
rect 9979 8227 10025 8273
rect 9979 8118 10025 8164
rect 9979 8009 10025 8055
rect 9979 7901 10025 7947
rect 9979 7793 10025 7839
rect 9979 7685 10025 7731
rect 9979 7577 10025 7623
rect 9979 7469 10025 7515
rect 9979 7361 10025 7407
rect 9979 7253 10025 7299
rect 9979 7145 10025 7191
rect 10203 8227 10249 8273
rect 10203 8118 10249 8164
rect 10203 8009 10249 8055
rect 10203 7901 10249 7947
rect 10203 7793 10249 7839
rect 10203 7685 10249 7731
rect 10203 7577 10249 7623
rect 10203 7469 10249 7515
rect 10203 7361 10249 7407
rect 10203 7253 10249 7299
rect 10203 7145 10249 7191
rect 10427 8227 10473 8273
rect 10427 8118 10473 8164
rect 10427 8009 10473 8055
rect 10427 7901 10473 7947
rect 10427 7793 10473 7839
rect 10427 7685 10473 7731
rect 10427 7577 10473 7623
rect 10427 7469 10473 7515
rect 10427 7361 10473 7407
rect 10427 7253 10473 7299
rect 10427 7145 10473 7191
rect 10717 8227 10763 8273
rect 10717 8118 10763 8164
rect 10717 8009 10763 8055
rect 10717 7901 10763 7947
rect 10717 7793 10763 7839
rect 10717 7685 10763 7731
rect 10717 7577 10763 7623
rect 10717 7469 10763 7515
rect 10717 7361 10763 7407
rect 10717 7253 10763 7299
rect 10717 7145 10763 7191
rect 10941 8227 10987 8273
rect 10941 8118 10987 8164
rect 10941 8009 10987 8055
rect 10941 7901 10987 7947
rect 10941 7793 10987 7839
rect 10941 7685 10987 7731
rect 10941 7577 10987 7623
rect 10941 7469 10987 7515
rect 10941 7361 10987 7407
rect 10941 7253 10987 7299
rect 10941 7145 10987 7191
rect 11165 8227 11211 8273
rect 11165 8118 11211 8164
rect 11165 8009 11211 8055
rect 11165 7901 11211 7947
rect 11165 7793 11211 7839
rect 11165 7685 11211 7731
rect 11165 7577 11211 7623
rect 11165 7469 11211 7515
rect 11165 7361 11211 7407
rect 11165 7253 11211 7299
rect 11165 7145 11211 7191
rect 11389 8227 11435 8273
rect 11389 8118 11435 8164
rect 11389 8009 11435 8055
rect 11389 7901 11435 7947
rect 11389 7793 11435 7839
rect 11389 7685 11435 7731
rect 11389 7577 11435 7623
rect 11389 7469 11435 7515
rect 11389 7361 11435 7407
rect 11389 7253 11435 7299
rect 11389 7145 11435 7191
rect 11613 8227 11659 8273
rect 11613 8118 11659 8164
rect 11613 8009 11659 8055
rect 11613 7901 11659 7947
rect 11613 7793 11659 7839
rect 11613 7685 11659 7731
rect 11613 7577 11659 7623
rect 11613 7469 11659 7515
rect 11613 7361 11659 7407
rect 11613 7253 11659 7299
rect 11613 7145 11659 7191
rect 11837 8227 11883 8273
rect 11837 8118 11883 8164
rect 11837 8009 11883 8055
rect 11837 7901 11883 7947
rect 11837 7793 11883 7839
rect 11837 7685 11883 7731
rect 11837 7577 11883 7623
rect 11837 7469 11883 7515
rect 11837 7361 11883 7407
rect 11837 7253 11883 7299
rect 11837 7145 11883 7191
rect 12061 8227 12107 8273
rect 12061 8118 12107 8164
rect 12061 8009 12107 8055
rect 12061 7901 12107 7947
rect 12061 7793 12107 7839
rect 12061 7685 12107 7731
rect 12061 7577 12107 7623
rect 12061 7469 12107 7515
rect 12061 7361 12107 7407
rect 12061 7253 12107 7299
rect 12061 7145 12107 7191
rect 12351 8227 12397 8273
rect 12351 8118 12397 8164
rect 12351 8009 12397 8055
rect 12351 7901 12397 7947
rect 12351 7793 12397 7839
rect 12351 7685 12397 7731
rect 12351 7577 12397 7623
rect 12351 7469 12397 7515
rect 12351 7361 12397 7407
rect 12351 7253 12397 7299
rect 12351 7145 12397 7191
rect 12575 8227 12621 8273
rect 12575 8118 12621 8164
rect 12575 8009 12621 8055
rect 12575 7901 12621 7947
rect 12575 7793 12621 7839
rect 12575 7685 12621 7731
rect 12575 7577 12621 7623
rect 12575 7469 12621 7515
rect 12575 7361 12621 7407
rect 12575 7253 12621 7299
rect 12575 7145 12621 7191
rect 12799 8227 12845 8273
rect 12799 8118 12845 8164
rect 12799 8009 12845 8055
rect 12799 7901 12845 7947
rect 12799 7793 12845 7839
rect 12799 7685 12845 7731
rect 12799 7577 12845 7623
rect 12799 7469 12845 7515
rect 12799 7361 12845 7407
rect 12799 7253 12845 7299
rect 12799 7145 12845 7191
rect 13023 8227 13069 8273
rect 13023 8118 13069 8164
rect 13023 8009 13069 8055
rect 13023 7901 13069 7947
rect 13023 7793 13069 7839
rect 13023 7685 13069 7731
rect 13023 7577 13069 7623
rect 13023 7469 13069 7515
rect 13023 7361 13069 7407
rect 13023 7253 13069 7299
rect 13023 7145 13069 7191
rect 13247 8227 13293 8273
rect 13247 8118 13293 8164
rect 13247 8009 13293 8055
rect 13247 7901 13293 7947
rect 13247 7793 13293 7839
rect 13247 7685 13293 7731
rect 13247 7577 13293 7623
rect 13247 7469 13293 7515
rect 13247 7361 13293 7407
rect 13247 7253 13293 7299
rect 13247 7145 13293 7191
rect 13471 8227 13517 8273
rect 13471 8118 13517 8164
rect 13471 8009 13517 8055
rect 13471 7901 13517 7947
rect 13471 7793 13517 7839
rect 13471 7685 13517 7731
rect 13471 7577 13517 7623
rect 13471 7469 13517 7515
rect 13471 7361 13517 7407
rect 13471 7253 13517 7299
rect 13471 7145 13517 7191
rect 13695 8227 13741 8273
rect 13695 8118 13741 8164
rect 13695 8009 13741 8055
rect 13695 7901 13741 7947
rect 13695 7793 13741 7839
rect 13695 7685 13741 7731
rect 13695 7577 13741 7623
rect 13695 7469 13741 7515
rect 13695 7361 13741 7407
rect 13695 7253 13741 7299
rect 13695 7145 13741 7191
rect 7450 6360 7496 6406
rect 7450 6254 7496 6300
rect 7450 6148 7496 6194
rect 7450 6042 7496 6088
rect 7450 5936 7496 5982
rect 7450 5830 7496 5876
rect 7450 5724 7496 5770
rect 7450 5618 7496 5664
rect 7450 5512 7496 5558
rect 7450 5405 7496 5451
rect 7450 5298 7496 5344
rect 7674 6360 7720 6406
rect 7674 6254 7720 6300
rect 7674 6148 7720 6194
rect 7674 6042 7720 6088
rect 7674 5936 7720 5982
rect 7674 5830 7720 5876
rect 7674 5724 7720 5770
rect 7674 5618 7720 5664
rect 7674 5512 7720 5558
rect 7674 5405 7720 5451
rect 7674 5298 7720 5344
rect 7898 6360 7944 6406
rect 7898 6254 7944 6300
rect 7898 6148 7944 6194
rect 7898 6042 7944 6088
rect 7898 5936 7944 5982
rect 7898 5830 7944 5876
rect 7898 5724 7944 5770
rect 7898 5618 7944 5664
rect 7898 5512 7944 5558
rect 7898 5405 7944 5451
rect 7898 5298 7944 5344
rect 8122 6360 8168 6406
rect 8122 6254 8168 6300
rect 8122 6148 8168 6194
rect 8122 6042 8168 6088
rect 8122 5936 8168 5982
rect 8122 5830 8168 5876
rect 8122 5724 8168 5770
rect 8122 5618 8168 5664
rect 8122 5512 8168 5558
rect 8122 5405 8168 5451
rect 8122 5298 8168 5344
rect 8346 6360 8392 6406
rect 8346 6254 8392 6300
rect 8346 6148 8392 6194
rect 8346 6042 8392 6088
rect 8346 5936 8392 5982
rect 8346 5830 8392 5876
rect 8346 5724 8392 5770
rect 8346 5618 8392 5664
rect 8346 5512 8392 5558
rect 8346 5405 8392 5451
rect 8346 5298 8392 5344
rect 8570 6360 8616 6406
rect 8570 6254 8616 6300
rect 8570 6148 8616 6194
rect 8570 6042 8616 6088
rect 8570 5936 8616 5982
rect 8570 5830 8616 5876
rect 8570 5724 8616 5770
rect 8570 5618 8616 5664
rect 8570 5512 8616 5558
rect 8570 5405 8616 5451
rect 8570 5298 8616 5344
rect 8794 6360 8840 6406
rect 8794 6254 8840 6300
rect 8794 6148 8840 6194
rect 8794 6042 8840 6088
rect 8794 5936 8840 5982
rect 8794 5830 8840 5876
rect 8794 5724 8840 5770
rect 8794 5618 8840 5664
rect 8794 5512 8840 5558
rect 8794 5405 8840 5451
rect 8794 5298 8840 5344
rect 9083 6360 9129 6406
rect 9083 6254 9129 6300
rect 9083 6148 9129 6194
rect 9083 6042 9129 6088
rect 9083 5936 9129 5982
rect 9083 5830 9129 5876
rect 9083 5724 9129 5770
rect 9083 5618 9129 5664
rect 9083 5512 9129 5558
rect 9083 5405 9129 5451
rect 9083 5298 9129 5344
rect 9307 6360 9353 6406
rect 9307 6254 9353 6300
rect 9307 6148 9353 6194
rect 9307 6042 9353 6088
rect 9307 5936 9353 5982
rect 9307 5830 9353 5876
rect 9307 5724 9353 5770
rect 9307 5618 9353 5664
rect 9307 5512 9353 5558
rect 9307 5405 9353 5451
rect 9307 5298 9353 5344
rect 9531 6360 9577 6406
rect 9531 6254 9577 6300
rect 9531 6148 9577 6194
rect 9531 6042 9577 6088
rect 9531 5936 9577 5982
rect 9531 5830 9577 5876
rect 9531 5724 9577 5770
rect 9531 5618 9577 5664
rect 9531 5512 9577 5558
rect 9531 5405 9577 5451
rect 9531 5298 9577 5344
rect 9755 6360 9801 6406
rect 9755 6254 9801 6300
rect 9755 6148 9801 6194
rect 9755 6042 9801 6088
rect 9755 5936 9801 5982
rect 9755 5830 9801 5876
rect 9755 5724 9801 5770
rect 9755 5618 9801 5664
rect 9755 5512 9801 5558
rect 9755 5405 9801 5451
rect 9755 5298 9801 5344
rect 9979 6360 10025 6406
rect 9979 6254 10025 6300
rect 9979 6148 10025 6194
rect 9979 6042 10025 6088
rect 9979 5936 10025 5982
rect 9979 5830 10025 5876
rect 9979 5724 10025 5770
rect 9979 5618 10025 5664
rect 9979 5512 10025 5558
rect 9979 5405 10025 5451
rect 9979 5298 10025 5344
rect 10203 6360 10249 6406
rect 10203 6254 10249 6300
rect 10203 6148 10249 6194
rect 10203 6042 10249 6088
rect 10203 5936 10249 5982
rect 10203 5830 10249 5876
rect 10203 5724 10249 5770
rect 10203 5618 10249 5664
rect 10203 5512 10249 5558
rect 10203 5405 10249 5451
rect 10203 5298 10249 5344
rect 10427 6360 10473 6406
rect 10427 6254 10473 6300
rect 10427 6148 10473 6194
rect 10427 6042 10473 6088
rect 10427 5936 10473 5982
rect 10427 5830 10473 5876
rect 10427 5724 10473 5770
rect 10427 5618 10473 5664
rect 10427 5512 10473 5558
rect 10427 5405 10473 5451
rect 10427 5298 10473 5344
rect 10717 6360 10763 6406
rect 10717 6254 10763 6300
rect 10717 6148 10763 6194
rect 10717 6042 10763 6088
rect 10717 5936 10763 5982
rect 10717 5830 10763 5876
rect 10717 5724 10763 5770
rect 10717 5618 10763 5664
rect 10717 5512 10763 5558
rect 10717 5405 10763 5451
rect 10717 5298 10763 5344
rect 10941 6360 10987 6406
rect 10941 6254 10987 6300
rect 10941 6148 10987 6194
rect 10941 6042 10987 6088
rect 10941 5936 10987 5982
rect 10941 5830 10987 5876
rect 10941 5724 10987 5770
rect 10941 5618 10987 5664
rect 10941 5512 10987 5558
rect 10941 5405 10987 5451
rect 10941 5298 10987 5344
rect 11165 6360 11211 6406
rect 11165 6254 11211 6300
rect 11165 6148 11211 6194
rect 11165 6042 11211 6088
rect 11165 5936 11211 5982
rect 11165 5830 11211 5876
rect 11165 5724 11211 5770
rect 11165 5618 11211 5664
rect 11165 5512 11211 5558
rect 11165 5405 11211 5451
rect 11165 5298 11211 5344
rect 11389 6360 11435 6406
rect 11389 6254 11435 6300
rect 11389 6148 11435 6194
rect 11389 6042 11435 6088
rect 11389 5936 11435 5982
rect 11389 5830 11435 5876
rect 11389 5724 11435 5770
rect 11389 5618 11435 5664
rect 11389 5512 11435 5558
rect 11389 5405 11435 5451
rect 11389 5298 11435 5344
rect 11613 6360 11659 6406
rect 11613 6254 11659 6300
rect 11613 6148 11659 6194
rect 11613 6042 11659 6088
rect 11613 5936 11659 5982
rect 11613 5830 11659 5876
rect 11613 5724 11659 5770
rect 11613 5618 11659 5664
rect 11613 5512 11659 5558
rect 11613 5405 11659 5451
rect 11613 5298 11659 5344
rect 11837 6360 11883 6406
rect 11837 6254 11883 6300
rect 11837 6148 11883 6194
rect 11837 6042 11883 6088
rect 11837 5936 11883 5982
rect 11837 5830 11883 5876
rect 11837 5724 11883 5770
rect 11837 5618 11883 5664
rect 11837 5512 11883 5558
rect 11837 5405 11883 5451
rect 11837 5298 11883 5344
rect 12061 6360 12107 6406
rect 12061 6254 12107 6300
rect 12061 6148 12107 6194
rect 12061 6042 12107 6088
rect 12061 5936 12107 5982
rect 12061 5830 12107 5876
rect 12061 5724 12107 5770
rect 12061 5618 12107 5664
rect 12061 5512 12107 5558
rect 12061 5405 12107 5451
rect 12061 5298 12107 5344
rect 12351 6360 12397 6406
rect 12351 6254 12397 6300
rect 12351 6148 12397 6194
rect 12351 6042 12397 6088
rect 12351 5936 12397 5982
rect 12351 5830 12397 5876
rect 12351 5724 12397 5770
rect 12351 5618 12397 5664
rect 12351 5512 12397 5558
rect 12351 5405 12397 5451
rect 12351 5298 12397 5344
rect 12575 6360 12621 6406
rect 12575 6254 12621 6300
rect 12575 6148 12621 6194
rect 12575 6042 12621 6088
rect 12575 5936 12621 5982
rect 12575 5830 12621 5876
rect 12575 5724 12621 5770
rect 12575 5618 12621 5664
rect 12575 5512 12621 5558
rect 12575 5405 12621 5451
rect 12575 5298 12621 5344
rect 12799 6360 12845 6406
rect 12799 6254 12845 6300
rect 12799 6148 12845 6194
rect 12799 6042 12845 6088
rect 12799 5936 12845 5982
rect 12799 5830 12845 5876
rect 12799 5724 12845 5770
rect 12799 5618 12845 5664
rect 12799 5512 12845 5558
rect 12799 5405 12845 5451
rect 12799 5298 12845 5344
rect 13023 6360 13069 6406
rect 13023 6254 13069 6300
rect 13023 6148 13069 6194
rect 13023 6042 13069 6088
rect 13023 5936 13069 5982
rect 13023 5830 13069 5876
rect 13023 5724 13069 5770
rect 13023 5618 13069 5664
rect 13023 5512 13069 5558
rect 13023 5405 13069 5451
rect 13023 5298 13069 5344
rect 13247 6360 13293 6406
rect 13247 6254 13293 6300
rect 13247 6148 13293 6194
rect 13247 6042 13293 6088
rect 13247 5936 13293 5982
rect 13247 5830 13293 5876
rect 13247 5724 13293 5770
rect 13247 5618 13293 5664
rect 13247 5512 13293 5558
rect 13247 5405 13293 5451
rect 13247 5298 13293 5344
rect 13471 6360 13517 6406
rect 13471 6254 13517 6300
rect 13471 6148 13517 6194
rect 13471 6042 13517 6088
rect 13471 5936 13517 5982
rect 13471 5830 13517 5876
rect 13471 5724 13517 5770
rect 13471 5618 13517 5664
rect 13471 5512 13517 5558
rect 13471 5405 13517 5451
rect 13471 5298 13517 5344
rect 13695 6360 13741 6406
rect 13695 6254 13741 6300
rect 13695 6148 13741 6194
rect 13695 6042 13741 6088
rect 13695 5936 13741 5982
rect 13695 5830 13741 5876
rect 13695 5724 13741 5770
rect 13695 5618 13741 5664
rect 13695 5512 13741 5558
rect 13695 5405 13741 5451
rect 13695 5298 13741 5344
rect 7732 1124 7778 1170
rect 7732 989 7778 1035
rect 7732 854 7778 900
rect 7956 1124 8002 1170
rect 7956 989 8002 1035
rect 7956 854 8002 900
rect 8180 1124 8226 1170
rect 8180 989 8226 1035
rect 8180 854 8226 900
rect 8761 1077 8807 1123
rect 8761 873 8807 919
rect 9209 1077 9255 1123
rect 9209 873 9255 919
rect 9657 1077 9703 1123
rect 9657 873 9703 919
<< mvpsubdiff >>
rect 5188 29015 9138 29037
rect 12567 29015 16517 29037
rect 1753 28996 16517 29015
rect 1753 28950 1772 28996
rect 5202 28980 9132 28996
rect 12562 28980 16517 28996
rect 5202 28950 5401 28980
rect 1753 28934 5401 28950
rect 5447 28934 5559 28980
rect 5605 28934 5717 28980
rect 5763 28934 5875 28980
rect 5921 28934 6033 28980
rect 6079 28934 6191 28980
rect 6237 28934 6349 28980
rect 6395 28934 6507 28980
rect 6553 28934 6666 28980
rect 6712 28934 6824 28980
rect 6870 28934 6982 28980
rect 7028 28934 7140 28980
rect 7186 28934 7298 28980
rect 7344 28934 7456 28980
rect 7502 28934 7614 28980
rect 7660 28934 7773 28980
rect 7819 28934 7931 28980
rect 7977 28934 8089 28980
rect 8135 28934 8247 28980
rect 8293 28934 8405 28980
rect 8451 28934 8563 28980
rect 8609 28934 8721 28980
rect 8767 28934 8879 28980
rect 8925 28934 9037 28980
rect 12562 28950 12780 28980
rect 9083 28934 12780 28950
rect 12826 28934 12938 28980
rect 12984 28934 13096 28980
rect 13142 28934 13254 28980
rect 13300 28934 13412 28980
rect 13458 28934 13570 28980
rect 13616 28934 13728 28980
rect 13774 28934 13886 28980
rect 13932 28934 14045 28980
rect 14091 28934 14203 28980
rect 14249 28934 14361 28980
rect 14407 28934 14519 28980
rect 14565 28934 14677 28980
rect 14723 28934 14835 28980
rect 14881 28934 14993 28980
rect 15039 28934 15152 28980
rect 15198 28934 15310 28980
rect 15356 28934 15468 28980
rect 15514 28934 15626 28980
rect 15672 28934 15784 28980
rect 15830 28934 15942 28980
rect 15988 28934 16100 28980
rect 16146 28934 16258 28980
rect 16304 28934 16416 28980
rect 16462 28934 16517 28980
rect 1753 28931 16517 28934
rect 5188 28877 9138 28931
rect 12567 28877 16517 28931
rect 16581 28411 23118 28470
rect 16581 28365 16812 28411
rect 16858 28365 16970 28411
rect 17016 28365 17128 28411
rect 17174 28365 17286 28411
rect 17332 28365 17466 28411
rect 17512 28365 17624 28411
rect 17670 28365 17782 28411
rect 17828 28365 17940 28411
rect 17986 28365 18446 28411
rect 18492 28365 18604 28411
rect 18650 28365 18762 28411
rect 18808 28365 18920 28411
rect 18966 28365 19100 28411
rect 19146 28365 19258 28411
rect 19304 28365 19416 28411
rect 19462 28365 19574 28411
rect 19620 28365 20079 28411
rect 20125 28365 20237 28411
rect 20283 28365 20395 28411
rect 20441 28365 20553 28411
rect 20599 28365 20733 28411
rect 20779 28365 20891 28411
rect 20937 28365 21049 28411
rect 21095 28365 21207 28411
rect 21253 28365 21713 28411
rect 21759 28365 21871 28411
rect 21917 28365 22029 28411
rect 22075 28365 22187 28411
rect 22233 28365 22367 28411
rect 22413 28365 22525 28411
rect 22571 28365 22683 28411
rect 22729 28365 22841 28411
rect 22887 28365 23118 28411
rect 16581 28306 23118 28365
rect 23212 28407 24518 28426
rect 23212 28361 23231 28407
rect 24499 28361 24518 28407
rect 23212 28342 24518 28361
rect 24596 28411 28525 28470
rect 24596 28365 24726 28411
rect 24772 28365 24884 28411
rect 24930 28365 25042 28411
rect 25088 28365 25200 28411
rect 25246 28365 25358 28411
rect 25404 28365 25516 28411
rect 25562 28365 25674 28411
rect 25720 28365 25833 28411
rect 25879 28365 25991 28411
rect 26037 28365 26149 28411
rect 26195 28365 26307 28411
rect 26353 28365 26465 28411
rect 26511 28365 26623 28411
rect 26669 28365 26781 28411
rect 26827 28365 26939 28411
rect 26985 28365 27097 28411
rect 27143 28365 27256 28411
rect 27302 28365 27414 28411
rect 27460 28365 27572 28411
rect 27618 28365 27730 28411
rect 27776 28365 27888 28411
rect 27934 28365 28046 28411
rect 28092 28365 28204 28411
rect 28250 28365 28362 28411
rect 28408 28365 28525 28411
rect 24596 28305 28525 28365
rect 5731 26545 5890 26604
rect 5731 26499 5787 26545
rect 5833 26499 5890 26545
rect 5731 26382 5890 26499
rect 5731 26336 5787 26382
rect 5833 26336 5890 26382
rect 5731 26218 5890 26336
rect 5731 26172 5787 26218
rect 5833 26172 5890 26218
rect 5731 26055 5890 26172
rect 5731 26009 5787 26055
rect 5833 26009 5890 26055
rect 5731 25892 5890 26009
rect 5731 25846 5787 25892
rect 5833 25846 5890 25892
rect 5731 25728 5890 25846
rect 5731 25682 5787 25728
rect 5833 25682 5890 25728
rect 5731 25565 5890 25682
rect 5731 25519 5787 25565
rect 5833 25519 5890 25565
rect 5731 25460 5890 25519
rect 7422 26545 7581 26604
rect 7422 26499 7478 26545
rect 7524 26499 7581 26545
rect 7422 26382 7581 26499
rect 7422 26336 7478 26382
rect 7524 26336 7581 26382
rect 7422 26218 7581 26336
rect 7422 26172 7478 26218
rect 7524 26172 7581 26218
rect 7422 26055 7581 26172
rect 7422 26009 7478 26055
rect 7524 26009 7581 26055
rect 7422 25892 7581 26009
rect 7422 25846 7478 25892
rect 7524 25846 7581 25892
rect 7422 25728 7581 25846
rect 7422 25682 7478 25728
rect 7524 25682 7581 25728
rect 7422 25565 7581 25682
rect 7422 25519 7478 25565
rect 7524 25519 7581 25565
rect 7422 25460 7581 25519
rect 13110 26545 13269 26604
rect 13110 26499 13166 26545
rect 13212 26499 13269 26545
rect 13110 26382 13269 26499
rect 13110 26336 13166 26382
rect 13212 26336 13269 26382
rect 13110 26218 13269 26336
rect 13110 26172 13166 26218
rect 13212 26172 13269 26218
rect 13110 26055 13269 26172
rect 13110 26009 13166 26055
rect 13212 26009 13269 26055
rect 13110 25892 13269 26009
rect 13110 25846 13166 25892
rect 13212 25846 13269 25892
rect 13110 25728 13269 25846
rect 13110 25682 13166 25728
rect 13212 25682 13269 25728
rect 13110 25565 13269 25682
rect 13110 25519 13166 25565
rect 13212 25519 13269 25565
rect 13110 25460 13269 25519
rect 14801 26545 14960 26604
rect 14801 26499 14857 26545
rect 14903 26499 14960 26545
rect 14801 26382 14960 26499
rect 14801 26336 14857 26382
rect 14903 26336 14960 26382
rect 14801 26218 14960 26336
rect 14801 26172 14857 26218
rect 14903 26172 14960 26218
rect 14801 26055 14960 26172
rect 14801 26009 14857 26055
rect 14903 26009 14960 26055
rect 14801 25892 14960 26009
rect 14801 25846 14857 25892
rect 14903 25846 14960 25892
rect 14801 25728 14960 25846
rect 14801 25682 14857 25728
rect 14903 25682 14960 25728
rect 14801 25565 14960 25682
rect 14801 25519 14857 25565
rect 14903 25519 14960 25565
rect 14801 25460 14960 25519
rect 23596 26636 23755 26695
rect 23596 26590 23652 26636
rect 23698 26590 23755 26636
rect 23596 26473 23755 26590
rect 23596 26427 23652 26473
rect 23698 26427 23755 26473
rect 23596 26309 23755 26427
rect 23596 26263 23652 26309
rect 23698 26263 23755 26309
rect 23596 26146 23755 26263
rect 23596 26100 23652 26146
rect 23698 26100 23755 26146
rect 23596 25983 23755 26100
rect 23596 25937 23652 25983
rect 23698 25937 23755 25983
rect 23596 25819 23755 25937
rect 23596 25773 23652 25819
rect 23698 25773 23755 25819
rect 23596 25656 23755 25773
rect 23596 25610 23652 25656
rect 23698 25610 23755 25656
rect 23596 25551 23755 25610
rect 25286 26636 25445 26695
rect 25286 26590 25342 26636
rect 25388 26590 25445 26636
rect 25286 26473 25445 26590
rect 25286 26427 25342 26473
rect 25388 26427 25445 26473
rect 25286 26309 25445 26427
rect 25286 26263 25342 26309
rect 25388 26263 25445 26309
rect 25286 26146 25445 26263
rect 25286 26100 25342 26146
rect 25388 26100 25445 26146
rect 25286 25983 25445 26100
rect 25286 25937 25342 25983
rect 25388 25937 25445 25983
rect 25286 25819 25445 25937
rect 25286 25773 25342 25819
rect 25388 25773 25445 25819
rect 25286 25656 25445 25773
rect 25286 25610 25342 25656
rect 25388 25610 25445 25656
rect 25286 25551 25445 25610
rect 26977 26636 27136 26695
rect 26977 26590 27033 26636
rect 27079 26590 27136 26636
rect 26977 26473 27136 26590
rect 26977 26427 27033 26473
rect 27079 26427 27136 26473
rect 26977 26309 27136 26427
rect 26977 26263 27033 26309
rect 27079 26263 27136 26309
rect 26977 26146 27136 26263
rect 26977 26100 27033 26146
rect 27079 26100 27136 26146
rect 26977 25983 27136 26100
rect 26977 25937 27033 25983
rect 27079 25937 27136 25983
rect 26977 25819 27136 25937
rect 26977 25773 27033 25819
rect 27079 25773 27136 25819
rect 26977 25656 27136 25773
rect 26977 25610 27033 25656
rect 27079 25610 27136 25656
rect 26977 25551 27136 25610
rect 2512 20492 2644 20551
rect 2512 20446 2555 20492
rect 2601 20446 2644 20492
rect 2512 20329 2644 20446
rect 2512 20283 2555 20329
rect 2601 20283 2644 20329
rect 2512 20166 2644 20283
rect 2512 20120 2555 20166
rect 2601 20120 2644 20166
rect 2512 20003 2644 20120
rect 2512 19957 2555 20003
rect 2601 19957 2644 20003
rect 2512 19840 2644 19957
rect 2512 19794 2555 19840
rect 2601 19794 2644 19840
rect 2512 19676 2644 19794
rect 2512 19630 2555 19676
rect 2601 19630 2644 19676
rect 2512 19513 2644 19630
rect 2512 19467 2555 19513
rect 2601 19467 2644 19513
rect 2512 19350 2644 19467
rect 2512 19304 2555 19350
rect 2601 19304 2644 19350
rect 2512 19187 2644 19304
rect 2512 19141 2555 19187
rect 2601 19141 2644 19187
rect 2512 19023 2644 19141
rect 2512 18977 2555 19023
rect 2601 18977 2644 19023
rect 2512 18860 2644 18977
rect 2512 18814 2555 18860
rect 2601 18814 2644 18860
rect 2512 18697 2644 18814
rect 2512 18651 2555 18697
rect 2601 18651 2644 18697
rect 2512 18534 2644 18651
rect 2512 18488 2555 18534
rect 2601 18488 2644 18534
rect 2512 18371 2644 18488
rect 2512 18325 2555 18371
rect 2601 18325 2644 18371
rect 2512 18207 2644 18325
rect 2512 18161 2555 18207
rect 2601 18161 2644 18207
rect 2512 18101 2644 18161
rect 4304 20492 4436 20551
rect 4304 20446 4347 20492
rect 4393 20446 4436 20492
rect 4304 20329 4436 20446
rect 4304 20283 4347 20329
rect 4393 20283 4436 20329
rect 4304 20166 4436 20283
rect 4304 20120 4347 20166
rect 4393 20120 4436 20166
rect 4304 20003 4436 20120
rect 4304 19957 4347 20003
rect 4393 19957 4436 20003
rect 4304 19840 4436 19957
rect 4304 19794 4347 19840
rect 4393 19794 4436 19840
rect 4304 19676 4436 19794
rect 4304 19630 4347 19676
rect 4393 19630 4436 19676
rect 4304 19513 4436 19630
rect 4304 19467 4347 19513
rect 4393 19467 4436 19513
rect 4304 19350 4436 19467
rect 4304 19304 4347 19350
rect 4393 19304 4436 19350
rect 4304 19187 4436 19304
rect 4304 19141 4347 19187
rect 4393 19141 4436 19187
rect 4304 19023 4436 19141
rect 4304 18977 4347 19023
rect 4393 18977 4436 19023
rect 4304 18860 4436 18977
rect 4304 18814 4347 18860
rect 4393 18814 4436 18860
rect 4304 18697 4436 18814
rect 4304 18651 4347 18697
rect 4393 18651 4436 18697
rect 4304 18534 4436 18651
rect 4304 18488 4347 18534
rect 4393 18488 4436 18534
rect 4304 18371 4436 18488
rect 4304 18325 4347 18371
rect 4393 18325 4436 18371
rect 4304 18207 4436 18325
rect 4304 18161 4347 18207
rect 4393 18161 4436 18207
rect 4304 18101 4436 18161
rect 9891 20492 10023 20551
rect 9891 20446 9934 20492
rect 9980 20446 10023 20492
rect 9891 20329 10023 20446
rect 9891 20283 9934 20329
rect 9980 20283 10023 20329
rect 9891 20166 10023 20283
rect 9891 20120 9934 20166
rect 9980 20120 10023 20166
rect 9891 20003 10023 20120
rect 9891 19957 9934 20003
rect 9980 19957 10023 20003
rect 9891 19840 10023 19957
rect 9891 19794 9934 19840
rect 9980 19794 10023 19840
rect 9891 19676 10023 19794
rect 9891 19630 9934 19676
rect 9980 19630 10023 19676
rect 9891 19513 10023 19630
rect 9891 19467 9934 19513
rect 9980 19467 10023 19513
rect 9891 19350 10023 19467
rect 9891 19304 9934 19350
rect 9980 19304 10023 19350
rect 9891 19187 10023 19304
rect 9891 19141 9934 19187
rect 9980 19141 10023 19187
rect 9891 19023 10023 19141
rect 9891 18977 9934 19023
rect 9980 18977 10023 19023
rect 9891 18860 10023 18977
rect 9891 18814 9934 18860
rect 9980 18814 10023 18860
rect 9891 18697 10023 18814
rect 9891 18651 9934 18697
rect 9980 18651 10023 18697
rect 9891 18534 10023 18651
rect 9891 18488 9934 18534
rect 9980 18488 10023 18534
rect 9891 18371 10023 18488
rect 9891 18325 9934 18371
rect 9980 18325 10023 18371
rect 9891 18207 10023 18325
rect 9891 18161 9934 18207
rect 9980 18161 10023 18207
rect 9891 18101 10023 18161
rect 11683 20492 11815 20551
rect 11683 20446 11726 20492
rect 11772 20446 11815 20492
rect 11683 20329 11815 20446
rect 11683 20283 11726 20329
rect 11772 20283 11815 20329
rect 11683 20166 11815 20283
rect 11683 20120 11726 20166
rect 11772 20120 11815 20166
rect 11683 20003 11815 20120
rect 11683 19957 11726 20003
rect 11772 19957 11815 20003
rect 11683 19840 11815 19957
rect 11683 19794 11726 19840
rect 11772 19794 11815 19840
rect 11683 19676 11815 19794
rect 11683 19630 11726 19676
rect 11772 19630 11815 19676
rect 11683 19513 11815 19630
rect 11683 19467 11726 19513
rect 11772 19467 11815 19513
rect 11683 19350 11815 19467
rect 11683 19304 11726 19350
rect 11772 19304 11815 19350
rect 11683 19187 11815 19304
rect 11683 19141 11726 19187
rect 11772 19141 11815 19187
rect 11683 19023 11815 19141
rect 11683 18977 11726 19023
rect 11772 18977 11815 19023
rect 11683 18860 11815 18977
rect 11683 18814 11726 18860
rect 11772 18814 11815 18860
rect 11683 18697 11815 18814
rect 11683 18651 11726 18697
rect 11772 18651 11815 18697
rect 11683 18534 11815 18651
rect 11683 18488 11726 18534
rect 11772 18488 11815 18534
rect 11683 18371 11815 18488
rect 11683 18325 11726 18371
rect 11772 18325 11815 18371
rect 11683 18207 11815 18325
rect 11683 18161 11726 18207
rect 11772 18161 11815 18207
rect 11683 18101 11815 18161
rect 1681 17833 5267 17879
rect 1681 17787 1763 17833
rect 1809 17787 1921 17833
rect 1967 17787 2079 17833
rect 2125 17787 2237 17833
rect 2283 17787 2395 17833
rect 2441 17787 2715 17833
rect 2761 17787 2873 17833
rect 2919 17787 3031 17833
rect 3077 17787 3189 17833
rect 3235 17787 3347 17833
rect 3393 17787 3555 17833
rect 3601 17787 3713 17833
rect 3759 17787 3871 17833
rect 3917 17787 4029 17833
rect 4075 17787 4187 17833
rect 4233 17787 4507 17833
rect 4553 17787 4665 17833
rect 4711 17787 4823 17833
rect 4869 17787 4981 17833
rect 5027 17787 5139 17833
rect 5185 17787 5267 17833
rect 1681 17741 5267 17787
rect 9060 17833 12646 17879
rect 9060 17787 9142 17833
rect 9188 17787 9300 17833
rect 9346 17787 9458 17833
rect 9504 17787 9616 17833
rect 9662 17787 9774 17833
rect 9820 17787 10094 17833
rect 10140 17787 10252 17833
rect 10298 17787 10410 17833
rect 10456 17787 10568 17833
rect 10614 17787 10726 17833
rect 10772 17787 10934 17833
rect 10980 17787 11092 17833
rect 11138 17787 11250 17833
rect 11296 17787 11408 17833
rect 11454 17787 11566 17833
rect 11612 17787 11886 17833
rect 11932 17787 12044 17833
rect 12090 17787 12202 17833
rect 12248 17787 12360 17833
rect 12406 17787 12518 17833
rect 12564 17787 12646 17833
rect 9060 17741 12646 17787
rect 16581 17767 23118 17826
rect 16581 17721 16812 17767
rect 16858 17721 16970 17767
rect 17016 17721 17128 17767
rect 17174 17721 17286 17767
rect 17332 17721 17466 17767
rect 17512 17721 17624 17767
rect 17670 17721 17782 17767
rect 17828 17721 17940 17767
rect 17986 17721 18446 17767
rect 18492 17721 18604 17767
rect 18650 17721 18762 17767
rect 18808 17721 18920 17767
rect 18966 17721 19100 17767
rect 19146 17721 19258 17767
rect 19304 17721 19416 17767
rect 19462 17721 19574 17767
rect 19620 17721 20079 17767
rect 20125 17721 20237 17767
rect 20283 17721 20395 17767
rect 20441 17721 20553 17767
rect 20599 17721 20733 17767
rect 20779 17721 20891 17767
rect 20937 17721 21049 17767
rect 21095 17721 21207 17767
rect 21253 17721 21713 17767
rect 21759 17721 21871 17767
rect 21917 17721 22029 17767
rect 22075 17721 22187 17767
rect 22233 17721 22367 17767
rect 22413 17721 22525 17767
rect 22571 17721 22683 17767
rect 22729 17721 22841 17767
rect 22887 17721 23118 17767
rect 16581 17662 23118 17721
rect 2037 9669 19916 9729
rect 2037 9623 2443 9669
rect 2489 9623 2601 9669
rect 2647 9623 2759 9669
rect 2805 9623 2917 9669
rect 2963 9623 3075 9669
rect 3121 9623 3233 9669
rect 3279 9623 3392 9669
rect 3438 9623 3550 9669
rect 3596 9623 3708 9669
rect 3754 9623 3866 9669
rect 3912 9623 4024 9669
rect 4070 9623 4182 9669
rect 4228 9623 4340 9669
rect 4386 9623 4498 9669
rect 4544 9623 4656 9669
rect 4702 9623 4815 9669
rect 4861 9623 4973 9669
rect 5019 9623 5131 9669
rect 5177 9623 5289 9669
rect 5335 9623 5447 9669
rect 5493 9623 5605 9669
rect 5651 9623 5763 9669
rect 5809 9623 5921 9669
rect 5967 9623 6079 9669
rect 6125 9623 6238 9669
rect 6284 9623 6396 9669
rect 6442 9623 6554 9669
rect 6600 9623 6712 9669
rect 6758 9623 6870 9669
rect 6916 9623 7028 9669
rect 7074 9623 7186 9669
rect 7232 9623 7344 9669
rect 7390 9623 7502 9669
rect 7548 9623 7661 9669
rect 7707 9623 7819 9669
rect 7865 9623 7977 9669
rect 8023 9623 8135 9669
rect 8181 9623 8293 9669
rect 8339 9623 8451 9669
rect 8497 9623 8609 9669
rect 8655 9623 8767 9669
rect 8813 9623 8925 9669
rect 8971 9623 9084 9669
rect 9130 9623 9242 9669
rect 9288 9623 9400 9669
rect 9446 9623 9558 9669
rect 9604 9623 9716 9669
rect 9762 9623 9874 9669
rect 9920 9623 10032 9669
rect 10078 9623 10190 9669
rect 10236 9623 10348 9669
rect 10394 9623 10507 9669
rect 10553 9623 10665 9669
rect 10711 9623 10823 9669
rect 10869 9623 10981 9669
rect 11027 9623 11139 9669
rect 11185 9623 11297 9669
rect 11343 9623 11455 9669
rect 11501 9623 11613 9669
rect 11659 9623 11771 9669
rect 11817 9623 11930 9669
rect 11976 9623 12088 9669
rect 12134 9623 12246 9669
rect 12292 9623 12404 9669
rect 12450 9623 12562 9669
rect 12608 9623 12720 9669
rect 12766 9623 12878 9669
rect 12924 9623 13036 9669
rect 13082 9623 13195 9669
rect 13241 9623 13353 9669
rect 13399 9623 13511 9669
rect 13557 9623 13669 9669
rect 13715 9623 13827 9669
rect 13873 9623 13985 9669
rect 14031 9623 14143 9669
rect 14189 9623 14301 9669
rect 14347 9623 14459 9669
rect 14505 9623 14618 9669
rect 14664 9623 14776 9669
rect 14822 9623 14934 9669
rect 14980 9623 15092 9669
rect 15138 9623 15250 9669
rect 15296 9623 15408 9669
rect 15454 9623 15566 9669
rect 15612 9623 15724 9669
rect 15770 9623 15882 9669
rect 15928 9623 16041 9669
rect 16087 9623 16199 9669
rect 16245 9623 16357 9669
rect 16403 9623 16515 9669
rect 16561 9623 16673 9669
rect 16719 9623 16831 9669
rect 16877 9623 16989 9669
rect 17035 9623 17147 9669
rect 17193 9623 17305 9669
rect 17351 9623 17464 9669
rect 17510 9623 17622 9669
rect 17668 9623 17780 9669
rect 17826 9623 17938 9669
rect 17984 9623 18096 9669
rect 18142 9623 18254 9669
rect 18300 9623 18412 9669
rect 18458 9623 18570 9669
rect 18616 9623 18728 9669
rect 18774 9623 18887 9669
rect 18933 9623 19045 9669
rect 19091 9623 19203 9669
rect 19249 9623 19361 9669
rect 19407 9623 19519 9669
rect 19565 9623 19677 9669
rect 19723 9623 19835 9669
rect 19881 9623 19916 9669
rect 2037 9564 19916 9623
rect 7327 9343 13864 9402
rect 7327 9297 7558 9343
rect 7604 9297 7716 9343
rect 7762 9297 7874 9343
rect 7920 9297 8032 9343
rect 8078 9297 8212 9343
rect 8258 9297 8370 9343
rect 8416 9297 8528 9343
rect 8574 9297 8686 9343
rect 8732 9297 9191 9343
rect 9237 9297 9349 9343
rect 9395 9297 9507 9343
rect 9553 9297 9665 9343
rect 9711 9297 9845 9343
rect 9891 9297 10003 9343
rect 10049 9297 10161 9343
rect 10207 9297 10319 9343
rect 10365 9297 10825 9343
rect 10871 9297 10983 9343
rect 11029 9297 11141 9343
rect 11187 9297 11299 9343
rect 11345 9297 11479 9343
rect 11525 9297 11637 9343
rect 11683 9297 11795 9343
rect 11841 9297 11953 9343
rect 11999 9297 12459 9343
rect 12505 9297 12617 9343
rect 12663 9297 12775 9343
rect 12821 9297 12933 9343
rect 12979 9297 13113 9343
rect 13159 9297 13271 9343
rect 13317 9297 13429 9343
rect 13475 9297 13587 9343
rect 13633 9297 13864 9343
rect 7327 9238 13864 9297
rect 2261 9107 2420 9166
rect 2261 9061 2317 9107
rect 2363 9061 2420 9107
rect 2261 8944 2420 9061
rect 2261 8898 2317 8944
rect 2363 8898 2420 8944
rect 2261 8780 2420 8898
rect 2261 8734 2317 8780
rect 2363 8734 2420 8780
rect 2261 8617 2420 8734
rect 2261 8571 2317 8617
rect 2363 8571 2420 8617
rect 2261 8512 2420 8571
rect 3952 9107 4111 9166
rect 3952 9061 4008 9107
rect 4054 9061 4111 9107
rect 3952 8944 4111 9061
rect 3952 8898 4008 8944
rect 4054 8898 4111 8944
rect 3952 8780 4111 8898
rect 3952 8734 4008 8780
rect 4054 8734 4111 8780
rect 3952 8617 4111 8734
rect 3952 8571 4008 8617
rect 4054 8571 4111 8617
rect 3952 8512 4111 8571
rect 5643 9107 5802 9166
rect 5643 9061 5699 9107
rect 5745 9061 5802 9107
rect 5643 8944 5802 9061
rect 5643 8898 5699 8944
rect 5745 8898 5802 8944
rect 5643 8780 5802 8898
rect 5643 8734 5699 8780
rect 5745 8734 5802 8780
rect 5643 8617 5802 8734
rect 5643 8571 5699 8617
rect 5745 8571 5802 8617
rect 5643 8512 5802 8571
rect 7327 2274 13864 2334
rect 7327 2228 7558 2274
rect 7604 2228 7716 2274
rect 7762 2228 7874 2274
rect 7920 2228 8032 2274
rect 8078 2228 8212 2274
rect 8258 2228 8370 2274
rect 8416 2228 8528 2274
rect 8574 2228 8686 2274
rect 8732 2228 9191 2274
rect 9237 2228 9349 2274
rect 9395 2228 9507 2274
rect 9553 2228 9665 2274
rect 9711 2228 9845 2274
rect 9891 2228 10003 2274
rect 10049 2228 10161 2274
rect 10207 2228 10319 2274
rect 10365 2228 10825 2274
rect 10871 2228 10983 2274
rect 11029 2228 11141 2274
rect 11187 2228 11299 2274
rect 11345 2228 11479 2274
rect 11525 2228 11637 2274
rect 11683 2228 11795 2274
rect 11841 2228 11953 2274
rect 11999 2228 12459 2274
rect 12505 2228 12617 2274
rect 12663 2228 12775 2274
rect 12821 2228 12933 2274
rect 12979 2228 13113 2274
rect 13159 2228 13271 2274
rect 13317 2228 13429 2274
rect 13475 2228 13587 2274
rect 13633 2228 13864 2274
rect 7327 2169 13864 2228
rect 9903 1948 13699 2169
rect 9903 1902 9960 1948
rect 10006 1902 10118 1948
rect 10164 1902 10276 1948
rect 10322 1902 10434 1948
rect 10480 1902 10592 1948
rect 10638 1902 10750 1948
rect 10796 1902 10908 1948
rect 10954 1902 11066 1948
rect 11112 1902 11224 1948
rect 11270 1902 11383 1948
rect 11429 1902 11541 1948
rect 11587 1902 11699 1948
rect 11745 1902 11857 1948
rect 11903 1902 12015 1948
rect 12061 1902 12173 1948
rect 12219 1902 12332 1948
rect 12378 1902 12490 1948
rect 12536 1902 12648 1948
rect 12694 1902 12806 1948
rect 12852 1902 12964 1948
rect 13010 1902 13122 1948
rect 13168 1902 13280 1948
rect 13326 1902 13438 1948
rect 13484 1902 13596 1948
rect 13642 1902 13699 1948
rect 9903 1784 13699 1902
rect 9903 1738 9960 1784
rect 10006 1738 10118 1784
rect 10164 1738 10276 1784
rect 10322 1738 10434 1784
rect 10480 1738 10592 1784
rect 10638 1738 10750 1784
rect 10796 1738 10908 1784
rect 10954 1738 11066 1784
rect 11112 1738 11224 1784
rect 11270 1738 11383 1784
rect 11429 1738 11541 1784
rect 11587 1738 11699 1784
rect 11745 1738 11857 1784
rect 11903 1738 12015 1784
rect 12061 1738 12173 1784
rect 12219 1738 12332 1784
rect 12378 1738 12490 1784
rect 12536 1738 12648 1784
rect 12694 1738 12806 1784
rect 12852 1738 12964 1784
rect 13010 1738 13122 1784
rect 13168 1738 13280 1784
rect 13326 1738 13438 1784
rect 13484 1738 13596 1784
rect 13642 1738 13699 1784
rect 9903 1679 13699 1738
<< mvnsubdiff >>
rect 5630 27378 5714 27397
rect 5630 27144 5649 27378
rect 5695 27144 5714 27378
rect 5630 27125 5714 27144
rect 8122 27378 8206 27397
rect 8122 27144 8141 27378
rect 8187 27144 8206 27378
rect 8122 27125 8206 27144
rect 13009 27378 13093 27397
rect 13009 27144 13028 27378
rect 13074 27144 13093 27378
rect 13009 27125 13093 27144
rect 15501 27378 15585 27397
rect 15501 27144 15520 27378
rect 15566 27144 15585 27378
rect 15501 27125 15585 27144
rect 24959 27384 25043 27403
rect 24959 27244 24978 27384
rect 25024 27244 25043 27384
rect 24959 27225 25043 27244
rect 25989 27328 26073 27347
rect 25989 27188 26008 27328
rect 26054 27188 26073 27328
rect 25989 27169 26073 27188
rect 1536 24854 5826 24911
rect 1536 24808 1659 24854
rect 1705 24808 1818 24854
rect 1864 24808 2266 24854
rect 2312 24808 2424 24854
rect 2470 24808 2686 24854
rect 2732 24808 2844 24854
rect 2890 24808 3292 24854
rect 3338 24808 3451 24854
rect 3497 24808 3610 24854
rect 3656 24808 4058 24854
rect 4104 24808 4216 24854
rect 4262 24808 4478 24854
rect 4524 24808 4636 24854
rect 4682 24808 5084 24854
rect 5130 24808 5243 24854
rect 5289 24808 5726 24854
rect 5772 24808 5826 24854
rect 1536 24751 5826 24808
rect 5671 24690 5826 24751
rect 5671 24644 5726 24690
rect 5772 24644 5826 24690
rect 2536 21989 2620 22008
rect 2536 21661 2555 21989
rect 2601 21661 2620 21989
rect 2536 21642 2620 21661
rect 4328 21989 4412 22008
rect 4328 21661 4347 21989
rect 4393 21661 4412 21989
rect 4328 21642 4412 21661
rect 5671 24527 5826 24644
rect 5671 24481 5726 24527
rect 5772 24481 5826 24527
rect 5671 24364 5826 24481
rect 5671 24318 5726 24364
rect 5772 24318 5826 24364
rect 5671 24201 5826 24318
rect 5671 24155 5726 24201
rect 5772 24155 5826 24201
rect 5671 24037 5826 24155
rect 5671 23991 5726 24037
rect 5772 23991 5826 24037
rect 5671 23874 5826 23991
rect 5671 23828 5726 23874
rect 5772 23828 5826 23874
rect 5671 23711 5826 23828
rect 5671 23665 5726 23711
rect 5772 23665 5826 23711
rect 5671 23548 5826 23665
rect 5671 23502 5726 23548
rect 5772 23502 5826 23548
rect 5671 23384 5826 23502
rect 5671 23338 5726 23384
rect 5772 23338 5826 23384
rect 5671 23221 5826 23338
rect 5671 23175 5726 23221
rect 5772 23175 5826 23221
rect 5671 23058 5826 23175
rect 5671 23012 5726 23058
rect 5772 23012 5826 23058
rect 5671 22894 5826 23012
rect 5671 22848 5726 22894
rect 5772 22848 5826 22894
rect 5671 22731 5826 22848
rect 5671 22685 5726 22731
rect 5772 22685 5826 22731
rect 5671 22568 5826 22685
rect 5671 22522 5726 22568
rect 5772 22522 5826 22568
rect 5671 22405 5826 22522
rect 5671 22359 5726 22405
rect 5772 22359 5826 22405
rect 5671 22241 5826 22359
rect 5671 22195 5726 22241
rect 5772 22195 5826 22241
rect 5671 22078 5826 22195
rect 5671 22032 5726 22078
rect 5772 22032 5826 22078
rect 5671 21915 5826 22032
rect 5671 21869 5726 21915
rect 5772 21869 5826 21915
rect 5671 21752 5826 21869
rect 5671 21706 5726 21752
rect 5772 21706 5826 21752
rect 5671 21588 5826 21706
rect 5671 21542 5726 21588
rect 5772 21542 5826 21588
rect 5671 21486 5826 21542
rect 7362 24854 7517 24911
rect 7362 24808 7417 24854
rect 7463 24808 7517 24854
rect 7362 24690 7517 24808
rect 7362 24644 7417 24690
rect 7463 24644 7517 24690
rect 7362 24527 7517 24644
rect 7362 24481 7417 24527
rect 7463 24481 7517 24527
rect 7362 24364 7517 24481
rect 7362 24318 7417 24364
rect 7463 24318 7517 24364
rect 7362 24201 7517 24318
rect 7362 24155 7417 24201
rect 7463 24155 7517 24201
rect 7362 24037 7517 24155
rect 7362 23991 7417 24037
rect 7463 23991 7517 24037
rect 7362 23874 7517 23991
rect 7362 23828 7417 23874
rect 7463 23828 7517 23874
rect 7362 23711 7517 23828
rect 7362 23665 7417 23711
rect 7463 23665 7517 23711
rect 7362 23548 7517 23665
rect 7362 23502 7417 23548
rect 7463 23502 7517 23548
rect 7362 23384 7517 23502
rect 7362 23338 7417 23384
rect 7463 23338 7517 23384
rect 7362 23221 7517 23338
rect 7362 23175 7417 23221
rect 7463 23175 7517 23221
rect 7362 23058 7517 23175
rect 7362 23012 7417 23058
rect 7463 23012 7517 23058
rect 7362 22894 7517 23012
rect 7362 22848 7417 22894
rect 7463 22848 7517 22894
rect 7362 22731 7517 22848
rect 7362 22685 7417 22731
rect 7463 22685 7517 22731
rect 7362 22568 7517 22685
rect 7362 22522 7417 22568
rect 7463 22522 7517 22568
rect 7362 22405 7517 22522
rect 7362 22359 7417 22405
rect 7463 22359 7517 22405
rect 7362 22241 7517 22359
rect 7362 22195 7417 22241
rect 7463 22195 7517 22241
rect 7362 22078 7517 22195
rect 7362 22032 7417 22078
rect 7463 22032 7517 22078
rect 7362 21915 7517 22032
rect 7362 21869 7417 21915
rect 7463 21869 7517 21915
rect 7362 21752 7517 21869
rect 7362 21706 7417 21752
rect 7463 21706 7517 21752
rect 7362 21588 7517 21706
rect 7362 21542 7417 21588
rect 7463 21542 7517 21588
rect 7362 21486 7517 21542
rect 8915 24854 13205 24911
rect 8915 24808 9038 24854
rect 9084 24808 9197 24854
rect 9243 24808 9645 24854
rect 9691 24808 9803 24854
rect 9849 24808 10065 24854
rect 10111 24808 10223 24854
rect 10269 24808 10671 24854
rect 10717 24808 10830 24854
rect 10876 24808 10989 24854
rect 11035 24808 11437 24854
rect 11483 24808 11595 24854
rect 11641 24808 11857 24854
rect 11903 24808 12015 24854
rect 12061 24808 12463 24854
rect 12509 24808 12622 24854
rect 12668 24808 13105 24854
rect 13151 24808 13205 24854
rect 8915 24751 13205 24808
rect 13050 24690 13205 24751
rect 13050 24644 13105 24690
rect 13151 24644 13205 24690
rect 9915 21989 9999 22008
rect 9915 21661 9934 21989
rect 9980 21661 9999 21989
rect 9915 21642 9999 21661
rect 11707 21989 11791 22008
rect 11707 21661 11726 21989
rect 11772 21661 11791 21989
rect 11707 21642 11791 21661
rect 13050 24527 13205 24644
rect 13050 24481 13105 24527
rect 13151 24481 13205 24527
rect 13050 24364 13205 24481
rect 13050 24318 13105 24364
rect 13151 24318 13205 24364
rect 13050 24201 13205 24318
rect 13050 24155 13105 24201
rect 13151 24155 13205 24201
rect 13050 24037 13205 24155
rect 13050 23991 13105 24037
rect 13151 23991 13205 24037
rect 13050 23874 13205 23991
rect 13050 23828 13105 23874
rect 13151 23828 13205 23874
rect 13050 23711 13205 23828
rect 13050 23665 13105 23711
rect 13151 23665 13205 23711
rect 13050 23548 13205 23665
rect 13050 23502 13105 23548
rect 13151 23502 13205 23548
rect 13050 23384 13205 23502
rect 13050 23338 13105 23384
rect 13151 23338 13205 23384
rect 13050 23221 13205 23338
rect 13050 23175 13105 23221
rect 13151 23175 13205 23221
rect 13050 23058 13205 23175
rect 13050 23012 13105 23058
rect 13151 23012 13205 23058
rect 13050 22894 13205 23012
rect 13050 22848 13105 22894
rect 13151 22848 13205 22894
rect 13050 22731 13205 22848
rect 13050 22685 13105 22731
rect 13151 22685 13205 22731
rect 13050 22568 13205 22685
rect 13050 22522 13105 22568
rect 13151 22522 13205 22568
rect 13050 22405 13205 22522
rect 13050 22359 13105 22405
rect 13151 22359 13205 22405
rect 13050 22241 13205 22359
rect 13050 22195 13105 22241
rect 13151 22195 13205 22241
rect 13050 22078 13205 22195
rect 13050 22032 13105 22078
rect 13151 22032 13205 22078
rect 13050 21915 13205 22032
rect 13050 21869 13105 21915
rect 13151 21869 13205 21915
rect 13050 21752 13205 21869
rect 13050 21706 13105 21752
rect 13151 21706 13205 21752
rect 13050 21588 13205 21706
rect 13050 21542 13105 21588
rect 13151 21542 13205 21588
rect 13050 21486 13205 21542
rect 14741 24854 14896 24911
rect 14741 24808 14796 24854
rect 14842 24808 14896 24854
rect 14741 24690 14896 24808
rect 14741 24644 14796 24690
rect 14842 24644 14896 24690
rect 14741 24527 14896 24644
rect 14741 24481 14796 24527
rect 14842 24481 14896 24527
rect 14741 24364 14896 24481
rect 14741 24318 14796 24364
rect 14842 24318 14896 24364
rect 14741 24201 14896 24318
rect 14741 24155 14796 24201
rect 14842 24155 14896 24201
rect 14741 24037 14896 24155
rect 14741 23991 14796 24037
rect 14842 23991 14896 24037
rect 14741 23874 14896 23991
rect 14741 23828 14796 23874
rect 14842 23828 14896 23874
rect 14741 23711 14896 23828
rect 14741 23665 14796 23711
rect 14842 23665 14896 23711
rect 14741 23548 14896 23665
rect 14741 23502 14796 23548
rect 14842 23502 14896 23548
rect 14741 23384 14896 23502
rect 14741 23338 14796 23384
rect 14842 23338 14896 23384
rect 14741 23221 14896 23338
rect 14741 23175 14796 23221
rect 14842 23175 14896 23221
rect 14741 23058 14896 23175
rect 14741 23012 14796 23058
rect 14842 23012 14896 23058
rect 14741 22894 14896 23012
rect 14741 22848 14796 22894
rect 14842 22848 14896 22894
rect 14741 22731 14896 22848
rect 14741 22685 14796 22731
rect 14842 22685 14896 22731
rect 14741 22568 14896 22685
rect 14741 22522 14796 22568
rect 14842 22522 14896 22568
rect 14741 22405 14896 22522
rect 14741 22359 14796 22405
rect 14842 22359 14896 22405
rect 14741 22241 14896 22359
rect 14741 22195 14796 22241
rect 14842 22195 14896 22241
rect 14741 22078 14896 22195
rect 14741 22032 14796 22078
rect 14842 22032 14896 22078
rect 14741 21915 14896 22032
rect 14741 21869 14796 21915
rect 14842 21869 14896 21915
rect 14741 21752 14896 21869
rect 14741 21706 14796 21752
rect 14842 21706 14896 21752
rect 14741 21588 14896 21706
rect 14741 21542 14796 21588
rect 14842 21542 14896 21588
rect 14741 21486 14896 21542
rect 23537 24766 23691 24822
rect 23537 24720 23591 24766
rect 23637 24720 23691 24766
rect 23537 24602 23691 24720
rect 23537 24556 23591 24602
rect 23637 24556 23691 24602
rect 23537 24439 23691 24556
rect 23537 24393 23591 24439
rect 23637 24393 23691 24439
rect 16581 24290 23118 24346
rect 16581 24244 16981 24290
rect 17027 24244 17139 24290
rect 17185 24244 17297 24290
rect 17343 24244 17455 24290
rect 17501 24244 17613 24290
rect 17659 24244 17771 24290
rect 17817 24244 18615 24290
rect 18661 24244 18773 24290
rect 18819 24244 18931 24290
rect 18977 24244 19089 24290
rect 19135 24244 19247 24290
rect 19293 24244 19405 24290
rect 19451 24244 20248 24290
rect 20294 24244 20406 24290
rect 20452 24244 20564 24290
rect 20610 24244 20722 24290
rect 20768 24244 20880 24290
rect 20926 24244 21038 24290
rect 21084 24244 21882 24290
rect 21928 24244 22040 24290
rect 22086 24244 22198 24290
rect 22244 24244 22356 24290
rect 22402 24244 22514 24290
rect 22560 24244 22672 24290
rect 22718 24244 23118 24290
rect 16581 24186 23118 24244
rect 23537 24276 23691 24393
rect 23537 24230 23591 24276
rect 23637 24230 23691 24276
rect 23537 24113 23691 24230
rect 23537 24067 23591 24113
rect 23637 24067 23691 24113
rect 23537 23950 23691 24067
rect 23537 23904 23591 23950
rect 23637 23904 23691 23950
rect 23537 23786 23691 23904
rect 23537 23740 23591 23786
rect 23637 23740 23691 23786
rect 23537 23623 23691 23740
rect 23537 23577 23591 23623
rect 23637 23577 23691 23623
rect 23537 23460 23691 23577
rect 23537 23414 23591 23460
rect 23637 23414 23691 23460
rect 23537 23296 23691 23414
rect 23537 23250 23591 23296
rect 23637 23250 23691 23296
rect 23537 23133 23691 23250
rect 23537 23087 23591 23133
rect 23637 23087 23691 23133
rect 23537 22970 23691 23087
rect 23537 22924 23591 22970
rect 23637 22924 23691 22970
rect 23537 22806 23691 22924
rect 23537 22760 23591 22806
rect 23637 22760 23691 22806
rect 23537 22643 23691 22760
rect 23537 22597 23591 22643
rect 23637 22597 23691 22643
rect 23537 22480 23691 22597
rect 23537 22434 23591 22480
rect 23637 22434 23691 22480
rect 23537 22317 23691 22434
rect 23537 22271 23591 22317
rect 23637 22271 23691 22317
rect 23537 22154 23691 22271
rect 23537 22108 23591 22154
rect 23637 22108 23691 22154
rect 23537 21990 23691 22108
rect 23537 21944 23591 21990
rect 23637 21944 23691 21990
rect 23537 21887 23691 21944
rect 25227 24766 25381 24822
rect 25227 24720 25281 24766
rect 25327 24720 25381 24766
rect 25227 24602 25381 24720
rect 25227 24556 25281 24602
rect 25327 24556 25381 24602
rect 25227 24439 25381 24556
rect 25227 24393 25281 24439
rect 25327 24393 25381 24439
rect 25227 24276 25381 24393
rect 25227 24230 25281 24276
rect 25327 24230 25381 24276
rect 25227 24113 25381 24230
rect 25227 24067 25281 24113
rect 25327 24067 25381 24113
rect 25227 23950 25381 24067
rect 25227 23904 25281 23950
rect 25327 23904 25381 23950
rect 25227 23786 25381 23904
rect 25227 23740 25281 23786
rect 25327 23740 25381 23786
rect 25227 23623 25381 23740
rect 25227 23577 25281 23623
rect 25327 23577 25381 23623
rect 25227 23460 25381 23577
rect 25227 23414 25281 23460
rect 25327 23414 25381 23460
rect 25227 23296 25381 23414
rect 25227 23250 25281 23296
rect 25327 23250 25381 23296
rect 25227 23133 25381 23250
rect 25227 23087 25281 23133
rect 25327 23087 25381 23133
rect 25227 22970 25381 23087
rect 25227 22924 25281 22970
rect 25327 22924 25381 22970
rect 25227 22806 25381 22924
rect 25227 22760 25281 22806
rect 25327 22760 25381 22806
rect 25227 22643 25381 22760
rect 25227 22597 25281 22643
rect 25327 22597 25381 22643
rect 25227 22480 25381 22597
rect 25227 22434 25281 22480
rect 25327 22434 25381 22480
rect 25227 22317 25381 22434
rect 25227 22271 25281 22317
rect 25327 22271 25381 22317
rect 25227 22154 25381 22271
rect 25227 22108 25281 22154
rect 25327 22108 25381 22154
rect 25227 21990 25381 22108
rect 25227 21944 25281 21990
rect 25327 21944 25381 21990
rect 25227 21887 25381 21944
rect 26918 24766 27072 24822
rect 26918 24720 26972 24766
rect 27018 24720 27072 24766
rect 26918 24602 27072 24720
rect 26918 24556 26972 24602
rect 27018 24556 27072 24602
rect 26918 24439 27072 24556
rect 26918 24393 26972 24439
rect 27018 24393 27072 24439
rect 26918 24276 27072 24393
rect 26918 24230 26972 24276
rect 27018 24230 27072 24276
rect 26918 24113 27072 24230
rect 26918 24067 26972 24113
rect 27018 24067 27072 24113
rect 26918 23950 27072 24067
rect 26918 23904 26972 23950
rect 27018 23904 27072 23950
rect 26918 23786 27072 23904
rect 26918 23740 26972 23786
rect 27018 23740 27072 23786
rect 26918 23623 27072 23740
rect 26918 23577 26972 23623
rect 27018 23577 27072 23623
rect 26918 23460 27072 23577
rect 26918 23414 26972 23460
rect 27018 23414 27072 23460
rect 26918 23296 27072 23414
rect 26918 23250 26972 23296
rect 27018 23250 27072 23296
rect 26918 23133 27072 23250
rect 26918 23087 26972 23133
rect 27018 23087 27072 23133
rect 26918 22970 27072 23087
rect 26918 22924 26972 22970
rect 27018 22924 27072 22970
rect 26918 22806 27072 22924
rect 26918 22760 26972 22806
rect 27018 22760 27072 22806
rect 26918 22643 27072 22760
rect 26918 22597 26972 22643
rect 27018 22597 27072 22643
rect 26918 22480 27072 22597
rect 26918 22434 26972 22480
rect 27018 22434 27072 22480
rect 26918 22317 27072 22434
rect 26918 22271 26972 22317
rect 27018 22271 27072 22317
rect 26918 22154 27072 22271
rect 26918 22108 26972 22154
rect 27018 22108 27072 22154
rect 26918 21990 27072 22108
rect 26918 21944 26972 21990
rect 27018 21944 27072 21990
rect 26918 21887 27072 21944
rect 20114 16944 20180 16945
rect 1958 16887 20180 16944
rect 1958 16841 2012 16887
rect 2058 16841 2171 16887
rect 2217 16841 2329 16887
rect 2375 16841 2487 16887
rect 2533 16841 2645 16887
rect 2691 16841 2803 16887
rect 2849 16841 2961 16887
rect 3007 16841 3119 16887
rect 3165 16841 3277 16887
rect 3323 16841 3435 16887
rect 3481 16841 3594 16887
rect 3640 16841 3752 16887
rect 3798 16841 3910 16887
rect 3956 16841 4068 16887
rect 4114 16841 4226 16887
rect 4272 16841 4384 16887
rect 4430 16841 4542 16887
rect 4588 16841 4700 16887
rect 4746 16841 4858 16887
rect 4904 16841 5017 16887
rect 5063 16841 5175 16887
rect 5221 16841 5333 16887
rect 5379 16841 5491 16887
rect 5537 16841 5649 16887
rect 5695 16841 5807 16887
rect 5853 16841 5965 16887
rect 6011 16841 6123 16887
rect 6169 16841 6282 16887
rect 6328 16841 6440 16887
rect 6486 16841 6598 16887
rect 6644 16841 6756 16887
rect 6802 16841 6914 16887
rect 6960 16841 7072 16887
rect 7118 16841 7230 16887
rect 7276 16841 7388 16887
rect 7434 16841 7546 16887
rect 7592 16841 7705 16887
rect 7751 16841 7863 16887
rect 7909 16841 8021 16887
rect 8067 16841 8179 16887
rect 8225 16841 8337 16887
rect 8383 16841 8495 16887
rect 8541 16841 8653 16887
rect 8699 16841 8811 16887
rect 8857 16841 8969 16887
rect 9015 16841 9128 16887
rect 9174 16841 9286 16887
rect 9332 16841 9444 16887
rect 9490 16841 9602 16887
rect 9648 16841 9760 16887
rect 9806 16841 9918 16887
rect 9964 16841 10076 16887
rect 10122 16841 10234 16887
rect 10280 16841 10392 16887
rect 10438 16841 10551 16887
rect 10597 16841 10709 16887
rect 10755 16841 10867 16887
rect 10913 16841 11025 16887
rect 11071 16841 11183 16887
rect 11229 16841 11341 16887
rect 11387 16841 11499 16887
rect 11545 16841 11658 16887
rect 11704 16841 11816 16887
rect 11862 16841 11974 16887
rect 12020 16841 12132 16887
rect 12178 16841 12290 16887
rect 12336 16841 12448 16887
rect 12494 16841 12606 16887
rect 12652 16841 12764 16887
rect 12810 16841 12922 16887
rect 12968 16841 13081 16887
rect 13127 16841 13239 16887
rect 13285 16841 13397 16887
rect 13443 16841 13555 16887
rect 13601 16841 13713 16887
rect 13759 16841 13871 16887
rect 13917 16841 14029 16887
rect 14075 16841 14187 16887
rect 14233 16841 14345 16887
rect 14391 16841 14504 16887
rect 14550 16841 14662 16887
rect 14708 16841 14820 16887
rect 14866 16841 14978 16887
rect 15024 16841 15136 16887
rect 15182 16841 15294 16887
rect 15340 16841 15452 16887
rect 15498 16841 15610 16887
rect 15656 16841 15768 16887
rect 15814 16841 15927 16887
rect 15973 16841 16085 16887
rect 16131 16841 16243 16887
rect 16289 16841 16401 16887
rect 16447 16841 16559 16887
rect 16605 16841 16717 16887
rect 16763 16841 16875 16887
rect 16921 16841 17033 16887
rect 17079 16841 17192 16887
rect 17238 16841 17350 16887
rect 17396 16841 17508 16887
rect 17554 16841 17666 16887
rect 17712 16841 17824 16887
rect 17870 16841 17982 16887
rect 18028 16841 18140 16887
rect 18186 16841 18298 16887
rect 18344 16841 18456 16887
rect 18502 16841 18615 16887
rect 18661 16841 18773 16887
rect 18819 16841 18931 16887
rect 18977 16841 19089 16887
rect 19135 16841 19247 16887
rect 19293 16841 19405 16887
rect 19451 16841 19563 16887
rect 19609 16841 19721 16887
rect 19767 16841 19879 16887
rect 19925 16841 20038 16887
rect 20084 16841 20180 16887
rect 1958 16784 20180 16841
rect 2567 12263 2839 12282
rect 2567 12217 2586 12263
rect 2820 12217 2839 12263
rect 2567 12198 2839 12217
rect 3687 12263 3959 12282
rect 3687 12217 3706 12263
rect 3940 12217 3959 12263
rect 3687 12198 3959 12217
rect 4807 12263 5079 12282
rect 4807 12217 4826 12263
rect 5060 12217 5079 12263
rect 4807 12198 5079 12217
rect 5927 12263 6199 12282
rect 5927 12217 5946 12263
rect 6180 12217 6199 12263
rect 5927 12198 6199 12217
rect 7047 12263 7319 12282
rect 7047 12217 7066 12263
rect 7300 12217 7319 12263
rect 7047 12198 7319 12217
rect 8167 12263 8439 12282
rect 8167 12217 8186 12263
rect 8420 12217 8439 12263
rect 8167 12198 8439 12217
rect 9287 12263 9559 12282
rect 9287 12217 9306 12263
rect 9540 12217 9559 12263
rect 9287 12198 9559 12217
rect 10407 12263 10679 12282
rect 10407 12217 10426 12263
rect 10660 12217 10679 12263
rect 10407 12198 10679 12217
rect 11527 12263 11799 12282
rect 11527 12217 11546 12263
rect 11780 12217 11799 12263
rect 11527 12198 11799 12217
rect 12647 12263 12919 12282
rect 12647 12217 12666 12263
rect 12900 12217 12919 12263
rect 12647 12198 12919 12217
rect 13767 12263 14039 12282
rect 13767 12217 13786 12263
rect 14020 12217 14039 12263
rect 13767 12198 14039 12217
rect 14887 12263 15159 12282
rect 14887 12217 14906 12263
rect 15140 12217 15159 12263
rect 14887 12198 15159 12217
rect 16007 12263 16279 12282
rect 16007 12217 16026 12263
rect 16260 12217 16279 12263
rect 16007 12198 16279 12217
rect 17127 12263 17399 12282
rect 17127 12217 17146 12263
rect 17380 12217 17399 12263
rect 17127 12198 17399 12217
rect 18247 12263 18519 12282
rect 18247 12217 18266 12263
rect 18500 12217 18519 12263
rect 18247 12198 18519 12217
rect 19367 12263 19639 12282
rect 19367 12217 19386 12263
rect 19620 12217 19639 12263
rect 19367 12198 19639 12217
rect 2202 7894 2357 7951
rect 2202 7848 2256 7894
rect 2302 7848 2357 7894
rect 2202 7731 2357 7848
rect 2202 7685 2256 7731
rect 2302 7685 2357 7731
rect 2202 7568 2357 7685
rect 2202 7522 2256 7568
rect 2302 7522 2357 7568
rect 2202 7405 2357 7522
rect 2202 7359 2256 7405
rect 2302 7359 2357 7405
rect 2202 7242 2357 7359
rect 2202 7196 2256 7242
rect 2302 7196 2357 7242
rect 2202 7078 2357 7196
rect 2202 7032 2256 7078
rect 2302 7032 2357 7078
rect 2202 6915 2357 7032
rect 2202 6869 2256 6915
rect 2302 6869 2357 6915
rect 2202 6752 2357 6869
rect 2202 6706 2256 6752
rect 2302 6706 2357 6752
rect 2202 6588 2357 6706
rect 2202 6542 2256 6588
rect 2302 6542 2357 6588
rect 2202 6425 2357 6542
rect 2202 6379 2256 6425
rect 2302 6379 2357 6425
rect 2202 6262 2357 6379
rect 2202 6216 2256 6262
rect 2302 6216 2357 6262
rect 2202 6098 2357 6216
rect 2202 6052 2256 6098
rect 2302 6052 2357 6098
rect 2202 5935 2357 6052
rect 2202 5889 2256 5935
rect 2302 5889 2357 5935
rect 2202 5772 2357 5889
rect 2202 5726 2256 5772
rect 2302 5726 2357 5772
rect 2202 5609 2357 5726
rect 2202 5563 2256 5609
rect 2302 5563 2357 5609
rect 2202 5446 2357 5563
rect 2202 5400 2256 5446
rect 2302 5400 2357 5446
rect 2202 5342 2357 5400
rect 3893 7894 4048 7951
rect 3893 7848 3947 7894
rect 3993 7848 4048 7894
rect 3893 7731 4048 7848
rect 3893 7685 3947 7731
rect 3993 7685 4048 7731
rect 3893 7568 4048 7685
rect 3893 7522 3947 7568
rect 3993 7522 4048 7568
rect 3893 7405 4048 7522
rect 3893 7359 3947 7405
rect 3993 7359 4048 7405
rect 3893 7242 4048 7359
rect 3893 7196 3947 7242
rect 3993 7196 4048 7242
rect 3893 7078 4048 7196
rect 3893 7032 3947 7078
rect 3993 7032 4048 7078
rect 3893 6915 4048 7032
rect 3893 6869 3947 6915
rect 3993 6869 4048 6915
rect 3893 6752 4048 6869
rect 3893 6706 3947 6752
rect 3993 6706 4048 6752
rect 3893 6588 4048 6706
rect 3893 6542 3947 6588
rect 3993 6542 4048 6588
rect 3893 6425 4048 6542
rect 3893 6379 3947 6425
rect 3993 6379 4048 6425
rect 3893 6262 4048 6379
rect 3893 6216 3947 6262
rect 3993 6216 4048 6262
rect 3893 6098 4048 6216
rect 3893 6052 3947 6098
rect 3993 6052 4048 6098
rect 3893 5935 4048 6052
rect 3893 5889 3947 5935
rect 3993 5889 4048 5935
rect 3893 5772 4048 5889
rect 3893 5726 3947 5772
rect 3993 5726 4048 5772
rect 3893 5609 4048 5726
rect 3893 5563 3947 5609
rect 3993 5563 4048 5609
rect 3893 5446 4048 5563
rect 3893 5400 3947 5446
rect 3993 5400 4048 5446
rect 3893 5342 4048 5400
rect 5584 7894 5739 7951
rect 5584 7848 5638 7894
rect 5684 7848 5739 7894
rect 5584 7731 5739 7848
rect 5584 7685 5638 7731
rect 5684 7685 5739 7731
rect 5584 7568 5739 7685
rect 5584 7522 5638 7568
rect 5684 7522 5739 7568
rect 5584 7405 5739 7522
rect 5584 7359 5638 7405
rect 5684 7359 5739 7405
rect 5584 7242 5739 7359
rect 5584 7196 5638 7242
rect 5684 7196 5739 7242
rect 5584 7078 5739 7196
rect 5584 7032 5638 7078
rect 5684 7032 5739 7078
rect 5584 6915 5739 7032
rect 5584 6869 5638 6915
rect 5684 6869 5739 6915
rect 5584 6752 5739 6869
rect 5584 6706 5638 6752
rect 5684 6706 5739 6752
rect 5584 6588 5739 6706
rect 5584 6542 5638 6588
rect 5684 6542 5739 6588
rect 5584 6425 5739 6542
rect 5584 6379 5638 6425
rect 5684 6379 5739 6425
rect 5584 6262 5739 6379
rect 5584 6216 5638 6262
rect 5684 6216 5739 6262
rect 5584 6098 5739 6216
rect 5584 6052 5638 6098
rect 5684 6052 5739 6098
rect 5584 5935 5739 6052
rect 5584 5889 5638 5935
rect 5684 5889 5739 5935
rect 5584 5772 5739 5889
rect 5584 5726 5638 5772
rect 5684 5726 5739 5772
rect 5584 5609 5739 5726
rect 5584 5563 5638 5609
rect 5684 5563 5739 5609
rect 5584 5446 5739 5563
rect 5584 5400 5638 5446
rect 5684 5400 5739 5446
rect 5584 5342 5739 5400
rect 7327 6808 13864 6865
rect 7327 6762 7727 6808
rect 7773 6762 7885 6808
rect 7931 6762 8043 6808
rect 8089 6762 8201 6808
rect 8247 6762 8359 6808
rect 8405 6762 8517 6808
rect 8563 6762 9360 6808
rect 9406 6762 9518 6808
rect 9564 6762 9676 6808
rect 9722 6762 9834 6808
rect 9880 6762 9992 6808
rect 10038 6762 10150 6808
rect 10196 6762 10994 6808
rect 11040 6762 11152 6808
rect 11198 6762 11310 6808
rect 11356 6762 11468 6808
rect 11514 6762 11626 6808
rect 11672 6762 11784 6808
rect 11830 6762 12628 6808
rect 12674 6762 12786 6808
rect 12832 6762 12944 6808
rect 12990 6762 13102 6808
rect 13148 6762 13260 6808
rect 13306 6762 13418 6808
rect 13464 6762 13864 6808
rect 7327 6705 13864 6762
rect 9877 1107 13668 1164
rect 9877 1061 9931 1107
rect 9977 1061 10089 1107
rect 10135 1061 10247 1107
rect 10293 1061 10405 1107
rect 10451 1061 10563 1107
rect 10609 1061 10721 1107
rect 10767 1061 10879 1107
rect 10925 1061 11037 1107
rect 11083 1061 11195 1107
rect 11241 1061 11354 1107
rect 11400 1061 11512 1107
rect 11558 1061 11670 1107
rect 11716 1061 11828 1107
rect 11874 1061 11986 1107
rect 12032 1061 12144 1107
rect 12190 1061 12303 1107
rect 12349 1061 12461 1107
rect 12507 1061 12619 1107
rect 12665 1061 12777 1107
rect 12823 1061 12935 1107
rect 12981 1061 13093 1107
rect 13139 1061 13251 1107
rect 13297 1061 13409 1107
rect 13455 1061 13567 1107
rect 13613 1061 13668 1107
rect 9877 943 13668 1061
rect 9877 897 9931 943
rect 9977 897 10089 943
rect 10135 897 10247 943
rect 10293 897 10405 943
rect 10451 897 10563 943
rect 10609 897 10721 943
rect 10767 897 10879 943
rect 10925 897 11037 943
rect 11083 897 11195 943
rect 11241 897 11354 943
rect 11400 897 11512 943
rect 11558 897 11670 943
rect 11716 897 11828 943
rect 11874 897 11986 943
rect 12032 897 12144 943
rect 12190 897 12303 943
rect 12349 897 12461 943
rect 12507 897 12619 943
rect 12665 897 12777 943
rect 12823 897 12935 943
rect 12981 897 13093 943
rect 13139 897 13251 943
rect 13297 897 13409 943
rect 13455 897 13567 943
rect 13613 897 13668 943
rect 9877 840 13668 897
<< mvpsubdiffcont >>
rect 1772 28950 5202 28996
rect 9132 28980 12562 28996
rect 5401 28934 5447 28980
rect 5559 28934 5605 28980
rect 5717 28934 5763 28980
rect 5875 28934 5921 28980
rect 6033 28934 6079 28980
rect 6191 28934 6237 28980
rect 6349 28934 6395 28980
rect 6507 28934 6553 28980
rect 6666 28934 6712 28980
rect 6824 28934 6870 28980
rect 6982 28934 7028 28980
rect 7140 28934 7186 28980
rect 7298 28934 7344 28980
rect 7456 28934 7502 28980
rect 7614 28934 7660 28980
rect 7773 28934 7819 28980
rect 7931 28934 7977 28980
rect 8089 28934 8135 28980
rect 8247 28934 8293 28980
rect 8405 28934 8451 28980
rect 8563 28934 8609 28980
rect 8721 28934 8767 28980
rect 8879 28934 8925 28980
rect 9037 28950 12562 28980
rect 9037 28934 9083 28950
rect 12780 28934 12826 28980
rect 12938 28934 12984 28980
rect 13096 28934 13142 28980
rect 13254 28934 13300 28980
rect 13412 28934 13458 28980
rect 13570 28934 13616 28980
rect 13728 28934 13774 28980
rect 13886 28934 13932 28980
rect 14045 28934 14091 28980
rect 14203 28934 14249 28980
rect 14361 28934 14407 28980
rect 14519 28934 14565 28980
rect 14677 28934 14723 28980
rect 14835 28934 14881 28980
rect 14993 28934 15039 28980
rect 15152 28934 15198 28980
rect 15310 28934 15356 28980
rect 15468 28934 15514 28980
rect 15626 28934 15672 28980
rect 15784 28934 15830 28980
rect 15942 28934 15988 28980
rect 16100 28934 16146 28980
rect 16258 28934 16304 28980
rect 16416 28934 16462 28980
rect 16812 28365 16858 28411
rect 16970 28365 17016 28411
rect 17128 28365 17174 28411
rect 17286 28365 17332 28411
rect 17466 28365 17512 28411
rect 17624 28365 17670 28411
rect 17782 28365 17828 28411
rect 17940 28365 17986 28411
rect 18446 28365 18492 28411
rect 18604 28365 18650 28411
rect 18762 28365 18808 28411
rect 18920 28365 18966 28411
rect 19100 28365 19146 28411
rect 19258 28365 19304 28411
rect 19416 28365 19462 28411
rect 19574 28365 19620 28411
rect 20079 28365 20125 28411
rect 20237 28365 20283 28411
rect 20395 28365 20441 28411
rect 20553 28365 20599 28411
rect 20733 28365 20779 28411
rect 20891 28365 20937 28411
rect 21049 28365 21095 28411
rect 21207 28365 21253 28411
rect 21713 28365 21759 28411
rect 21871 28365 21917 28411
rect 22029 28365 22075 28411
rect 22187 28365 22233 28411
rect 22367 28365 22413 28411
rect 22525 28365 22571 28411
rect 22683 28365 22729 28411
rect 22841 28365 22887 28411
rect 23231 28361 24499 28407
rect 24726 28365 24772 28411
rect 24884 28365 24930 28411
rect 25042 28365 25088 28411
rect 25200 28365 25246 28411
rect 25358 28365 25404 28411
rect 25516 28365 25562 28411
rect 25674 28365 25720 28411
rect 25833 28365 25879 28411
rect 25991 28365 26037 28411
rect 26149 28365 26195 28411
rect 26307 28365 26353 28411
rect 26465 28365 26511 28411
rect 26623 28365 26669 28411
rect 26781 28365 26827 28411
rect 26939 28365 26985 28411
rect 27097 28365 27143 28411
rect 27256 28365 27302 28411
rect 27414 28365 27460 28411
rect 27572 28365 27618 28411
rect 27730 28365 27776 28411
rect 27888 28365 27934 28411
rect 28046 28365 28092 28411
rect 28204 28365 28250 28411
rect 28362 28365 28408 28411
rect 5787 26499 5833 26545
rect 5787 26336 5833 26382
rect 5787 26172 5833 26218
rect 5787 26009 5833 26055
rect 5787 25846 5833 25892
rect 5787 25682 5833 25728
rect 5787 25519 5833 25565
rect 7478 26499 7524 26545
rect 7478 26336 7524 26382
rect 7478 26172 7524 26218
rect 7478 26009 7524 26055
rect 7478 25846 7524 25892
rect 7478 25682 7524 25728
rect 7478 25519 7524 25565
rect 13166 26499 13212 26545
rect 13166 26336 13212 26382
rect 13166 26172 13212 26218
rect 13166 26009 13212 26055
rect 13166 25846 13212 25892
rect 13166 25682 13212 25728
rect 13166 25519 13212 25565
rect 14857 26499 14903 26545
rect 14857 26336 14903 26382
rect 14857 26172 14903 26218
rect 14857 26009 14903 26055
rect 14857 25846 14903 25892
rect 14857 25682 14903 25728
rect 14857 25519 14903 25565
rect 23652 26590 23698 26636
rect 23652 26427 23698 26473
rect 23652 26263 23698 26309
rect 23652 26100 23698 26146
rect 23652 25937 23698 25983
rect 23652 25773 23698 25819
rect 23652 25610 23698 25656
rect 25342 26590 25388 26636
rect 25342 26427 25388 26473
rect 25342 26263 25388 26309
rect 25342 26100 25388 26146
rect 25342 25937 25388 25983
rect 25342 25773 25388 25819
rect 25342 25610 25388 25656
rect 27033 26590 27079 26636
rect 27033 26427 27079 26473
rect 27033 26263 27079 26309
rect 27033 26100 27079 26146
rect 27033 25937 27079 25983
rect 27033 25773 27079 25819
rect 27033 25610 27079 25656
rect 2555 20446 2601 20492
rect 2555 20283 2601 20329
rect 2555 20120 2601 20166
rect 2555 19957 2601 20003
rect 2555 19794 2601 19840
rect 2555 19630 2601 19676
rect 2555 19467 2601 19513
rect 2555 19304 2601 19350
rect 2555 19141 2601 19187
rect 2555 18977 2601 19023
rect 2555 18814 2601 18860
rect 2555 18651 2601 18697
rect 2555 18488 2601 18534
rect 2555 18325 2601 18371
rect 2555 18161 2601 18207
rect 4347 20446 4393 20492
rect 4347 20283 4393 20329
rect 4347 20120 4393 20166
rect 4347 19957 4393 20003
rect 4347 19794 4393 19840
rect 4347 19630 4393 19676
rect 4347 19467 4393 19513
rect 4347 19304 4393 19350
rect 4347 19141 4393 19187
rect 4347 18977 4393 19023
rect 4347 18814 4393 18860
rect 4347 18651 4393 18697
rect 4347 18488 4393 18534
rect 4347 18325 4393 18371
rect 4347 18161 4393 18207
rect 9934 20446 9980 20492
rect 9934 20283 9980 20329
rect 9934 20120 9980 20166
rect 9934 19957 9980 20003
rect 9934 19794 9980 19840
rect 9934 19630 9980 19676
rect 9934 19467 9980 19513
rect 9934 19304 9980 19350
rect 9934 19141 9980 19187
rect 9934 18977 9980 19023
rect 9934 18814 9980 18860
rect 9934 18651 9980 18697
rect 9934 18488 9980 18534
rect 9934 18325 9980 18371
rect 9934 18161 9980 18207
rect 11726 20446 11772 20492
rect 11726 20283 11772 20329
rect 11726 20120 11772 20166
rect 11726 19957 11772 20003
rect 11726 19794 11772 19840
rect 11726 19630 11772 19676
rect 11726 19467 11772 19513
rect 11726 19304 11772 19350
rect 11726 19141 11772 19187
rect 11726 18977 11772 19023
rect 11726 18814 11772 18860
rect 11726 18651 11772 18697
rect 11726 18488 11772 18534
rect 11726 18325 11772 18371
rect 11726 18161 11772 18207
rect 1763 17787 1809 17833
rect 1921 17787 1967 17833
rect 2079 17787 2125 17833
rect 2237 17787 2283 17833
rect 2395 17787 2441 17833
rect 2715 17787 2761 17833
rect 2873 17787 2919 17833
rect 3031 17787 3077 17833
rect 3189 17787 3235 17833
rect 3347 17787 3393 17833
rect 3555 17787 3601 17833
rect 3713 17787 3759 17833
rect 3871 17787 3917 17833
rect 4029 17787 4075 17833
rect 4187 17787 4233 17833
rect 4507 17787 4553 17833
rect 4665 17787 4711 17833
rect 4823 17787 4869 17833
rect 4981 17787 5027 17833
rect 5139 17787 5185 17833
rect 9142 17787 9188 17833
rect 9300 17787 9346 17833
rect 9458 17787 9504 17833
rect 9616 17787 9662 17833
rect 9774 17787 9820 17833
rect 10094 17787 10140 17833
rect 10252 17787 10298 17833
rect 10410 17787 10456 17833
rect 10568 17787 10614 17833
rect 10726 17787 10772 17833
rect 10934 17787 10980 17833
rect 11092 17787 11138 17833
rect 11250 17787 11296 17833
rect 11408 17787 11454 17833
rect 11566 17787 11612 17833
rect 11886 17787 11932 17833
rect 12044 17787 12090 17833
rect 12202 17787 12248 17833
rect 12360 17787 12406 17833
rect 12518 17787 12564 17833
rect 16812 17721 16858 17767
rect 16970 17721 17016 17767
rect 17128 17721 17174 17767
rect 17286 17721 17332 17767
rect 17466 17721 17512 17767
rect 17624 17721 17670 17767
rect 17782 17721 17828 17767
rect 17940 17721 17986 17767
rect 18446 17721 18492 17767
rect 18604 17721 18650 17767
rect 18762 17721 18808 17767
rect 18920 17721 18966 17767
rect 19100 17721 19146 17767
rect 19258 17721 19304 17767
rect 19416 17721 19462 17767
rect 19574 17721 19620 17767
rect 20079 17721 20125 17767
rect 20237 17721 20283 17767
rect 20395 17721 20441 17767
rect 20553 17721 20599 17767
rect 20733 17721 20779 17767
rect 20891 17721 20937 17767
rect 21049 17721 21095 17767
rect 21207 17721 21253 17767
rect 21713 17721 21759 17767
rect 21871 17721 21917 17767
rect 22029 17721 22075 17767
rect 22187 17721 22233 17767
rect 22367 17721 22413 17767
rect 22525 17721 22571 17767
rect 22683 17721 22729 17767
rect 22841 17721 22887 17767
rect 2443 9623 2489 9669
rect 2601 9623 2647 9669
rect 2759 9623 2805 9669
rect 2917 9623 2963 9669
rect 3075 9623 3121 9669
rect 3233 9623 3279 9669
rect 3392 9623 3438 9669
rect 3550 9623 3596 9669
rect 3708 9623 3754 9669
rect 3866 9623 3912 9669
rect 4024 9623 4070 9669
rect 4182 9623 4228 9669
rect 4340 9623 4386 9669
rect 4498 9623 4544 9669
rect 4656 9623 4702 9669
rect 4815 9623 4861 9669
rect 4973 9623 5019 9669
rect 5131 9623 5177 9669
rect 5289 9623 5335 9669
rect 5447 9623 5493 9669
rect 5605 9623 5651 9669
rect 5763 9623 5809 9669
rect 5921 9623 5967 9669
rect 6079 9623 6125 9669
rect 6238 9623 6284 9669
rect 6396 9623 6442 9669
rect 6554 9623 6600 9669
rect 6712 9623 6758 9669
rect 6870 9623 6916 9669
rect 7028 9623 7074 9669
rect 7186 9623 7232 9669
rect 7344 9623 7390 9669
rect 7502 9623 7548 9669
rect 7661 9623 7707 9669
rect 7819 9623 7865 9669
rect 7977 9623 8023 9669
rect 8135 9623 8181 9669
rect 8293 9623 8339 9669
rect 8451 9623 8497 9669
rect 8609 9623 8655 9669
rect 8767 9623 8813 9669
rect 8925 9623 8971 9669
rect 9084 9623 9130 9669
rect 9242 9623 9288 9669
rect 9400 9623 9446 9669
rect 9558 9623 9604 9669
rect 9716 9623 9762 9669
rect 9874 9623 9920 9669
rect 10032 9623 10078 9669
rect 10190 9623 10236 9669
rect 10348 9623 10394 9669
rect 10507 9623 10553 9669
rect 10665 9623 10711 9669
rect 10823 9623 10869 9669
rect 10981 9623 11027 9669
rect 11139 9623 11185 9669
rect 11297 9623 11343 9669
rect 11455 9623 11501 9669
rect 11613 9623 11659 9669
rect 11771 9623 11817 9669
rect 11930 9623 11976 9669
rect 12088 9623 12134 9669
rect 12246 9623 12292 9669
rect 12404 9623 12450 9669
rect 12562 9623 12608 9669
rect 12720 9623 12766 9669
rect 12878 9623 12924 9669
rect 13036 9623 13082 9669
rect 13195 9623 13241 9669
rect 13353 9623 13399 9669
rect 13511 9623 13557 9669
rect 13669 9623 13715 9669
rect 13827 9623 13873 9669
rect 13985 9623 14031 9669
rect 14143 9623 14189 9669
rect 14301 9623 14347 9669
rect 14459 9623 14505 9669
rect 14618 9623 14664 9669
rect 14776 9623 14822 9669
rect 14934 9623 14980 9669
rect 15092 9623 15138 9669
rect 15250 9623 15296 9669
rect 15408 9623 15454 9669
rect 15566 9623 15612 9669
rect 15724 9623 15770 9669
rect 15882 9623 15928 9669
rect 16041 9623 16087 9669
rect 16199 9623 16245 9669
rect 16357 9623 16403 9669
rect 16515 9623 16561 9669
rect 16673 9623 16719 9669
rect 16831 9623 16877 9669
rect 16989 9623 17035 9669
rect 17147 9623 17193 9669
rect 17305 9623 17351 9669
rect 17464 9623 17510 9669
rect 17622 9623 17668 9669
rect 17780 9623 17826 9669
rect 17938 9623 17984 9669
rect 18096 9623 18142 9669
rect 18254 9623 18300 9669
rect 18412 9623 18458 9669
rect 18570 9623 18616 9669
rect 18728 9623 18774 9669
rect 18887 9623 18933 9669
rect 19045 9623 19091 9669
rect 19203 9623 19249 9669
rect 19361 9623 19407 9669
rect 19519 9623 19565 9669
rect 19677 9623 19723 9669
rect 19835 9623 19881 9669
rect 7558 9297 7604 9343
rect 7716 9297 7762 9343
rect 7874 9297 7920 9343
rect 8032 9297 8078 9343
rect 8212 9297 8258 9343
rect 8370 9297 8416 9343
rect 8528 9297 8574 9343
rect 8686 9297 8732 9343
rect 9191 9297 9237 9343
rect 9349 9297 9395 9343
rect 9507 9297 9553 9343
rect 9665 9297 9711 9343
rect 9845 9297 9891 9343
rect 10003 9297 10049 9343
rect 10161 9297 10207 9343
rect 10319 9297 10365 9343
rect 10825 9297 10871 9343
rect 10983 9297 11029 9343
rect 11141 9297 11187 9343
rect 11299 9297 11345 9343
rect 11479 9297 11525 9343
rect 11637 9297 11683 9343
rect 11795 9297 11841 9343
rect 11953 9297 11999 9343
rect 12459 9297 12505 9343
rect 12617 9297 12663 9343
rect 12775 9297 12821 9343
rect 12933 9297 12979 9343
rect 13113 9297 13159 9343
rect 13271 9297 13317 9343
rect 13429 9297 13475 9343
rect 13587 9297 13633 9343
rect 2317 9061 2363 9107
rect 2317 8898 2363 8944
rect 2317 8734 2363 8780
rect 2317 8571 2363 8617
rect 4008 9061 4054 9107
rect 4008 8898 4054 8944
rect 4008 8734 4054 8780
rect 4008 8571 4054 8617
rect 5699 9061 5745 9107
rect 5699 8898 5745 8944
rect 5699 8734 5745 8780
rect 5699 8571 5745 8617
rect 7558 2228 7604 2274
rect 7716 2228 7762 2274
rect 7874 2228 7920 2274
rect 8032 2228 8078 2274
rect 8212 2228 8258 2274
rect 8370 2228 8416 2274
rect 8528 2228 8574 2274
rect 8686 2228 8732 2274
rect 9191 2228 9237 2274
rect 9349 2228 9395 2274
rect 9507 2228 9553 2274
rect 9665 2228 9711 2274
rect 9845 2228 9891 2274
rect 10003 2228 10049 2274
rect 10161 2228 10207 2274
rect 10319 2228 10365 2274
rect 10825 2228 10871 2274
rect 10983 2228 11029 2274
rect 11141 2228 11187 2274
rect 11299 2228 11345 2274
rect 11479 2228 11525 2274
rect 11637 2228 11683 2274
rect 11795 2228 11841 2274
rect 11953 2228 11999 2274
rect 12459 2228 12505 2274
rect 12617 2228 12663 2274
rect 12775 2228 12821 2274
rect 12933 2228 12979 2274
rect 13113 2228 13159 2274
rect 13271 2228 13317 2274
rect 13429 2228 13475 2274
rect 13587 2228 13633 2274
rect 9960 1902 10006 1948
rect 10118 1902 10164 1948
rect 10276 1902 10322 1948
rect 10434 1902 10480 1948
rect 10592 1902 10638 1948
rect 10750 1902 10796 1948
rect 10908 1902 10954 1948
rect 11066 1902 11112 1948
rect 11224 1902 11270 1948
rect 11383 1902 11429 1948
rect 11541 1902 11587 1948
rect 11699 1902 11745 1948
rect 11857 1902 11903 1948
rect 12015 1902 12061 1948
rect 12173 1902 12219 1948
rect 12332 1902 12378 1948
rect 12490 1902 12536 1948
rect 12648 1902 12694 1948
rect 12806 1902 12852 1948
rect 12964 1902 13010 1948
rect 13122 1902 13168 1948
rect 13280 1902 13326 1948
rect 13438 1902 13484 1948
rect 13596 1902 13642 1948
rect 9960 1738 10006 1784
rect 10118 1738 10164 1784
rect 10276 1738 10322 1784
rect 10434 1738 10480 1784
rect 10592 1738 10638 1784
rect 10750 1738 10796 1784
rect 10908 1738 10954 1784
rect 11066 1738 11112 1784
rect 11224 1738 11270 1784
rect 11383 1738 11429 1784
rect 11541 1738 11587 1784
rect 11699 1738 11745 1784
rect 11857 1738 11903 1784
rect 12015 1738 12061 1784
rect 12173 1738 12219 1784
rect 12332 1738 12378 1784
rect 12490 1738 12536 1784
rect 12648 1738 12694 1784
rect 12806 1738 12852 1784
rect 12964 1738 13010 1784
rect 13122 1738 13168 1784
rect 13280 1738 13326 1784
rect 13438 1738 13484 1784
rect 13596 1738 13642 1784
<< mvnsubdiffcont >>
rect 5649 27144 5695 27378
rect 8141 27144 8187 27378
rect 13028 27144 13074 27378
rect 15520 27144 15566 27378
rect 24978 27244 25024 27384
rect 26008 27188 26054 27328
rect 1659 24808 1705 24854
rect 1818 24808 1864 24854
rect 2266 24808 2312 24854
rect 2424 24808 2470 24854
rect 2686 24808 2732 24854
rect 2844 24808 2890 24854
rect 3292 24808 3338 24854
rect 3451 24808 3497 24854
rect 3610 24808 3656 24854
rect 4058 24808 4104 24854
rect 4216 24808 4262 24854
rect 4478 24808 4524 24854
rect 4636 24808 4682 24854
rect 5084 24808 5130 24854
rect 5243 24808 5289 24854
rect 5726 24808 5772 24854
rect 5726 24644 5772 24690
rect 2555 21661 2601 21989
rect 4347 21661 4393 21989
rect 5726 24481 5772 24527
rect 5726 24318 5772 24364
rect 5726 24155 5772 24201
rect 5726 23991 5772 24037
rect 5726 23828 5772 23874
rect 5726 23665 5772 23711
rect 5726 23502 5772 23548
rect 5726 23338 5772 23384
rect 5726 23175 5772 23221
rect 5726 23012 5772 23058
rect 5726 22848 5772 22894
rect 5726 22685 5772 22731
rect 5726 22522 5772 22568
rect 5726 22359 5772 22405
rect 5726 22195 5772 22241
rect 5726 22032 5772 22078
rect 5726 21869 5772 21915
rect 5726 21706 5772 21752
rect 5726 21542 5772 21588
rect 7417 24808 7463 24854
rect 7417 24644 7463 24690
rect 7417 24481 7463 24527
rect 7417 24318 7463 24364
rect 7417 24155 7463 24201
rect 7417 23991 7463 24037
rect 7417 23828 7463 23874
rect 7417 23665 7463 23711
rect 7417 23502 7463 23548
rect 7417 23338 7463 23384
rect 7417 23175 7463 23221
rect 7417 23012 7463 23058
rect 7417 22848 7463 22894
rect 7417 22685 7463 22731
rect 7417 22522 7463 22568
rect 7417 22359 7463 22405
rect 7417 22195 7463 22241
rect 7417 22032 7463 22078
rect 7417 21869 7463 21915
rect 7417 21706 7463 21752
rect 7417 21542 7463 21588
rect 9038 24808 9084 24854
rect 9197 24808 9243 24854
rect 9645 24808 9691 24854
rect 9803 24808 9849 24854
rect 10065 24808 10111 24854
rect 10223 24808 10269 24854
rect 10671 24808 10717 24854
rect 10830 24808 10876 24854
rect 10989 24808 11035 24854
rect 11437 24808 11483 24854
rect 11595 24808 11641 24854
rect 11857 24808 11903 24854
rect 12015 24808 12061 24854
rect 12463 24808 12509 24854
rect 12622 24808 12668 24854
rect 13105 24808 13151 24854
rect 13105 24644 13151 24690
rect 9934 21661 9980 21989
rect 11726 21661 11772 21989
rect 13105 24481 13151 24527
rect 13105 24318 13151 24364
rect 13105 24155 13151 24201
rect 13105 23991 13151 24037
rect 13105 23828 13151 23874
rect 13105 23665 13151 23711
rect 13105 23502 13151 23548
rect 13105 23338 13151 23384
rect 13105 23175 13151 23221
rect 13105 23012 13151 23058
rect 13105 22848 13151 22894
rect 13105 22685 13151 22731
rect 13105 22522 13151 22568
rect 13105 22359 13151 22405
rect 13105 22195 13151 22241
rect 13105 22032 13151 22078
rect 13105 21869 13151 21915
rect 13105 21706 13151 21752
rect 13105 21542 13151 21588
rect 14796 24808 14842 24854
rect 14796 24644 14842 24690
rect 14796 24481 14842 24527
rect 14796 24318 14842 24364
rect 14796 24155 14842 24201
rect 14796 23991 14842 24037
rect 14796 23828 14842 23874
rect 14796 23665 14842 23711
rect 14796 23502 14842 23548
rect 14796 23338 14842 23384
rect 14796 23175 14842 23221
rect 14796 23012 14842 23058
rect 14796 22848 14842 22894
rect 14796 22685 14842 22731
rect 14796 22522 14842 22568
rect 14796 22359 14842 22405
rect 14796 22195 14842 22241
rect 14796 22032 14842 22078
rect 14796 21869 14842 21915
rect 14796 21706 14842 21752
rect 14796 21542 14842 21588
rect 23591 24720 23637 24766
rect 23591 24556 23637 24602
rect 23591 24393 23637 24439
rect 16981 24244 17027 24290
rect 17139 24244 17185 24290
rect 17297 24244 17343 24290
rect 17455 24244 17501 24290
rect 17613 24244 17659 24290
rect 17771 24244 17817 24290
rect 18615 24244 18661 24290
rect 18773 24244 18819 24290
rect 18931 24244 18977 24290
rect 19089 24244 19135 24290
rect 19247 24244 19293 24290
rect 19405 24244 19451 24290
rect 20248 24244 20294 24290
rect 20406 24244 20452 24290
rect 20564 24244 20610 24290
rect 20722 24244 20768 24290
rect 20880 24244 20926 24290
rect 21038 24244 21084 24290
rect 21882 24244 21928 24290
rect 22040 24244 22086 24290
rect 22198 24244 22244 24290
rect 22356 24244 22402 24290
rect 22514 24244 22560 24290
rect 22672 24244 22718 24290
rect 23591 24230 23637 24276
rect 23591 24067 23637 24113
rect 23591 23904 23637 23950
rect 23591 23740 23637 23786
rect 23591 23577 23637 23623
rect 23591 23414 23637 23460
rect 23591 23250 23637 23296
rect 23591 23087 23637 23133
rect 23591 22924 23637 22970
rect 23591 22760 23637 22806
rect 23591 22597 23637 22643
rect 23591 22434 23637 22480
rect 23591 22271 23637 22317
rect 23591 22108 23637 22154
rect 23591 21944 23637 21990
rect 25281 24720 25327 24766
rect 25281 24556 25327 24602
rect 25281 24393 25327 24439
rect 25281 24230 25327 24276
rect 25281 24067 25327 24113
rect 25281 23904 25327 23950
rect 25281 23740 25327 23786
rect 25281 23577 25327 23623
rect 25281 23414 25327 23460
rect 25281 23250 25327 23296
rect 25281 23087 25327 23133
rect 25281 22924 25327 22970
rect 25281 22760 25327 22806
rect 25281 22597 25327 22643
rect 25281 22434 25327 22480
rect 25281 22271 25327 22317
rect 25281 22108 25327 22154
rect 25281 21944 25327 21990
rect 26972 24720 27018 24766
rect 26972 24556 27018 24602
rect 26972 24393 27018 24439
rect 26972 24230 27018 24276
rect 26972 24067 27018 24113
rect 26972 23904 27018 23950
rect 26972 23740 27018 23786
rect 26972 23577 27018 23623
rect 26972 23414 27018 23460
rect 26972 23250 27018 23296
rect 26972 23087 27018 23133
rect 26972 22924 27018 22970
rect 26972 22760 27018 22806
rect 26972 22597 27018 22643
rect 26972 22434 27018 22480
rect 26972 22271 27018 22317
rect 26972 22108 27018 22154
rect 26972 21944 27018 21990
rect 2012 16841 2058 16887
rect 2171 16841 2217 16887
rect 2329 16841 2375 16887
rect 2487 16841 2533 16887
rect 2645 16841 2691 16887
rect 2803 16841 2849 16887
rect 2961 16841 3007 16887
rect 3119 16841 3165 16887
rect 3277 16841 3323 16887
rect 3435 16841 3481 16887
rect 3594 16841 3640 16887
rect 3752 16841 3798 16887
rect 3910 16841 3956 16887
rect 4068 16841 4114 16887
rect 4226 16841 4272 16887
rect 4384 16841 4430 16887
rect 4542 16841 4588 16887
rect 4700 16841 4746 16887
rect 4858 16841 4904 16887
rect 5017 16841 5063 16887
rect 5175 16841 5221 16887
rect 5333 16841 5379 16887
rect 5491 16841 5537 16887
rect 5649 16841 5695 16887
rect 5807 16841 5853 16887
rect 5965 16841 6011 16887
rect 6123 16841 6169 16887
rect 6282 16841 6328 16887
rect 6440 16841 6486 16887
rect 6598 16841 6644 16887
rect 6756 16841 6802 16887
rect 6914 16841 6960 16887
rect 7072 16841 7118 16887
rect 7230 16841 7276 16887
rect 7388 16841 7434 16887
rect 7546 16841 7592 16887
rect 7705 16841 7751 16887
rect 7863 16841 7909 16887
rect 8021 16841 8067 16887
rect 8179 16841 8225 16887
rect 8337 16841 8383 16887
rect 8495 16841 8541 16887
rect 8653 16841 8699 16887
rect 8811 16841 8857 16887
rect 8969 16841 9015 16887
rect 9128 16841 9174 16887
rect 9286 16841 9332 16887
rect 9444 16841 9490 16887
rect 9602 16841 9648 16887
rect 9760 16841 9806 16887
rect 9918 16841 9964 16887
rect 10076 16841 10122 16887
rect 10234 16841 10280 16887
rect 10392 16841 10438 16887
rect 10551 16841 10597 16887
rect 10709 16841 10755 16887
rect 10867 16841 10913 16887
rect 11025 16841 11071 16887
rect 11183 16841 11229 16887
rect 11341 16841 11387 16887
rect 11499 16841 11545 16887
rect 11658 16841 11704 16887
rect 11816 16841 11862 16887
rect 11974 16841 12020 16887
rect 12132 16841 12178 16887
rect 12290 16841 12336 16887
rect 12448 16841 12494 16887
rect 12606 16841 12652 16887
rect 12764 16841 12810 16887
rect 12922 16841 12968 16887
rect 13081 16841 13127 16887
rect 13239 16841 13285 16887
rect 13397 16841 13443 16887
rect 13555 16841 13601 16887
rect 13713 16841 13759 16887
rect 13871 16841 13917 16887
rect 14029 16841 14075 16887
rect 14187 16841 14233 16887
rect 14345 16841 14391 16887
rect 14504 16841 14550 16887
rect 14662 16841 14708 16887
rect 14820 16841 14866 16887
rect 14978 16841 15024 16887
rect 15136 16841 15182 16887
rect 15294 16841 15340 16887
rect 15452 16841 15498 16887
rect 15610 16841 15656 16887
rect 15768 16841 15814 16887
rect 15927 16841 15973 16887
rect 16085 16841 16131 16887
rect 16243 16841 16289 16887
rect 16401 16841 16447 16887
rect 16559 16841 16605 16887
rect 16717 16841 16763 16887
rect 16875 16841 16921 16887
rect 17033 16841 17079 16887
rect 17192 16841 17238 16887
rect 17350 16841 17396 16887
rect 17508 16841 17554 16887
rect 17666 16841 17712 16887
rect 17824 16841 17870 16887
rect 17982 16841 18028 16887
rect 18140 16841 18186 16887
rect 18298 16841 18344 16887
rect 18456 16841 18502 16887
rect 18615 16841 18661 16887
rect 18773 16841 18819 16887
rect 18931 16841 18977 16887
rect 19089 16841 19135 16887
rect 19247 16841 19293 16887
rect 19405 16841 19451 16887
rect 19563 16841 19609 16887
rect 19721 16841 19767 16887
rect 19879 16841 19925 16887
rect 20038 16841 20084 16887
rect 2586 12217 2820 12263
rect 3706 12217 3940 12263
rect 4826 12217 5060 12263
rect 5946 12217 6180 12263
rect 7066 12217 7300 12263
rect 8186 12217 8420 12263
rect 9306 12217 9540 12263
rect 10426 12217 10660 12263
rect 11546 12217 11780 12263
rect 12666 12217 12900 12263
rect 13786 12217 14020 12263
rect 14906 12217 15140 12263
rect 16026 12217 16260 12263
rect 17146 12217 17380 12263
rect 18266 12217 18500 12263
rect 19386 12217 19620 12263
rect 2256 7848 2302 7894
rect 2256 7685 2302 7731
rect 2256 7522 2302 7568
rect 2256 7359 2302 7405
rect 2256 7196 2302 7242
rect 2256 7032 2302 7078
rect 2256 6869 2302 6915
rect 2256 6706 2302 6752
rect 2256 6542 2302 6588
rect 2256 6379 2302 6425
rect 2256 6216 2302 6262
rect 2256 6052 2302 6098
rect 2256 5889 2302 5935
rect 2256 5726 2302 5772
rect 2256 5563 2302 5609
rect 2256 5400 2302 5446
rect 3947 7848 3993 7894
rect 3947 7685 3993 7731
rect 3947 7522 3993 7568
rect 3947 7359 3993 7405
rect 3947 7196 3993 7242
rect 3947 7032 3993 7078
rect 3947 6869 3993 6915
rect 3947 6706 3993 6752
rect 3947 6542 3993 6588
rect 3947 6379 3993 6425
rect 3947 6216 3993 6262
rect 3947 6052 3993 6098
rect 3947 5889 3993 5935
rect 3947 5726 3993 5772
rect 3947 5563 3993 5609
rect 3947 5400 3993 5446
rect 5638 7848 5684 7894
rect 5638 7685 5684 7731
rect 5638 7522 5684 7568
rect 5638 7359 5684 7405
rect 5638 7196 5684 7242
rect 5638 7032 5684 7078
rect 5638 6869 5684 6915
rect 5638 6706 5684 6752
rect 5638 6542 5684 6588
rect 5638 6379 5684 6425
rect 5638 6216 5684 6262
rect 5638 6052 5684 6098
rect 5638 5889 5684 5935
rect 5638 5726 5684 5772
rect 5638 5563 5684 5609
rect 5638 5400 5684 5446
rect 7727 6762 7773 6808
rect 7885 6762 7931 6808
rect 8043 6762 8089 6808
rect 8201 6762 8247 6808
rect 8359 6762 8405 6808
rect 8517 6762 8563 6808
rect 9360 6762 9406 6808
rect 9518 6762 9564 6808
rect 9676 6762 9722 6808
rect 9834 6762 9880 6808
rect 9992 6762 10038 6808
rect 10150 6762 10196 6808
rect 10994 6762 11040 6808
rect 11152 6762 11198 6808
rect 11310 6762 11356 6808
rect 11468 6762 11514 6808
rect 11626 6762 11672 6808
rect 11784 6762 11830 6808
rect 12628 6762 12674 6808
rect 12786 6762 12832 6808
rect 12944 6762 12990 6808
rect 13102 6762 13148 6808
rect 13260 6762 13306 6808
rect 13418 6762 13464 6808
rect 9931 1061 9977 1107
rect 10089 1061 10135 1107
rect 10247 1061 10293 1107
rect 10405 1061 10451 1107
rect 10563 1061 10609 1107
rect 10721 1061 10767 1107
rect 10879 1061 10925 1107
rect 11037 1061 11083 1107
rect 11195 1061 11241 1107
rect 11354 1061 11400 1107
rect 11512 1061 11558 1107
rect 11670 1061 11716 1107
rect 11828 1061 11874 1107
rect 11986 1061 12032 1107
rect 12144 1061 12190 1107
rect 12303 1061 12349 1107
rect 12461 1061 12507 1107
rect 12619 1061 12665 1107
rect 12777 1061 12823 1107
rect 12935 1061 12981 1107
rect 13093 1061 13139 1107
rect 13251 1061 13297 1107
rect 13409 1061 13455 1107
rect 13567 1061 13613 1107
rect 9931 897 9977 943
rect 10089 897 10135 943
rect 10247 897 10293 943
rect 10405 897 10451 943
rect 10563 897 10609 943
rect 10721 897 10767 943
rect 10879 897 10925 943
rect 11037 897 11083 943
rect 11195 897 11241 943
rect 11354 897 11400 943
rect 11512 897 11558 943
rect 11670 897 11716 943
rect 11828 897 11874 943
rect 11986 897 12032 943
rect 12144 897 12190 943
rect 12303 897 12349 943
rect 12461 897 12507 943
rect 12619 897 12665 943
rect 12777 897 12823 943
rect 12935 897 12981 943
rect 13093 897 13139 943
rect 13251 897 13297 943
rect 13409 897 13455 943
rect 13567 897 13613 943
<< polysilicon >>
rect 1735 28697 1854 28726
rect 1959 28697 2078 28726
rect 2183 28697 2302 28726
rect 2407 28697 2526 28726
rect 1734 28653 1854 28697
rect 1958 28653 2078 28697
rect 2182 28653 2302 28697
rect 2406 28653 2526 28697
rect 2630 28697 2749 28726
rect 2854 28697 2973 28726
rect 3078 28697 3197 28726
rect 3302 28697 3421 28726
rect 3527 28697 3646 28726
rect 3751 28697 3870 28726
rect 3975 28697 4094 28726
rect 4199 28697 4318 28726
rect 2630 28653 2750 28697
rect 2854 28653 2974 28697
rect 3078 28653 3198 28697
rect 3302 28653 3422 28697
rect 3526 28653 3646 28697
rect 3750 28653 3870 28697
rect 3974 28653 4094 28697
rect 4198 28653 4318 28697
rect 4422 28697 4541 28726
rect 4646 28697 4765 28726
rect 4870 28697 4989 28726
rect 5094 28697 5213 28726
rect 9114 28697 9233 28726
rect 9338 28697 9457 28726
rect 9562 28697 9681 28726
rect 9786 28697 9905 28726
rect 4422 28653 4542 28697
rect 4646 28653 4766 28697
rect 4870 28653 4990 28697
rect 5094 28653 5214 28697
rect 9113 28653 9233 28697
rect 9337 28653 9457 28697
rect 9561 28653 9681 28697
rect 9785 28653 9905 28697
rect 10009 28697 10128 28726
rect 10233 28697 10352 28726
rect 10457 28697 10576 28726
rect 10681 28697 10800 28726
rect 10906 28697 11025 28726
rect 11130 28697 11249 28726
rect 11354 28697 11473 28726
rect 11578 28697 11697 28726
rect 10009 28653 10129 28697
rect 10233 28653 10353 28697
rect 10457 28653 10577 28697
rect 10681 28653 10801 28697
rect 10905 28653 11025 28697
rect 11129 28653 11249 28697
rect 11353 28653 11473 28697
rect 11577 28653 11697 28697
rect 11801 28697 11920 28726
rect 12025 28697 12144 28726
rect 12249 28697 12368 28726
rect 12473 28697 12592 28726
rect 11801 28653 11921 28697
rect 12025 28653 12145 28697
rect 12249 28653 12369 28697
rect 12473 28653 12593 28697
rect 6008 28095 6128 28139
rect 6232 28095 6352 28139
rect 6568 28026 6652 28045
rect 6568 27886 6587 28026
rect 6633 27886 6652 28026
rect 7602 28009 7722 28081
rect 1734 27674 1854 27745
rect 1958 27674 2078 27745
rect 2182 27674 2302 27745
rect 2406 27674 2526 27745
rect 1734 27537 2526 27674
rect 1734 27465 1854 27537
rect 1958 27465 2078 27537
rect 2182 27465 2302 27537
rect 2406 27465 2526 27537
rect 2630 27674 2750 27745
rect 2854 27674 2974 27745
rect 3078 27674 3198 27745
rect 3302 27674 3422 27745
rect 2630 27537 3422 27674
rect 2630 27465 2750 27537
rect 2854 27465 2974 27537
rect 3078 27465 3198 27537
rect 3302 27465 3422 27537
rect 3526 27674 3646 27745
rect 3750 27674 3870 27745
rect 3974 27674 4094 27745
rect 4198 27674 4318 27745
rect 3526 27537 4318 27674
rect 3526 27465 3646 27537
rect 3750 27465 3870 27537
rect 3974 27465 4094 27537
rect 4198 27465 4318 27537
rect 4422 27674 4542 27745
rect 4646 27674 4766 27745
rect 4870 27674 4990 27745
rect 5094 27674 5214 27745
rect 6008 27702 6128 27821
rect 6232 27761 6352 27821
rect 6568 27761 6652 27886
rect 6232 27748 6652 27761
rect 4422 27537 5214 27674
rect 5835 27683 6128 27702
rect 5835 27637 5854 27683
rect 5994 27637 6128 27683
rect 5835 27618 6128 27637
rect 4422 27465 4542 27537
rect 4646 27465 4766 27537
rect 4870 27465 4990 27537
rect 5094 27465 5214 27537
rect 6008 27427 6128 27618
rect 6231 27655 6652 27748
rect 6231 27427 6351 27655
rect 6456 27644 6652 27655
rect 6456 27427 6576 27644
rect 6763 27574 6957 27632
rect 6763 27548 6782 27574
rect 6679 27528 6782 27548
rect 6922 27528 6957 27574
rect 6679 27488 6957 27528
rect 6679 27427 6799 27488
rect 7602 27463 7722 27817
rect 23872 28203 23992 28247
rect 24096 28203 24216 28247
rect 13387 28095 13507 28139
rect 13611 28095 13731 28139
rect 16780 28133 16898 28162
rect 17004 28133 17122 28162
rect 17228 28133 17346 28162
rect 17452 28133 17570 28162
rect 17676 28133 17794 28162
rect 17900 28133 18018 28162
rect 18414 28133 18532 28162
rect 18638 28133 18756 28162
rect 18862 28133 18980 28162
rect 19086 28133 19204 28162
rect 19310 28133 19428 28162
rect 19534 28133 19652 28162
rect 20047 28133 20165 28162
rect 20271 28133 20389 28162
rect 20495 28133 20613 28162
rect 20719 28133 20837 28162
rect 20943 28133 21061 28162
rect 21167 28133 21285 28162
rect 21681 28133 21799 28162
rect 21905 28133 22023 28162
rect 22129 28133 22247 28162
rect 22353 28133 22471 28162
rect 22577 28133 22695 28162
rect 22801 28133 22919 28162
rect 16779 28089 16899 28133
rect 17003 28089 17123 28133
rect 17227 28089 17347 28133
rect 17451 28089 17571 28133
rect 17675 28089 17795 28133
rect 17899 28089 18019 28133
rect 18413 28089 18533 28133
rect 18637 28089 18757 28133
rect 18861 28089 18981 28133
rect 19085 28089 19205 28133
rect 19309 28089 19429 28133
rect 19533 28089 19653 28133
rect 20046 28089 20166 28133
rect 20270 28089 20390 28133
rect 20494 28089 20614 28133
rect 20718 28089 20838 28133
rect 20942 28089 21062 28133
rect 21166 28089 21286 28133
rect 21680 28089 21800 28133
rect 21904 28089 22024 28133
rect 22128 28089 22248 28133
rect 22352 28089 22472 28133
rect 22576 28089 22696 28133
rect 22800 28089 22920 28133
rect 13947 28026 14031 28045
rect 13947 27886 13966 28026
rect 14012 27886 14031 28026
rect 14981 28009 15101 28081
rect 9113 27674 9233 27745
rect 9337 27674 9457 27745
rect 9561 27674 9681 27745
rect 9785 27674 9905 27745
rect 9113 27537 9905 27674
rect 9113 27465 9233 27537
rect 9337 27465 9457 27537
rect 9561 27465 9681 27537
rect 9785 27465 9905 27537
rect 10009 27674 10129 27745
rect 10233 27674 10353 27745
rect 10457 27674 10577 27745
rect 10681 27674 10801 27745
rect 10009 27537 10801 27674
rect 10009 27465 10129 27537
rect 10233 27465 10353 27537
rect 10457 27465 10577 27537
rect 10681 27465 10801 27537
rect 10905 27674 11025 27745
rect 11129 27674 11249 27745
rect 11353 27674 11473 27745
rect 11577 27674 11697 27745
rect 10905 27537 11697 27674
rect 10905 27465 11025 27537
rect 11129 27465 11249 27537
rect 11353 27465 11473 27537
rect 11577 27465 11697 27537
rect 11801 27674 11921 27745
rect 12025 27674 12145 27745
rect 12249 27674 12369 27745
rect 12473 27674 12593 27745
rect 13387 27702 13507 27821
rect 13611 27761 13731 27821
rect 13947 27761 14031 27886
rect 13611 27748 14031 27761
rect 11801 27537 12593 27674
rect 13214 27683 13507 27702
rect 13214 27637 13233 27683
rect 13373 27637 13507 27683
rect 13214 27618 13507 27637
rect 11801 27465 11921 27537
rect 12025 27465 12145 27537
rect 12249 27465 12369 27537
rect 12473 27465 12593 27537
rect 7484 27388 7828 27463
rect 7484 27328 7604 27388
rect 7708 27328 7828 27388
rect 6008 27013 6128 27086
rect 6231 27013 6351 27086
rect 6456 27013 6576 27086
rect 6679 27013 6799 27086
rect 7484 27040 7604 27100
rect 7708 27040 7828 27100
rect 7484 27021 7828 27040
rect 7484 26975 7550 27021
rect 7784 26975 7828 27021
rect 7484 26956 7828 26975
rect 6166 26744 6286 26788
rect 7857 26744 7977 26788
rect 6680 26503 6799 26531
rect 6680 26459 6800 26503
rect 6166 25264 6286 25336
rect 6680 25264 6800 25415
rect 8371 26503 8490 26531
rect 8371 26459 8491 26503
rect 7857 25264 7977 25336
rect 8371 25264 8491 25415
rect 5880 25218 6286 25264
rect 1734 25135 1854 25197
rect 1958 25135 2078 25197
rect 2182 25135 2302 25197
rect 2406 25135 2526 25197
rect 1734 25088 2526 25135
rect 1734 25042 1895 25088
rect 2317 25042 2526 25088
rect 1734 24998 2526 25042
rect 2630 25135 2750 25197
rect 2854 25135 2974 25197
rect 3078 25135 3198 25197
rect 3302 25135 3422 25197
rect 2630 25088 3422 25135
rect 2630 25042 2839 25088
rect 3261 25042 3422 25088
rect 2630 24998 3422 25042
rect 3526 25135 3646 25197
rect 3750 25135 3870 25197
rect 3974 25135 4094 25197
rect 4198 25135 4318 25197
rect 3526 25088 4318 25135
rect 3526 25042 3687 25088
rect 4109 25042 4318 25088
rect 3526 24998 4318 25042
rect 4422 25135 4542 25197
rect 4646 25135 4766 25197
rect 4870 25135 4990 25197
rect 5094 25135 5214 25197
rect 4422 25088 5214 25135
rect 5880 25172 5954 25218
rect 6000 25172 6112 25218
rect 6158 25172 6286 25218
rect 5880 25126 6286 25172
rect 6390 25218 6800 25264
rect 6390 25172 6464 25218
rect 6510 25172 6622 25218
rect 6668 25172 6800 25218
rect 6390 25126 6800 25172
rect 7571 25218 7977 25264
rect 7571 25172 7645 25218
rect 7691 25172 7803 25218
rect 7849 25172 7977 25218
rect 7571 25126 7977 25172
rect 8081 25218 8491 25264
rect 8081 25172 8155 25218
rect 8201 25172 8313 25218
rect 8359 25172 8491 25218
rect 13387 27427 13507 27618
rect 13610 27655 14031 27748
rect 13610 27427 13730 27655
rect 13835 27644 14031 27655
rect 13835 27427 13955 27644
rect 14142 27574 14336 27632
rect 14142 27548 14161 27574
rect 14058 27528 14161 27548
rect 14301 27528 14336 27574
rect 14058 27488 14336 27528
rect 14058 27427 14178 27488
rect 14981 27463 15101 27817
rect 14863 27388 15207 27463
rect 14863 27328 14983 27388
rect 15087 27328 15207 27388
rect 25467 28089 25587 28133
rect 24404 28037 24488 28056
rect 24404 27897 24423 28037
rect 24469 27897 24488 28037
rect 23872 27740 23992 27821
rect 23587 27694 23992 27740
rect 23587 27648 23661 27694
rect 23707 27648 23819 27694
rect 23865 27648 23992 27694
rect 23587 27602 23992 27648
rect 23872 27541 23992 27602
rect 24096 27761 24216 27821
rect 24404 27761 24488 27897
rect 24096 27698 24488 27761
rect 24096 27676 24440 27698
rect 24096 27541 24216 27676
rect 24320 27541 24440 27676
rect 24544 27666 24748 27685
rect 24544 27620 24683 27666
rect 24729 27620 24748 27666
rect 24544 27601 24748 27620
rect 24544 27541 24664 27601
rect 25467 27577 25587 27817
rect 16779 27110 16899 27181
rect 17003 27110 17123 27181
rect 17227 27110 17347 27181
rect 13387 27013 13507 27086
rect 13610 27013 13730 27086
rect 13835 27013 13955 27086
rect 14058 27013 14178 27086
rect 14863 27040 14983 27100
rect 15087 27040 15207 27100
rect 14863 27021 15207 27040
rect 14863 26975 14929 27021
rect 15163 26975 15207 27021
rect 14863 26956 15207 26975
rect 16779 26973 17347 27110
rect 16779 26901 16899 26973
rect 17003 26901 17123 26973
rect 17227 26901 17347 26973
rect 17451 27110 17571 27181
rect 17675 27110 17795 27181
rect 17899 27110 18019 27181
rect 17451 26973 18019 27110
rect 17451 26901 17571 26973
rect 17675 26901 17795 26973
rect 17899 26901 18019 26973
rect 18413 27110 18533 27181
rect 18637 27110 18757 27181
rect 18861 27110 18981 27181
rect 18413 26973 18981 27110
rect 18413 26901 18533 26973
rect 18637 26901 18757 26973
rect 18861 26901 18981 26973
rect 19085 27110 19205 27181
rect 19309 27110 19429 27181
rect 19533 27110 19653 27181
rect 19085 26973 19653 27110
rect 19085 26901 19205 26973
rect 19309 26901 19429 26973
rect 19533 26901 19653 26973
rect 20046 27110 20166 27181
rect 20270 27110 20390 27181
rect 20494 27110 20614 27181
rect 20046 26973 20614 27110
rect 20046 26901 20166 26973
rect 20270 26901 20390 26973
rect 20494 26901 20614 26973
rect 20718 27110 20838 27181
rect 20942 27110 21062 27181
rect 21166 27110 21286 27181
rect 20718 26973 21286 27110
rect 20718 26901 20838 26973
rect 20942 26901 21062 26973
rect 21166 26901 21286 26973
rect 21680 27110 21800 27181
rect 21904 27110 22024 27181
rect 22128 27110 22248 27181
rect 21680 26973 22248 27110
rect 21680 26901 21800 26973
rect 21904 26901 22024 26973
rect 22128 26901 22248 26973
rect 22352 27110 22472 27181
rect 22576 27110 22696 27181
rect 22800 27110 22920 27181
rect 22352 26973 22920 27110
rect 25348 27502 25692 27577
rect 25348 27442 25468 27502
rect 25572 27442 25692 27502
rect 23872 27013 23992 27086
rect 24096 27013 24216 27086
rect 24320 27013 24440 27086
rect 24544 27013 24664 27086
rect 25348 27040 25468 27100
rect 25572 27040 25692 27100
rect 25348 27021 25692 27040
rect 22352 26901 22472 26973
rect 22576 26901 22696 26973
rect 22800 26901 22920 26973
rect 25348 26975 25392 27021
rect 25626 26975 25692 27021
rect 25348 26956 25692 26975
rect 13545 26744 13665 26788
rect 15236 26744 15356 26788
rect 14059 26503 14178 26531
rect 14059 26459 14179 26503
rect 13545 25264 13665 25336
rect 14059 25264 14179 25415
rect 15750 26503 15869 26531
rect 15750 26459 15870 26503
rect 15236 25264 15356 25336
rect 15750 25264 15870 25415
rect 13259 25218 13665 25264
rect 8081 25126 8491 25172
rect 4422 25042 4631 25088
rect 5053 25042 5214 25088
rect 4422 24998 5214 25042
rect 6166 25015 6286 25126
rect 6680 25016 6800 25126
rect 1893 24607 2012 24634
rect 2117 24607 2236 24634
rect 1892 24563 2012 24607
rect 2116 24563 2236 24607
rect 2920 24607 3039 24634
rect 3144 24607 3263 24634
rect 3685 24607 3804 24634
rect 3909 24607 4028 24634
rect 2920 24563 3040 24607
rect 3144 24563 3264 24607
rect 3684 24563 3804 24607
rect 3908 24563 4028 24607
rect 4712 24607 4831 24634
rect 4936 24607 5055 24634
rect 4712 24563 4832 24607
rect 4936 24563 5056 24607
rect 1892 21408 2012 21523
rect 1855 21363 2048 21408
rect 1855 21317 1929 21363
rect 1975 21317 2048 21363
rect 1855 21271 2048 21317
rect 1892 20551 2012 21271
rect 2116 21000 2236 21523
rect 2079 20955 2272 21000
rect 2079 20909 2153 20955
rect 2199 20909 2272 20955
rect 2079 20863 2272 20909
rect 2116 20551 2236 20863
rect 2920 20800 3040 21523
rect 3144 21408 3264 21523
rect 3107 21363 3300 21408
rect 3107 21317 3181 21363
rect 3227 21317 3300 21363
rect 3107 21271 3300 21317
rect 2883 20755 3076 20800
rect 2883 20709 2957 20755
rect 3003 20709 3076 20755
rect 2883 20663 3076 20709
rect 2920 20551 3040 20663
rect 3144 20551 3264 21271
rect 3684 21204 3804 21523
rect 3647 21159 3840 21204
rect 3647 21113 3721 21159
rect 3767 21113 3840 21159
rect 3647 21067 3840 21113
rect 3684 20551 3804 21067
rect 3908 21000 4028 21523
rect 3871 20955 4064 21000
rect 3871 20909 3945 20955
rect 3991 20909 4064 20955
rect 3871 20863 4064 20909
rect 3908 20551 4028 20863
rect 4712 20800 4832 21523
rect 4936 21204 5056 21523
rect 7857 25015 7977 25126
rect 8371 25016 8491 25126
rect 9113 25135 9233 25197
rect 9337 25135 9457 25197
rect 9561 25135 9681 25197
rect 9785 25135 9905 25197
rect 9113 25088 9905 25135
rect 9113 25042 9274 25088
rect 9696 25042 9905 25088
rect 6680 22340 6800 22384
rect 6680 22311 6799 22340
rect 9113 24998 9905 25042
rect 10009 25135 10129 25197
rect 10233 25135 10353 25197
rect 10457 25135 10577 25197
rect 10681 25135 10801 25197
rect 10009 25088 10801 25135
rect 10009 25042 10218 25088
rect 10640 25042 10801 25088
rect 10009 24998 10801 25042
rect 10905 25135 11025 25197
rect 11129 25135 11249 25197
rect 11353 25135 11473 25197
rect 11577 25135 11697 25197
rect 10905 25088 11697 25135
rect 10905 25042 11066 25088
rect 11488 25042 11697 25088
rect 10905 24998 11697 25042
rect 11801 25135 11921 25197
rect 12025 25135 12145 25197
rect 12249 25135 12369 25197
rect 12473 25135 12593 25197
rect 11801 25088 12593 25135
rect 13259 25172 13333 25218
rect 13379 25172 13491 25218
rect 13537 25172 13665 25218
rect 13259 25126 13665 25172
rect 13769 25218 14179 25264
rect 13769 25172 13843 25218
rect 13889 25172 14001 25218
rect 14047 25172 14179 25218
rect 13769 25126 14179 25172
rect 14950 25218 15356 25264
rect 14950 25172 15024 25218
rect 15070 25172 15182 25218
rect 15228 25172 15356 25218
rect 14950 25126 15356 25172
rect 15460 25218 15870 25264
rect 15460 25172 15534 25218
rect 15580 25172 15692 25218
rect 15738 25172 15870 25218
rect 15460 25126 15870 25172
rect 11801 25042 12010 25088
rect 12432 25042 12593 25088
rect 11801 24998 12593 25042
rect 13545 25015 13665 25126
rect 14059 25016 14179 25126
rect 9272 24607 9391 24634
rect 9496 24607 9615 24634
rect 9271 24563 9391 24607
rect 9495 24563 9615 24607
rect 10299 24607 10418 24634
rect 10523 24607 10642 24634
rect 11064 24607 11183 24634
rect 11288 24607 11407 24634
rect 10299 24563 10419 24607
rect 10523 24563 10643 24607
rect 11063 24563 11183 24607
rect 11287 24563 11407 24607
rect 12091 24607 12210 24634
rect 12315 24607 12434 24634
rect 12091 24563 12211 24607
rect 12315 24563 12435 24607
rect 8371 22340 8491 22384
rect 8371 22311 8490 22340
rect 6166 21433 6286 21477
rect 7857 21433 7977 21477
rect 6166 21404 6285 21433
rect 7857 21404 7976 21433
rect 9271 21408 9391 21523
rect 9234 21363 9427 21408
rect 9234 21317 9308 21363
rect 9354 21317 9427 21363
rect 9234 21271 9427 21317
rect 4899 21159 5092 21204
rect 4899 21113 4973 21159
rect 5019 21113 5092 21159
rect 4899 21067 5092 21113
rect 4675 20755 4868 20800
rect 4675 20709 4749 20755
rect 4795 20709 4868 20755
rect 4675 20663 4868 20709
rect 4712 20551 4832 20663
rect 4936 20551 5056 21067
rect 9271 20551 9391 21271
rect 9495 21000 9615 21523
rect 9458 20955 9651 21000
rect 9458 20909 9532 20955
rect 9578 20909 9651 20955
rect 9458 20863 9651 20909
rect 9495 20551 9615 20863
rect 10299 20800 10419 21523
rect 10523 21408 10643 21523
rect 10486 21363 10679 21408
rect 10486 21317 10560 21363
rect 10606 21317 10679 21363
rect 10486 21271 10679 21317
rect 10262 20755 10455 20800
rect 10262 20709 10336 20755
rect 10382 20709 10455 20755
rect 10262 20663 10455 20709
rect 10299 20551 10419 20663
rect 10523 20551 10643 21271
rect 11063 21204 11183 21523
rect 11026 21159 11219 21204
rect 11026 21113 11100 21159
rect 11146 21113 11219 21159
rect 11026 21067 11219 21113
rect 11063 20551 11183 21067
rect 11287 21000 11407 21523
rect 11250 20955 11443 21000
rect 11250 20909 11324 20955
rect 11370 20909 11443 20955
rect 11250 20863 11443 20909
rect 11287 20551 11407 20863
rect 12091 20800 12211 21523
rect 12315 21204 12435 21523
rect 15236 25015 15356 25126
rect 15750 25016 15870 25126
rect 14059 22340 14179 22384
rect 14059 22311 14178 22340
rect 24031 26787 24150 26815
rect 24545 26787 24664 26815
rect 25721 26787 25840 26815
rect 26235 26787 26354 26815
rect 27412 26787 27531 26815
rect 27926 26787 28045 26815
rect 24031 26743 24151 26787
rect 24545 26743 24665 26787
rect 25721 26743 25841 26787
rect 26235 26743 26355 26787
rect 27412 26743 27532 26787
rect 27926 26743 28046 26787
rect 24031 25383 24151 25427
rect 24545 25383 24665 25427
rect 25721 25383 25841 25427
rect 26235 25383 26355 25427
rect 27412 25383 27532 25427
rect 27926 25383 28046 25427
rect 24031 25355 24150 25383
rect 24545 25355 24664 25383
rect 25721 25355 25840 25383
rect 26235 25355 26354 25383
rect 27412 25355 27531 25383
rect 27926 25355 28045 25383
rect 23745 25309 24150 25355
rect 23745 25263 23819 25309
rect 23865 25263 23977 25309
rect 24023 25263 24150 25309
rect 23745 25217 24150 25263
rect 24255 25309 24664 25355
rect 24255 25263 24329 25309
rect 24375 25263 24487 25309
rect 24533 25263 24664 25309
rect 24255 25217 24664 25263
rect 25435 25309 25840 25355
rect 25435 25263 25509 25309
rect 25555 25263 25667 25309
rect 25713 25263 25840 25309
rect 25435 25217 25840 25263
rect 25945 25309 26354 25355
rect 25945 25263 26019 25309
rect 26065 25263 26177 25309
rect 26223 25263 26354 25309
rect 25945 25217 26354 25263
rect 27126 25309 27531 25355
rect 27126 25263 27200 25309
rect 27246 25263 27358 25309
rect 27404 25263 27531 25309
rect 27126 25217 27531 25263
rect 27636 25309 28045 25355
rect 27636 25263 27710 25309
rect 27756 25263 27868 25309
rect 27914 25263 28045 25309
rect 27636 25217 28045 25263
rect 24031 25191 24150 25217
rect 24545 25191 24664 25217
rect 25721 25191 25840 25217
rect 26235 25191 26354 25217
rect 27412 25191 27531 25217
rect 27926 25191 28045 25217
rect 24031 25147 24151 25191
rect 24545 25147 24665 25191
rect 25721 25147 25841 25191
rect 26235 25147 26355 25191
rect 27412 25147 27532 25191
rect 27926 25147 28046 25191
rect 16779 24571 16899 24633
rect 17003 24571 17123 24633
rect 17227 24571 17347 24633
rect 16779 24527 17347 24571
rect 16779 24481 16889 24527
rect 17217 24481 17347 24527
rect 16779 24434 17347 24481
rect 17451 24571 17571 24633
rect 17675 24571 17795 24633
rect 17899 24571 18019 24633
rect 17451 24527 18019 24571
rect 17451 24481 17581 24527
rect 17909 24481 18019 24527
rect 17451 24434 18019 24481
rect 18413 24571 18533 24633
rect 18637 24571 18757 24633
rect 18861 24571 18981 24633
rect 18413 24527 18981 24571
rect 18413 24481 18523 24527
rect 18851 24481 18981 24527
rect 18413 24434 18981 24481
rect 19085 24571 19205 24633
rect 19309 24571 19429 24633
rect 19533 24571 19653 24633
rect 19085 24527 19653 24571
rect 19085 24481 19215 24527
rect 19543 24481 19653 24527
rect 19085 24434 19653 24481
rect 20046 24571 20166 24633
rect 20270 24571 20390 24633
rect 20494 24571 20614 24633
rect 20046 24527 20614 24571
rect 20046 24481 20156 24527
rect 20484 24481 20614 24527
rect 20046 24434 20614 24481
rect 20718 24571 20838 24633
rect 20942 24571 21062 24633
rect 21166 24571 21286 24633
rect 20718 24527 21286 24571
rect 20718 24481 20848 24527
rect 21176 24481 21286 24527
rect 20718 24434 21286 24481
rect 21680 24571 21800 24633
rect 21904 24571 22024 24633
rect 22128 24571 22248 24633
rect 21680 24527 22248 24571
rect 21680 24481 21790 24527
rect 22118 24481 22248 24527
rect 21680 24434 22248 24481
rect 22352 24571 22472 24633
rect 22576 24571 22696 24633
rect 22800 24571 22920 24633
rect 22352 24527 22920 24571
rect 22352 24481 22482 24527
rect 22810 24481 22920 24527
rect 22352 24434 22920 24481
rect 16780 24041 16898 24070
rect 17004 24041 17122 24070
rect 17228 24041 17346 24070
rect 17452 24041 17570 24070
rect 17676 24041 17794 24070
rect 17900 24041 18018 24070
rect 18414 24041 18532 24070
rect 18638 24041 18756 24070
rect 18862 24041 18980 24070
rect 19086 24041 19204 24070
rect 19310 24041 19428 24070
rect 19534 24041 19652 24070
rect 20047 24041 20165 24070
rect 20271 24041 20389 24070
rect 20495 24041 20613 24070
rect 20719 24041 20837 24070
rect 20943 24041 21061 24070
rect 21167 24041 21285 24070
rect 21681 24041 21799 24070
rect 21905 24041 22023 24070
rect 22129 24041 22247 24070
rect 22353 24041 22471 24070
rect 22577 24041 22695 24070
rect 22801 24041 22919 24070
rect 16779 23997 16899 24041
rect 17003 23997 17123 24041
rect 17227 23997 17347 24041
rect 17451 23997 17571 24041
rect 17675 23997 17795 24041
rect 17899 23997 18019 24041
rect 18413 23997 18533 24041
rect 18637 23997 18757 24041
rect 18861 23997 18981 24041
rect 19085 23997 19205 24041
rect 19309 23997 19429 24041
rect 19533 23997 19653 24041
rect 20046 23997 20166 24041
rect 20270 23997 20390 24041
rect 20494 23997 20614 24041
rect 20718 23997 20838 24041
rect 20942 23997 21062 24041
rect 21166 23997 21286 24041
rect 21680 23997 21800 24041
rect 21904 23997 22024 24041
rect 22128 23997 22248 24041
rect 22352 23997 22472 24041
rect 22576 23997 22696 24041
rect 22800 23997 22920 24041
rect 15750 22340 15870 22384
rect 15750 22311 15869 22340
rect 16779 21809 16899 21911
rect 16742 21764 16935 21809
rect 16742 21718 16816 21764
rect 16862 21718 16935 21764
rect 16742 21672 16935 21718
rect 13545 21433 13665 21477
rect 15236 21433 15356 21477
rect 13545 21404 13664 21433
rect 15236 21404 15355 21433
rect 12278 21159 12471 21204
rect 12278 21113 12352 21159
rect 12398 21113 12471 21159
rect 12278 21067 12471 21113
rect 12054 20755 12247 20800
rect 12054 20709 12128 20755
rect 12174 20709 12247 20755
rect 12054 20663 12247 20709
rect 12091 20551 12211 20663
rect 12315 20551 12435 21067
rect 16779 20538 16899 21672
rect 17003 21609 17123 21911
rect 16966 21564 17159 21609
rect 16966 21518 17040 21564
rect 17086 21518 17159 21564
rect 16966 21472 17159 21518
rect 17003 20538 17123 21472
rect 17227 21405 17347 21911
rect 17451 21405 17571 21911
rect 17675 21609 17795 21911
rect 17899 21809 18019 21911
rect 18413 21809 18533 21911
rect 17862 21764 18055 21809
rect 17862 21718 17936 21764
rect 17982 21718 18055 21764
rect 17862 21672 18055 21718
rect 18375 21764 18568 21809
rect 18375 21718 18449 21764
rect 18495 21718 18568 21764
rect 18375 21672 18568 21718
rect 17638 21564 17831 21609
rect 17638 21518 17712 21564
rect 17758 21518 17831 21564
rect 17638 21472 17831 21518
rect 17190 21360 17383 21405
rect 17190 21314 17264 21360
rect 17310 21314 17383 21360
rect 17190 21268 17383 21314
rect 17451 21268 17572 21405
rect 17227 20538 17347 21268
rect 17451 20800 17571 21268
rect 17414 20755 17607 20800
rect 17414 20709 17488 20755
rect 17534 20709 17607 20755
rect 17414 20663 17607 20709
rect 17451 20538 17571 20663
rect 17675 20538 17795 21472
rect 17899 20538 18019 21672
rect 18413 20538 18533 21672
rect 18637 21002 18757 21911
rect 18861 21405 18981 21911
rect 19085 21405 19205 21911
rect 18823 21360 19016 21405
rect 18823 21314 18897 21360
rect 18943 21314 19016 21360
rect 18823 21268 19016 21314
rect 19085 21268 19206 21405
rect 18599 20957 18792 21002
rect 18599 20911 18673 20957
rect 18719 20911 18792 20957
rect 18599 20865 18792 20911
rect 18637 20538 18757 20865
rect 18861 20538 18981 21268
rect 19085 20800 19205 21268
rect 19309 21002 19429 21911
rect 19533 21809 19653 21911
rect 19495 21764 19688 21809
rect 19495 21718 19569 21764
rect 19615 21718 19688 21764
rect 19495 21672 19688 21718
rect 19271 20957 19464 21002
rect 19271 20911 19345 20957
rect 19391 20911 19464 20957
rect 19271 20865 19464 20911
rect 19047 20755 19240 20800
rect 19047 20709 19121 20755
rect 19167 20709 19240 20755
rect 19047 20663 19240 20709
rect 19085 20538 19205 20663
rect 19309 20538 19429 20865
rect 19533 20538 19653 21672
rect 20046 21204 20166 21911
rect 20270 21609 20390 21911
rect 20233 21564 20426 21609
rect 20233 21518 20307 21564
rect 20353 21518 20426 21564
rect 20233 21472 20426 21518
rect 20009 21159 20202 21204
rect 20009 21113 20083 21159
rect 20129 21113 20202 21159
rect 20009 21067 20202 21113
rect 20046 20538 20166 21067
rect 20270 20538 20390 21472
rect 20494 21405 20614 21911
rect 20718 21405 20838 21911
rect 20942 21609 21062 21911
rect 20905 21564 21098 21609
rect 20905 21518 20979 21564
rect 21025 21518 21098 21564
rect 20905 21472 21098 21518
rect 20457 21360 20650 21405
rect 20457 21314 20531 21360
rect 20577 21314 20650 21360
rect 20457 21268 20650 21314
rect 20718 21268 20839 21405
rect 20494 20538 20614 21268
rect 20718 20800 20838 21268
rect 20681 20755 20874 20800
rect 20681 20709 20755 20755
rect 20801 20709 20874 20755
rect 20681 20663 20874 20709
rect 20718 20538 20838 20663
rect 20942 20538 21062 21472
rect 21166 21204 21286 21911
rect 21680 21204 21800 21911
rect 21129 21159 21322 21204
rect 21129 21113 21203 21159
rect 21249 21113 21322 21159
rect 21129 21067 21322 21113
rect 21643 21159 21836 21204
rect 21643 21113 21717 21159
rect 21763 21113 21836 21159
rect 21643 21067 21836 21113
rect 21166 20538 21286 21067
rect 21680 20538 21800 21067
rect 21904 21002 22024 21911
rect 22128 21405 22248 21911
rect 22352 21405 22472 21911
rect 22091 21360 22284 21405
rect 22091 21314 22165 21360
rect 22211 21314 22284 21360
rect 22091 21268 22284 21314
rect 22352 21268 22473 21405
rect 21867 20957 22060 21002
rect 21867 20911 21941 20957
rect 21987 20911 22060 20957
rect 21867 20865 22060 20911
rect 21904 20538 22024 20865
rect 22128 20538 22248 21268
rect 22352 20800 22472 21268
rect 22576 21002 22696 21911
rect 22800 21204 22920 21911
rect 24031 21837 24151 21881
rect 24545 21837 24665 21881
rect 25721 21837 25841 21881
rect 26235 21837 26355 21881
rect 27412 21837 27532 21881
rect 27926 21837 28046 21881
rect 24031 21808 24150 21837
rect 24545 21808 24664 21837
rect 25721 21808 25840 21837
rect 26235 21808 26354 21837
rect 27412 21808 27531 21837
rect 27926 21808 28045 21837
rect 22763 21159 22956 21204
rect 22763 21113 22837 21159
rect 22883 21113 22956 21159
rect 22763 21067 22956 21113
rect 22539 20957 22732 21002
rect 22539 20911 22613 20957
rect 22659 20911 22732 20957
rect 22539 20865 22732 20911
rect 22315 20755 22508 20800
rect 22315 20709 22389 20755
rect 22435 20709 22508 20755
rect 22315 20663 22508 20709
rect 22352 20538 22472 20663
rect 22576 20538 22696 20865
rect 22800 20538 22920 21067
rect 1892 18029 2012 18101
rect 2116 18029 2236 18101
rect 2920 18029 3040 18101
rect 3144 18029 3264 18101
rect 3684 18029 3804 18101
rect 3908 18029 4028 18101
rect 4712 18029 4832 18101
rect 4936 18029 5056 18101
rect 9271 18029 9391 18101
rect 9495 18029 9615 18101
rect 10299 18029 10419 18101
rect 10523 18029 10643 18101
rect 11063 18029 11183 18101
rect 11287 18029 11407 18101
rect 12091 18029 12211 18101
rect 12315 18029 12435 18101
rect 16779 17970 16899 18043
rect 17003 17970 17123 18043
rect 17227 17970 17347 18043
rect 17451 17970 17571 18043
rect 17675 17970 17795 18043
rect 17899 17970 18019 18043
rect 18413 17970 18533 18043
rect 18637 17970 18757 18043
rect 18861 17970 18981 18043
rect 19085 17970 19205 18043
rect 19309 17970 19429 18043
rect 19533 17970 19653 18043
rect 20046 17970 20166 18043
rect 20270 17970 20390 18043
rect 20494 17970 20614 18043
rect 20718 17970 20838 18043
rect 20942 17970 21062 18043
rect 21166 17970 21286 18043
rect 21680 17970 21800 18043
rect 21904 17970 22024 18043
rect 22128 17970 22248 18043
rect 22352 17970 22472 18043
rect 22576 17970 22696 18043
rect 22800 17970 22920 18043
rect 2070 16585 2190 16629
rect 2518 16585 2638 16629
rect 2742 16585 2862 16629
rect 2966 16585 3086 16629
rect 3190 16585 3310 16629
rect 3638 16585 3758 16629
rect 3862 16585 3982 16629
rect 4086 16585 4206 16629
rect 4310 16585 4430 16629
rect 4758 16585 4878 16629
rect 4982 16585 5102 16629
rect 5206 16585 5326 16629
rect 5430 16585 5550 16629
rect 5878 16585 5998 16629
rect 6102 16585 6222 16629
rect 6326 16585 6446 16629
rect 6550 16585 6670 16629
rect 6998 16585 7118 16629
rect 7222 16585 7342 16629
rect 7446 16585 7566 16629
rect 7670 16585 7790 16629
rect 8118 16585 8238 16629
rect 8342 16585 8462 16629
rect 8566 16585 8686 16629
rect 8790 16585 8910 16629
rect 9238 16585 9358 16629
rect 9462 16585 9582 16629
rect 9686 16585 9806 16629
rect 9910 16585 10030 16629
rect 10358 16585 10478 16629
rect 10582 16585 10702 16629
rect 10806 16585 10926 16629
rect 11030 16585 11150 16629
rect 11478 16585 11598 16629
rect 11702 16585 11822 16629
rect 11926 16585 12046 16629
rect 12150 16585 12270 16629
rect 12598 16585 12718 16629
rect 12822 16585 12942 16629
rect 13046 16585 13166 16629
rect 13270 16585 13390 16629
rect 13718 16585 13838 16629
rect 13942 16585 14062 16629
rect 14166 16585 14286 16629
rect 14390 16585 14510 16629
rect 14838 16585 14958 16629
rect 15062 16585 15182 16629
rect 15286 16585 15406 16629
rect 15510 16585 15630 16629
rect 15958 16585 16078 16629
rect 16182 16585 16302 16629
rect 16406 16585 16526 16629
rect 16630 16585 16750 16629
rect 17078 16585 17198 16629
rect 17302 16585 17422 16629
rect 17526 16585 17646 16629
rect 17750 16585 17870 16629
rect 18198 16585 18318 16629
rect 18422 16585 18542 16629
rect 18646 16585 18766 16629
rect 18870 16585 18990 16629
rect 19318 16585 19438 16629
rect 19542 16585 19662 16629
rect 19766 16585 19886 16629
rect 2070 12427 2190 12585
rect 2070 12381 2089 12427
rect 2135 12381 2190 12427
rect 2518 12477 2638 12585
rect 2742 12477 2862 12585
rect 2966 12477 3086 12585
rect 2518 12458 3086 12477
rect 2518 12412 2916 12458
rect 3056 12412 3086 12458
rect 2518 12393 3086 12412
rect 3190 12427 3310 12585
rect 2070 12362 2190 12381
rect 3190 12381 3209 12427
rect 3255 12381 3310 12427
rect 3638 12477 3758 12585
rect 3862 12477 3982 12585
rect 4086 12477 4206 12585
rect 3638 12458 4206 12477
rect 3638 12412 4036 12458
rect 4176 12412 4206 12458
rect 3638 12393 4206 12412
rect 4310 12427 4430 12585
rect 3190 12362 3310 12381
rect 4310 12381 4329 12427
rect 4375 12381 4430 12427
rect 4758 12477 4878 12585
rect 4982 12477 5102 12585
rect 5206 12477 5326 12585
rect 4758 12458 5326 12477
rect 4758 12412 5156 12458
rect 5296 12412 5326 12458
rect 4758 12393 5326 12412
rect 5430 12427 5550 12585
rect 4310 12362 4430 12381
rect 5430 12381 5449 12427
rect 5495 12381 5550 12427
rect 5878 12477 5998 12585
rect 6102 12477 6222 12585
rect 6326 12477 6446 12585
rect 5878 12458 6446 12477
rect 5878 12412 6276 12458
rect 6416 12412 6446 12458
rect 5878 12393 6446 12412
rect 6550 12427 6670 12585
rect 5430 12362 5550 12381
rect 6550 12381 6569 12427
rect 6615 12381 6670 12427
rect 6998 12477 7118 12585
rect 7222 12477 7342 12585
rect 7446 12477 7566 12585
rect 6998 12458 7566 12477
rect 6998 12412 7396 12458
rect 7536 12412 7566 12458
rect 6998 12393 7566 12412
rect 7670 12427 7790 12585
rect 6550 12362 6670 12381
rect 7670 12381 7689 12427
rect 7735 12381 7790 12427
rect 8118 12477 8238 12585
rect 8342 12477 8462 12585
rect 8566 12477 8686 12585
rect 8118 12458 8686 12477
rect 8118 12412 8516 12458
rect 8656 12412 8686 12458
rect 8118 12393 8686 12412
rect 8790 12427 8910 12585
rect 7670 12362 7790 12381
rect 8790 12381 8809 12427
rect 8855 12381 8910 12427
rect 9238 12477 9358 12585
rect 9462 12477 9582 12585
rect 9686 12477 9806 12585
rect 9238 12458 9806 12477
rect 9238 12412 9636 12458
rect 9776 12412 9806 12458
rect 9238 12393 9806 12412
rect 9910 12427 10030 12585
rect 8790 12362 8910 12381
rect 9910 12381 9929 12427
rect 9975 12381 10030 12427
rect 10358 12477 10478 12585
rect 10582 12477 10702 12585
rect 10806 12477 10926 12585
rect 10358 12458 10926 12477
rect 10358 12412 10756 12458
rect 10896 12412 10926 12458
rect 10358 12393 10926 12412
rect 11030 12427 11150 12585
rect 9910 12362 10030 12381
rect 11030 12381 11049 12427
rect 11095 12381 11150 12427
rect 11478 12477 11598 12585
rect 11702 12477 11822 12585
rect 11926 12477 12046 12585
rect 11478 12458 12046 12477
rect 11478 12412 11876 12458
rect 12016 12412 12046 12458
rect 11478 12393 12046 12412
rect 12150 12427 12270 12585
rect 11030 12362 11150 12381
rect 12150 12381 12169 12427
rect 12215 12381 12270 12427
rect 12598 12477 12718 12585
rect 12822 12477 12942 12585
rect 13046 12477 13166 12585
rect 12598 12458 13166 12477
rect 12598 12412 12996 12458
rect 13136 12412 13166 12458
rect 12598 12393 13166 12412
rect 13270 12427 13390 12585
rect 12150 12362 12270 12381
rect 13270 12381 13289 12427
rect 13335 12381 13390 12427
rect 13718 12477 13838 12585
rect 13942 12477 14062 12585
rect 14166 12477 14286 12585
rect 13718 12458 14286 12477
rect 13718 12412 14116 12458
rect 14256 12412 14286 12458
rect 13718 12393 14286 12412
rect 14390 12427 14510 12585
rect 13270 12362 13390 12381
rect 14390 12381 14409 12427
rect 14455 12381 14510 12427
rect 14838 12477 14958 12585
rect 15062 12477 15182 12585
rect 15286 12477 15406 12585
rect 14838 12458 15406 12477
rect 14838 12412 15236 12458
rect 15376 12412 15406 12458
rect 14838 12393 15406 12412
rect 15510 12427 15630 12585
rect 14390 12362 14510 12381
rect 15510 12381 15529 12427
rect 15575 12381 15630 12427
rect 15958 12477 16078 12585
rect 16182 12477 16302 12585
rect 16406 12477 16526 12585
rect 15958 12458 16526 12477
rect 15958 12412 16356 12458
rect 16496 12412 16526 12458
rect 15958 12393 16526 12412
rect 16630 12427 16750 12585
rect 15510 12362 15630 12381
rect 16630 12381 16649 12427
rect 16695 12381 16750 12427
rect 17078 12477 17198 12585
rect 17302 12477 17422 12585
rect 17526 12477 17646 12585
rect 17078 12458 17646 12477
rect 17078 12412 17476 12458
rect 17616 12412 17646 12458
rect 17078 12393 17646 12412
rect 17750 12427 17870 12585
rect 16630 12362 16750 12381
rect 17750 12381 17769 12427
rect 17815 12381 17870 12427
rect 18198 12477 18318 12585
rect 18422 12477 18542 12585
rect 18646 12477 18766 12585
rect 18198 12458 18766 12477
rect 18198 12412 18596 12458
rect 18736 12412 18766 12458
rect 18198 12393 18766 12412
rect 18870 12427 18990 12585
rect 17750 12362 17870 12381
rect 18870 12381 18889 12427
rect 18935 12381 18990 12427
rect 19318 12477 19438 12585
rect 19542 12477 19662 12585
rect 19766 12477 19886 12585
rect 19318 12458 19886 12477
rect 19318 12412 19716 12458
rect 19856 12412 19886 12458
rect 19318 12393 19886 12412
rect 18870 12362 18990 12381
rect 2518 11947 3086 11966
rect 2070 11905 2190 11924
rect 2070 11859 2089 11905
rect 2135 11859 2190 11905
rect 2070 11770 2190 11859
rect 2518 11901 2916 11947
rect 3056 11901 3086 11947
rect 3638 11947 4206 11966
rect 2518 11849 3086 11901
rect 2518 11770 2638 11849
rect 2742 11770 2862 11849
rect 2966 11770 3086 11849
rect 3190 11905 3310 11924
rect 3190 11859 3209 11905
rect 3255 11859 3310 11905
rect 3190 11770 3310 11859
rect 3638 11901 4036 11947
rect 4176 11901 4206 11947
rect 4758 11947 5326 11966
rect 3638 11849 4206 11901
rect 3638 11770 3758 11849
rect 3862 11770 3982 11849
rect 4086 11770 4206 11849
rect 4310 11905 4430 11924
rect 4310 11859 4329 11905
rect 4375 11859 4430 11905
rect 4310 11770 4430 11859
rect 4758 11901 5156 11947
rect 5296 11901 5326 11947
rect 5878 11947 6446 11966
rect 4758 11849 5326 11901
rect 4758 11770 4878 11849
rect 4982 11770 5102 11849
rect 5206 11770 5326 11849
rect 5430 11905 5550 11924
rect 5430 11859 5449 11905
rect 5495 11859 5550 11905
rect 5430 11770 5550 11859
rect 5878 11901 6276 11947
rect 6416 11901 6446 11947
rect 6998 11947 7566 11966
rect 5878 11849 6446 11901
rect 5878 11770 5998 11849
rect 6102 11770 6222 11849
rect 6326 11770 6446 11849
rect 6550 11905 6670 11924
rect 6550 11859 6569 11905
rect 6615 11859 6670 11905
rect 6550 11770 6670 11859
rect 6998 11901 7396 11947
rect 7536 11901 7566 11947
rect 8118 11947 8686 11966
rect 6998 11849 7566 11901
rect 6998 11770 7118 11849
rect 7222 11770 7342 11849
rect 7446 11770 7566 11849
rect 7670 11905 7790 11924
rect 7670 11859 7689 11905
rect 7735 11859 7790 11905
rect 7670 11770 7790 11859
rect 8118 11901 8516 11947
rect 8656 11901 8686 11947
rect 9238 11947 9806 11966
rect 8118 11849 8686 11901
rect 8118 11770 8238 11849
rect 8342 11770 8462 11849
rect 8566 11770 8686 11849
rect 8790 11905 8910 11924
rect 8790 11859 8809 11905
rect 8855 11859 8910 11905
rect 8790 11770 8910 11859
rect 9238 11901 9636 11947
rect 9776 11901 9806 11947
rect 10358 11947 10926 11966
rect 9238 11849 9806 11901
rect 9238 11770 9358 11849
rect 9462 11770 9582 11849
rect 9686 11770 9806 11849
rect 9910 11905 10030 11924
rect 9910 11859 9929 11905
rect 9975 11859 10030 11905
rect 9910 11770 10030 11859
rect 10358 11901 10756 11947
rect 10896 11901 10926 11947
rect 11478 11947 12046 11966
rect 10358 11849 10926 11901
rect 10358 11770 10478 11849
rect 10582 11770 10702 11849
rect 10806 11770 10926 11849
rect 11030 11905 11150 11924
rect 11030 11859 11049 11905
rect 11095 11859 11150 11905
rect 11030 11770 11150 11859
rect 11478 11901 11876 11947
rect 12016 11901 12046 11947
rect 12598 11947 13166 11966
rect 11478 11849 12046 11901
rect 11478 11770 11598 11849
rect 11702 11770 11822 11849
rect 11926 11770 12046 11849
rect 12150 11905 12270 11924
rect 12150 11859 12169 11905
rect 12215 11859 12270 11905
rect 12150 11770 12270 11859
rect 12598 11901 12996 11947
rect 13136 11901 13166 11947
rect 13718 11947 14286 11966
rect 12598 11849 13166 11901
rect 12598 11770 12718 11849
rect 12822 11770 12942 11849
rect 13046 11770 13166 11849
rect 13270 11905 13390 11924
rect 13270 11859 13289 11905
rect 13335 11859 13390 11905
rect 13270 11770 13390 11859
rect 13718 11901 14116 11947
rect 14256 11901 14286 11947
rect 14838 11947 15406 11966
rect 13718 11849 14286 11901
rect 13718 11770 13838 11849
rect 13942 11770 14062 11849
rect 14166 11770 14286 11849
rect 14390 11905 14510 11924
rect 14390 11859 14409 11905
rect 14455 11859 14510 11905
rect 14390 11770 14510 11859
rect 14838 11901 15236 11947
rect 15376 11901 15406 11947
rect 15958 11947 16526 11966
rect 14838 11849 15406 11901
rect 14838 11770 14958 11849
rect 15062 11770 15182 11849
rect 15286 11770 15406 11849
rect 15510 11905 15630 11924
rect 15510 11859 15529 11905
rect 15575 11859 15630 11905
rect 15510 11770 15630 11859
rect 15958 11901 16356 11947
rect 16496 11901 16526 11947
rect 17078 11947 17646 11966
rect 15958 11849 16526 11901
rect 15958 11770 16078 11849
rect 16182 11770 16302 11849
rect 16406 11770 16526 11849
rect 16630 11905 16750 11924
rect 16630 11859 16649 11905
rect 16695 11859 16750 11905
rect 16630 11770 16750 11859
rect 17078 11901 17476 11947
rect 17616 11901 17646 11947
rect 18198 11947 18766 11966
rect 17078 11849 17646 11901
rect 17078 11770 17198 11849
rect 17302 11770 17422 11849
rect 17526 11770 17646 11849
rect 17750 11905 17870 11924
rect 17750 11859 17769 11905
rect 17815 11859 17870 11905
rect 17750 11770 17870 11859
rect 18198 11901 18596 11947
rect 18736 11901 18766 11947
rect 19318 11947 19886 11966
rect 18198 11849 18766 11901
rect 18198 11770 18318 11849
rect 18422 11770 18542 11849
rect 18646 11770 18766 11849
rect 18870 11905 18990 11924
rect 18870 11859 18889 11905
rect 18935 11859 18990 11905
rect 18870 11770 18990 11859
rect 19318 11901 19716 11947
rect 19856 11901 19886 11947
rect 19318 11849 19886 11901
rect 19318 11770 19438 11849
rect 19542 11770 19662 11849
rect 19766 11770 19886 11849
rect 2070 9910 2190 9954
rect 2518 9910 2638 9954
rect 2742 9910 2862 9954
rect 2966 9910 3086 9954
rect 3190 9910 3310 9954
rect 3638 9910 3758 9954
rect 3862 9910 3982 9954
rect 4086 9910 4206 9954
rect 4310 9910 4430 9954
rect 4758 9910 4878 9954
rect 4982 9910 5102 9954
rect 5206 9910 5326 9954
rect 5430 9910 5550 9954
rect 5878 9910 5998 9954
rect 6102 9910 6222 9954
rect 6326 9910 6446 9954
rect 6550 9910 6670 9954
rect 6998 9910 7118 9954
rect 7222 9910 7342 9954
rect 7446 9910 7566 9954
rect 7670 9910 7790 9954
rect 8118 9910 8238 9954
rect 8342 9910 8462 9954
rect 8566 9910 8686 9954
rect 8790 9910 8910 9954
rect 9238 9910 9358 9954
rect 9462 9910 9582 9954
rect 9686 9910 9806 9954
rect 9910 9910 10030 9954
rect 10358 9910 10478 9954
rect 10582 9910 10702 9954
rect 10806 9910 10926 9954
rect 11030 9910 11150 9954
rect 11478 9910 11598 9954
rect 11702 9910 11822 9954
rect 11926 9910 12046 9954
rect 12150 9910 12270 9954
rect 12598 9910 12718 9954
rect 12822 9910 12942 9954
rect 13046 9910 13166 9954
rect 13270 9910 13390 9954
rect 13718 9910 13838 9954
rect 13942 9910 14062 9954
rect 14166 9910 14286 9954
rect 14390 9910 14510 9954
rect 14838 9910 14958 9954
rect 15062 9910 15182 9954
rect 15286 9910 15406 9954
rect 15510 9910 15630 9954
rect 15958 9910 16078 9954
rect 16182 9910 16302 9954
rect 16406 9910 16526 9954
rect 16630 9910 16750 9954
rect 17078 9910 17198 9954
rect 17302 9910 17422 9954
rect 17526 9910 17646 9954
rect 17750 9910 17870 9954
rect 18198 9910 18318 9954
rect 18422 9910 18542 9954
rect 18646 9910 18766 9954
rect 18870 9910 18990 9954
rect 19318 9910 19438 9954
rect 19542 9910 19662 9954
rect 19766 9910 19886 9954
rect 2697 9209 2815 9237
rect 3211 9209 3329 9237
rect 4388 9209 4506 9237
rect 4902 9209 5020 9237
rect 6079 9209 6197 9237
rect 6593 9209 6711 9237
rect 2696 9165 2816 9209
rect 3210 9165 3330 9209
rect 4387 9165 4507 9209
rect 4901 9165 5021 9209
rect 6078 9165 6198 9209
rect 6592 9165 6712 9209
rect 7525 9021 7645 9094
rect 7749 9021 7869 9094
rect 7973 9021 8093 9094
rect 8197 9021 8317 9094
rect 8421 9021 8541 9094
rect 8645 9021 8765 9094
rect 9158 9021 9278 9094
rect 9382 9021 9502 9094
rect 9606 9021 9726 9094
rect 9830 9021 9950 9094
rect 10054 9021 10174 9094
rect 10278 9021 10398 9094
rect 10792 9021 10912 9094
rect 11016 9021 11136 9094
rect 11240 9021 11360 9094
rect 11464 9021 11584 9094
rect 11688 9021 11808 9094
rect 11912 9021 12032 9094
rect 12426 9021 12546 9094
rect 12650 9021 12770 9094
rect 12874 9021 12994 9094
rect 13098 9021 13218 9094
rect 13322 9021 13442 9094
rect 13546 9021 13666 9094
rect 7525 8495 7645 8567
rect 7749 8495 7869 8567
rect 7973 8495 8093 8567
rect 7525 8358 8093 8495
rect 7525 8286 7645 8358
rect 7749 8286 7869 8358
rect 7973 8286 8093 8358
rect 8197 8495 8317 8567
rect 8421 8495 8541 8567
rect 8645 8495 8765 8567
rect 8197 8358 8765 8495
rect 8197 8286 8317 8358
rect 8421 8286 8541 8358
rect 8645 8286 8765 8358
rect 9158 8495 9278 8567
rect 9382 8495 9502 8567
rect 9606 8495 9726 8567
rect 9158 8358 9726 8495
rect 9158 8286 9278 8358
rect 9382 8286 9502 8358
rect 9606 8286 9726 8358
rect 9830 8495 9950 8567
rect 10054 8495 10174 8567
rect 10278 8495 10398 8567
rect 9830 8358 10398 8495
rect 9830 8286 9950 8358
rect 10054 8286 10174 8358
rect 10278 8286 10398 8358
rect 10792 8495 10912 8567
rect 11016 8495 11136 8567
rect 11240 8495 11360 8567
rect 10792 8358 11360 8495
rect 10792 8286 10912 8358
rect 11016 8286 11136 8358
rect 11240 8286 11360 8358
rect 11464 8495 11584 8567
rect 11688 8495 11808 8567
rect 11912 8495 12032 8567
rect 11464 8358 12032 8495
rect 11464 8286 11584 8358
rect 11688 8286 11808 8358
rect 11912 8286 12032 8358
rect 12426 8495 12546 8567
rect 12650 8495 12770 8567
rect 12874 8495 12994 8567
rect 12426 8358 12994 8495
rect 12426 8286 12546 8358
rect 12650 8286 12770 8358
rect 12874 8286 12994 8358
rect 13098 8495 13218 8567
rect 13322 8495 13442 8567
rect 13546 8495 13666 8567
rect 13098 8358 13666 8495
rect 13098 8286 13218 8358
rect 13322 8286 13442 8358
rect 13546 8286 13666 8358
rect 2696 8213 2816 8257
rect 3210 8213 3330 8257
rect 4387 8213 4507 8257
rect 4901 8213 5021 8257
rect 6078 8213 6198 8257
rect 6592 8213 6712 8257
rect 2696 8185 2815 8213
rect 3210 8185 3329 8213
rect 4387 8185 4506 8213
rect 4901 8185 5020 8213
rect 6078 8185 6197 8213
rect 6592 8185 6711 8213
rect 2410 8139 2815 8185
rect 2410 8093 2484 8139
rect 2530 8093 2642 8139
rect 2688 8093 2815 8139
rect 2410 8047 2815 8093
rect 2920 8139 3329 8185
rect 2920 8093 2994 8139
rect 3040 8093 3152 8139
rect 3198 8093 3329 8139
rect 2920 8047 3329 8093
rect 4101 8139 4506 8185
rect 4101 8093 4175 8139
rect 4221 8093 4333 8139
rect 4379 8093 4506 8139
rect 4101 8047 4506 8093
rect 4611 8139 5020 8185
rect 4611 8093 4685 8139
rect 4731 8093 4843 8139
rect 4889 8093 5020 8139
rect 4611 8047 5020 8093
rect 5792 8139 6197 8185
rect 5792 8093 5866 8139
rect 5912 8093 6024 8139
rect 6070 8093 6197 8139
rect 5792 8047 6197 8093
rect 6302 8139 6711 8185
rect 6302 8093 6376 8139
rect 6422 8093 6534 8139
rect 6580 8093 6711 8139
rect 6302 8047 6711 8093
rect 2696 8021 2815 8047
rect 3210 8021 3329 8047
rect 4387 8021 4506 8047
rect 4901 8021 5020 8047
rect 6078 8021 6197 8047
rect 6592 8021 6711 8047
rect 2696 7977 2816 8021
rect 3210 7977 3330 8021
rect 4387 7977 4507 8021
rect 4901 7977 5021 8021
rect 6078 7977 6198 8021
rect 6592 7977 6712 8021
rect 7525 7063 7645 7132
rect 7749 7063 7869 7132
rect 7973 7063 8093 7132
rect 7525 7044 8093 7063
rect 7525 6998 7678 7044
rect 7912 6998 8093 7044
rect 7525 6979 8093 6998
rect 8197 7063 8317 7132
rect 8421 7063 8541 7132
rect 8645 7063 8765 7132
rect 8197 7044 8765 7063
rect 8197 6998 8378 7044
rect 8612 6998 8765 7044
rect 8197 6979 8765 6998
rect 9158 7063 9278 7132
rect 9382 7063 9502 7132
rect 9606 7063 9726 7132
rect 9158 7044 9726 7063
rect 9158 6998 9311 7044
rect 9545 6998 9726 7044
rect 9158 6979 9726 6998
rect 9830 7063 9950 7132
rect 10054 7063 10174 7132
rect 10278 7063 10398 7132
rect 9830 7044 10398 7063
rect 9830 6998 10011 7044
rect 10245 6998 10398 7044
rect 9830 6979 10398 6998
rect 10792 7063 10912 7132
rect 11016 7063 11136 7132
rect 11240 7063 11360 7132
rect 10792 7044 11360 7063
rect 10792 6998 10945 7044
rect 11179 6998 11360 7044
rect 10792 6979 11360 6998
rect 11464 7063 11584 7132
rect 11688 7063 11808 7132
rect 11912 7063 12032 7132
rect 11464 7044 12032 7063
rect 11464 6998 11645 7044
rect 11879 6998 12032 7044
rect 11464 6979 12032 6998
rect 12426 7063 12546 7132
rect 12650 7063 12770 7132
rect 12874 7063 12994 7132
rect 12426 7044 12994 7063
rect 12426 6998 12579 7044
rect 12813 6998 12994 7044
rect 12426 6979 12994 6998
rect 13098 7063 13218 7132
rect 13322 7063 13442 7132
rect 13546 7063 13666 7132
rect 13098 7044 13666 7063
rect 13098 6998 13279 7044
rect 13513 6998 13666 7044
rect 13098 6979 13666 6998
rect 7525 6419 7645 6491
rect 7749 6419 7869 6491
rect 7973 6419 8093 6491
rect 8197 6419 8317 6491
rect 8421 6419 8541 6491
rect 8645 6419 8765 6491
rect 9158 6419 9278 6491
rect 9382 6419 9502 6491
rect 9606 6419 9726 6491
rect 9830 6419 9950 6491
rect 10054 6419 10174 6491
rect 10278 6419 10398 6491
rect 10792 6419 10912 6491
rect 11016 6419 11136 6491
rect 11240 6419 11360 6491
rect 11464 6419 11584 6491
rect 11688 6419 11808 6491
rect 11912 6419 12032 6491
rect 12426 6419 12546 6491
rect 12650 6419 12770 6491
rect 12874 6419 12994 6491
rect 13098 6419 13218 6491
rect 13322 6419 13442 6491
rect 13546 6419 13666 6491
rect 2696 5211 2816 5255
rect 3210 5211 3330 5255
rect 4387 5211 4507 5255
rect 4901 5211 5021 5255
rect 6078 5211 6198 5255
rect 6592 5211 6712 5255
rect 2696 5181 2815 5211
rect 3210 5181 3329 5211
rect 4387 5181 4506 5211
rect 4901 5181 5020 5211
rect 6078 5181 6197 5211
rect 6592 5181 6711 5211
rect 7525 5182 7645 5285
rect 7488 5137 7681 5182
rect 7488 5091 7562 5137
rect 7608 5091 7681 5137
rect 7488 5045 7681 5091
rect 7526 4578 7645 5045
rect 7749 4983 7869 5285
rect 7973 5211 8093 5285
rect 8197 5211 8317 5285
rect 7712 4938 7905 4983
rect 7712 4892 7786 4938
rect 7832 4892 7905 4938
rect 7712 4846 7905 4892
rect 7526 3912 7646 4578
rect 7748 3912 7868 4846
rect 7974 4780 8092 5211
rect 7973 4779 8092 4780
rect 8198 4780 8316 5211
rect 8421 4983 8541 5285
rect 8645 5182 8765 5285
rect 9158 5182 9278 5285
rect 8608 5137 8801 5182
rect 8608 5091 8682 5137
rect 8728 5091 8801 5137
rect 8608 5045 8801 5091
rect 9121 5137 9314 5182
rect 9121 5091 9195 5137
rect 9241 5091 9314 5137
rect 9121 5045 9314 5091
rect 8384 4938 8577 4983
rect 8384 4892 8458 4938
rect 8504 4892 8577 4938
rect 8384 4846 8577 4892
rect 7936 4734 8129 4779
rect 7936 4688 8010 4734
rect 8056 4688 8129 4734
rect 7936 4642 8129 4688
rect 8198 4642 8317 4780
rect 7972 4175 8092 4642
rect 8198 4175 8318 4642
rect 7972 4037 8093 4175
rect 8197 4174 8318 4175
rect 8160 4129 8353 4174
rect 8160 4083 8234 4129
rect 8280 4083 8353 4129
rect 8160 4037 8353 4083
rect 7972 3912 8092 4037
rect 8198 3912 8318 4037
rect 8422 3912 8542 4846
rect 8645 4578 8764 5045
rect 8644 3912 8764 4578
rect 9159 4578 9278 5045
rect 9382 4933 9502 5285
rect 9606 5211 9726 5285
rect 9830 5211 9950 5285
rect 9381 4846 9502 4933
rect 9159 3912 9279 4578
rect 9381 4375 9501 4846
rect 9607 4780 9725 5211
rect 9606 4779 9725 4780
rect 9831 4780 9949 5211
rect 10054 4933 10174 5285
rect 10278 5182 10398 5285
rect 10241 5137 10434 5182
rect 10241 5091 10315 5137
rect 10361 5091 10434 5137
rect 10241 5045 10434 5091
rect 10792 5080 10912 5285
rect 10054 4846 10175 4933
rect 9569 4734 9762 4779
rect 9569 4688 9643 4734
rect 9689 4688 9762 4734
rect 9569 4642 9762 4688
rect 9831 4642 9950 4780
rect 9345 4330 9538 4375
rect 9345 4284 9419 4330
rect 9465 4284 9538 4330
rect 9345 4238 9538 4284
rect 9381 3912 9501 4238
rect 9605 4175 9725 4642
rect 9831 4175 9951 4642
rect 10055 4375 10175 4846
rect 10278 4578 10397 5045
rect 10017 4330 10210 4375
rect 10017 4284 10091 4330
rect 10137 4284 10210 4330
rect 10017 4238 10210 4284
rect 9605 4037 9726 4175
rect 9830 4174 9951 4175
rect 9793 4129 9986 4174
rect 9793 4083 9867 4129
rect 9913 4083 9986 4129
rect 9793 4037 9986 4083
rect 9605 3912 9725 4037
rect 9831 3912 9951 4037
rect 10055 3912 10175 4238
rect 10277 3912 10397 4578
rect 10793 4578 10912 5080
rect 11016 4983 11136 5285
rect 11240 5211 11360 5285
rect 11464 5211 11584 5285
rect 10979 4938 11172 4983
rect 10979 4892 11053 4938
rect 11099 4892 11172 4938
rect 10979 4846 11172 4892
rect 10793 4577 10913 4578
rect 10755 4532 10948 4577
rect 10755 4486 10829 4532
rect 10875 4486 10948 4532
rect 10755 4440 10948 4486
rect 10793 3912 10913 4440
rect 11015 3912 11135 4846
rect 11241 4780 11359 5211
rect 11240 4779 11359 4780
rect 11465 4780 11583 5211
rect 11688 4983 11808 5285
rect 11912 5080 12032 5285
rect 12426 5080 12546 5285
rect 11651 4938 11844 4983
rect 11651 4892 11725 4938
rect 11771 4892 11844 4938
rect 11651 4846 11844 4892
rect 11203 4734 11396 4779
rect 11203 4688 11277 4734
rect 11323 4688 11396 4734
rect 11203 4642 11396 4688
rect 11465 4642 11584 4780
rect 11239 4175 11359 4642
rect 11465 4175 11585 4642
rect 11239 4037 11360 4175
rect 11464 4174 11585 4175
rect 11427 4129 11620 4174
rect 11427 4083 11501 4129
rect 11547 4083 11620 4129
rect 11427 4037 11620 4083
rect 11239 3912 11359 4037
rect 11465 3912 11585 4037
rect 11689 3912 11809 4846
rect 11912 4578 12031 5080
rect 11911 4577 12031 4578
rect 12427 4578 12546 5080
rect 12650 4933 12770 5285
rect 12874 5211 12994 5285
rect 13098 5211 13218 5285
rect 12649 4846 12770 4933
rect 12427 4577 12547 4578
rect 11875 4532 12068 4577
rect 11875 4486 11949 4532
rect 11995 4486 12068 4532
rect 11875 4440 12068 4486
rect 12389 4532 12582 4577
rect 12389 4486 12463 4532
rect 12509 4486 12582 4532
rect 12389 4440 12582 4486
rect 11911 3912 12031 4440
rect 12427 3912 12547 4440
rect 12649 4375 12769 4846
rect 12875 4780 12993 5211
rect 12874 4779 12993 4780
rect 13099 4780 13217 5211
rect 13322 4933 13442 5285
rect 13546 5080 13666 5285
rect 13322 4846 13443 4933
rect 12837 4734 13030 4779
rect 12837 4688 12911 4734
rect 12957 4688 13030 4734
rect 12837 4642 13030 4688
rect 13099 4642 13218 4780
rect 12613 4330 12806 4375
rect 12613 4284 12687 4330
rect 12733 4284 12806 4330
rect 12613 4238 12806 4284
rect 12649 3912 12769 4238
rect 12873 4175 12993 4642
rect 13099 4175 13219 4642
rect 13323 4375 13443 4846
rect 13546 4578 13665 5080
rect 13545 4577 13665 4578
rect 13509 4532 13702 4577
rect 13509 4486 13583 4532
rect 13629 4486 13702 4532
rect 13509 4440 13702 4486
rect 13285 4330 13478 4375
rect 13285 4284 13359 4330
rect 13405 4284 13478 4330
rect 13285 4238 13478 4284
rect 12873 4037 12994 4175
rect 13098 4174 13219 4175
rect 13061 4129 13254 4174
rect 13061 4083 13135 4129
rect 13181 4083 13254 4129
rect 13061 4037 13254 4083
rect 12873 3912 12993 4037
rect 13099 3912 13219 4037
rect 13323 3912 13443 4238
rect 13545 3912 13665 4440
rect 7526 2477 7646 2550
rect 7748 2477 7868 2550
rect 7972 2477 8092 2550
rect 8198 2477 8318 2550
rect 8422 2477 8542 2550
rect 8644 2477 8764 2550
rect 9159 2477 9279 2550
rect 9381 2477 9501 2550
rect 9605 2477 9725 2550
rect 9831 2477 9951 2550
rect 10055 2477 10175 2550
rect 10277 2477 10397 2550
rect 10793 2477 10913 2550
rect 11015 2477 11135 2550
rect 11239 2477 11359 2550
rect 11465 2477 11585 2550
rect 11689 2477 11809 2550
rect 11911 2477 12031 2550
rect 12427 2477 12547 2550
rect 12649 2477 12769 2550
rect 12873 2477 12993 2550
rect 13099 2477 13219 2550
rect 13323 2477 13443 2550
rect 13545 2477 13665 2550
rect 9283 1944 9403 1988
rect 9507 1944 9627 1988
rect 7913 1829 8033 1873
rect 8990 1771 9127 1790
rect 8990 1631 9009 1771
rect 9055 1631 9127 1771
rect 8990 1612 9127 1631
rect 7913 1318 8033 1557
rect 9060 1502 9127 1612
rect 9283 1502 9403 1562
rect 8735 1432 8956 1451
rect 8735 1386 8754 1432
rect 8800 1386 8956 1432
rect 8735 1367 8956 1386
rect 7807 1243 8151 1318
rect 8836 1282 8956 1367
rect 9060 1436 9403 1502
rect 9507 1467 9627 1562
rect 9507 1451 9801 1467
rect 9508 1448 9801 1451
rect 9060 1380 9404 1436
rect 9060 1282 9180 1380
rect 9284 1282 9404 1380
rect 9508 1402 9642 1448
rect 9782 1402 9801 1448
rect 9508 1383 9801 1402
rect 9508 1282 9628 1383
rect 7807 1183 7927 1243
rect 8031 1183 8151 1243
rect 7807 781 7927 841
rect 8031 781 8151 841
rect 7807 762 8151 781
rect 7807 716 7868 762
rect 8102 716 8151 762
rect 8836 754 8956 827
rect 9060 754 9180 827
rect 9284 754 9404 827
rect 9508 754 9628 827
rect 7807 697 8151 716
<< polycontact >>
rect 6587 27886 6633 28026
rect 5854 27637 5994 27683
rect 6782 27528 6922 27574
rect 13966 27886 14012 28026
rect 13233 27637 13373 27683
rect 7550 26975 7784 27021
rect 1895 25042 2317 25088
rect 2839 25042 3261 25088
rect 3687 25042 4109 25088
rect 5954 25172 6000 25218
rect 6112 25172 6158 25218
rect 6464 25172 6510 25218
rect 6622 25172 6668 25218
rect 7645 25172 7691 25218
rect 7803 25172 7849 25218
rect 8155 25172 8201 25218
rect 8313 25172 8359 25218
rect 14161 27528 14301 27574
rect 24423 27897 24469 28037
rect 23661 27648 23707 27694
rect 23819 27648 23865 27694
rect 24683 27620 24729 27666
rect 14929 26975 15163 27021
rect 25392 26975 25626 27021
rect 4631 25042 5053 25088
rect 1929 21317 1975 21363
rect 2153 20909 2199 20955
rect 3181 21317 3227 21363
rect 2957 20709 3003 20755
rect 3721 21113 3767 21159
rect 3945 20909 3991 20955
rect 9274 25042 9696 25088
rect 10218 25042 10640 25088
rect 11066 25042 11488 25088
rect 13333 25172 13379 25218
rect 13491 25172 13537 25218
rect 13843 25172 13889 25218
rect 14001 25172 14047 25218
rect 15024 25172 15070 25218
rect 15182 25172 15228 25218
rect 15534 25172 15580 25218
rect 15692 25172 15738 25218
rect 12010 25042 12432 25088
rect 9308 21317 9354 21363
rect 4973 21113 5019 21159
rect 4749 20709 4795 20755
rect 9532 20909 9578 20955
rect 10560 21317 10606 21363
rect 10336 20709 10382 20755
rect 11100 21113 11146 21159
rect 11324 20909 11370 20955
rect 23819 25263 23865 25309
rect 23977 25263 24023 25309
rect 24329 25263 24375 25309
rect 24487 25263 24533 25309
rect 25509 25263 25555 25309
rect 25667 25263 25713 25309
rect 26019 25263 26065 25309
rect 26177 25263 26223 25309
rect 27200 25263 27246 25309
rect 27358 25263 27404 25309
rect 27710 25263 27756 25309
rect 27868 25263 27914 25309
rect 16889 24481 17217 24527
rect 17581 24481 17909 24527
rect 18523 24481 18851 24527
rect 19215 24481 19543 24527
rect 20156 24481 20484 24527
rect 20848 24481 21176 24527
rect 21790 24481 22118 24527
rect 22482 24481 22810 24527
rect 16816 21718 16862 21764
rect 12352 21113 12398 21159
rect 12128 20709 12174 20755
rect 17040 21518 17086 21564
rect 17936 21718 17982 21764
rect 18449 21718 18495 21764
rect 17712 21518 17758 21564
rect 17264 21314 17310 21360
rect 17488 20709 17534 20755
rect 18897 21314 18943 21360
rect 18673 20911 18719 20957
rect 19569 21718 19615 21764
rect 19345 20911 19391 20957
rect 19121 20709 19167 20755
rect 20307 21518 20353 21564
rect 20083 21113 20129 21159
rect 20979 21518 21025 21564
rect 20531 21314 20577 21360
rect 20755 20709 20801 20755
rect 21203 21113 21249 21159
rect 21717 21113 21763 21159
rect 22165 21314 22211 21360
rect 21941 20911 21987 20957
rect 22837 21113 22883 21159
rect 22613 20911 22659 20957
rect 22389 20709 22435 20755
rect 2089 12381 2135 12427
rect 2916 12412 3056 12458
rect 3209 12381 3255 12427
rect 4036 12412 4176 12458
rect 4329 12381 4375 12427
rect 5156 12412 5296 12458
rect 5449 12381 5495 12427
rect 6276 12412 6416 12458
rect 6569 12381 6615 12427
rect 7396 12412 7536 12458
rect 7689 12381 7735 12427
rect 8516 12412 8656 12458
rect 8809 12381 8855 12427
rect 9636 12412 9776 12458
rect 9929 12381 9975 12427
rect 10756 12412 10896 12458
rect 11049 12381 11095 12427
rect 11876 12412 12016 12458
rect 12169 12381 12215 12427
rect 12996 12412 13136 12458
rect 13289 12381 13335 12427
rect 14116 12412 14256 12458
rect 14409 12381 14455 12427
rect 15236 12412 15376 12458
rect 15529 12381 15575 12427
rect 16356 12412 16496 12458
rect 16649 12381 16695 12427
rect 17476 12412 17616 12458
rect 17769 12381 17815 12427
rect 18596 12412 18736 12458
rect 18889 12381 18935 12427
rect 19716 12412 19856 12458
rect 2089 11859 2135 11905
rect 2916 11901 3056 11947
rect 3209 11859 3255 11905
rect 4036 11901 4176 11947
rect 4329 11859 4375 11905
rect 5156 11901 5296 11947
rect 5449 11859 5495 11905
rect 6276 11901 6416 11947
rect 6569 11859 6615 11905
rect 7396 11901 7536 11947
rect 7689 11859 7735 11905
rect 8516 11901 8656 11947
rect 8809 11859 8855 11905
rect 9636 11901 9776 11947
rect 9929 11859 9975 11905
rect 10756 11901 10896 11947
rect 11049 11859 11095 11905
rect 11876 11901 12016 11947
rect 12169 11859 12215 11905
rect 12996 11901 13136 11947
rect 13289 11859 13335 11905
rect 14116 11901 14256 11947
rect 14409 11859 14455 11905
rect 15236 11901 15376 11947
rect 15529 11859 15575 11905
rect 16356 11901 16496 11947
rect 16649 11859 16695 11905
rect 17476 11901 17616 11947
rect 17769 11859 17815 11905
rect 18596 11901 18736 11947
rect 18889 11859 18935 11905
rect 19716 11901 19856 11947
rect 2484 8093 2530 8139
rect 2642 8093 2688 8139
rect 2994 8093 3040 8139
rect 3152 8093 3198 8139
rect 4175 8093 4221 8139
rect 4333 8093 4379 8139
rect 4685 8093 4731 8139
rect 4843 8093 4889 8139
rect 5866 8093 5912 8139
rect 6024 8093 6070 8139
rect 6376 8093 6422 8139
rect 6534 8093 6580 8139
rect 7678 6998 7912 7044
rect 8378 6998 8612 7044
rect 9311 6998 9545 7044
rect 10011 6998 10245 7044
rect 10945 6998 11179 7044
rect 11645 6998 11879 7044
rect 12579 6998 12813 7044
rect 13279 6998 13513 7044
rect 7562 5091 7608 5137
rect 7786 4892 7832 4938
rect 8682 5091 8728 5137
rect 9195 5091 9241 5137
rect 8458 4892 8504 4938
rect 8010 4688 8056 4734
rect 8234 4083 8280 4129
rect 10315 5091 10361 5137
rect 9643 4688 9689 4734
rect 9419 4284 9465 4330
rect 10091 4284 10137 4330
rect 9867 4083 9913 4129
rect 11053 4892 11099 4938
rect 10829 4486 10875 4532
rect 11725 4892 11771 4938
rect 11277 4688 11323 4734
rect 11501 4083 11547 4129
rect 11949 4486 11995 4532
rect 12463 4486 12509 4532
rect 12911 4688 12957 4734
rect 12687 4284 12733 4330
rect 13583 4486 13629 4532
rect 13359 4284 13405 4330
rect 13135 4083 13181 4129
rect 9009 1631 9055 1771
rect 8754 1386 8800 1432
rect 9642 1402 9782 1448
rect 7868 716 8102 762
<< metal1 >>
rect 403 28996 537 29037
rect 403 28944 444 28996
rect 496 28944 537 28996
rect 403 28778 537 28944
rect 403 28726 444 28778
rect 496 28726 537 28778
rect 403 1155 537 28726
rect 1624 29007 1740 29016
rect 2072 29007 2188 29016
rect 2520 29007 2636 29016
rect 2968 29007 3084 29016
rect 3416 29007 3532 29016
rect 3864 29007 3980 29016
rect 4312 29007 4428 29016
rect 4760 29007 4876 29016
rect 5208 29007 9119 29016
rect 9451 29007 9567 29016
rect 9899 29007 10015 29016
rect 10347 29007 10463 29016
rect 10795 29007 10911 29016
rect 11243 29007 11359 29016
rect 11691 29007 11807 29016
rect 12139 29007 12255 29016
rect 12587 29007 16497 29016
rect 1624 28996 16497 29007
rect 1624 28950 1772 28996
rect 5202 28980 9132 28996
rect 12562 28980 16497 28996
rect 5202 28950 5401 28980
rect 1624 28939 5401 28950
rect 1624 28640 1740 28939
rect 1624 28594 1659 28640
rect 1705 28594 1740 28640
rect 1624 28540 1740 28594
rect 1883 28640 1929 28653
rect 1618 28535 1746 28540
rect 1618 28500 1659 28535
rect 1705 28500 1746 28535
rect 1618 28448 1656 28500
rect 1708 28448 1746 28500
rect 1618 28430 1746 28448
rect 1618 28384 1659 28430
rect 1705 28384 1746 28430
rect 1618 28325 1746 28384
rect 1618 28282 1659 28325
rect 1705 28282 1746 28325
rect 1618 28230 1656 28282
rect 1708 28230 1746 28282
rect 1618 28220 1746 28230
rect 1618 28174 1659 28220
rect 1705 28174 1746 28220
rect 1618 28116 1746 28174
rect 1618 28070 1659 28116
rect 1705 28070 1746 28116
rect 1618 28064 1746 28070
rect 1618 28012 1656 28064
rect 1708 28012 1746 28064
rect 1618 27966 1659 28012
rect 1705 27966 1746 28012
rect 1618 27908 1746 27966
rect 1618 27862 1659 27908
rect 1705 27862 1746 27908
rect 1618 27846 1746 27862
rect 1618 27794 1656 27846
rect 1708 27794 1746 27846
rect 1883 28535 1929 28594
rect 2072 28640 2188 28939
rect 2072 28594 2107 28640
rect 2153 28594 2188 28640
rect 2072 28540 2188 28594
rect 2331 28640 2377 28653
rect 2331 28540 2377 28594
rect 2520 28640 2636 28939
rect 2520 28594 2555 28640
rect 2601 28594 2636 28640
rect 1883 28430 1929 28489
rect 1883 28325 1929 28384
rect 1883 28220 1929 28279
rect 1883 28116 1929 28174
rect 1883 28012 1929 28070
rect 1883 27908 1929 27966
rect 1883 27804 1929 27862
rect 1618 27758 1659 27794
rect 1705 27758 1746 27794
rect 1618 27754 1746 27758
rect 1848 27758 1883 27795
rect 2058 28539 2188 28540
rect 2058 28535 2186 28539
rect 2058 28500 2107 28535
rect 2058 28448 2096 28500
rect 2153 28489 2186 28535
rect 2148 28448 2186 28489
rect 2058 28430 2186 28448
rect 2058 28384 2107 28430
rect 2153 28384 2186 28430
rect 2058 28325 2186 28384
rect 2058 28282 2107 28325
rect 2058 28230 2096 28282
rect 2153 28279 2186 28325
rect 2148 28230 2186 28279
rect 2058 28220 2186 28230
rect 2058 28174 2107 28220
rect 2153 28174 2186 28220
rect 2058 28116 2186 28174
rect 2058 28070 2107 28116
rect 2153 28070 2186 28116
rect 2058 28064 2186 28070
rect 2058 28012 2096 28064
rect 2148 28012 2186 28064
rect 2058 27966 2107 28012
rect 2153 27966 2186 28012
rect 2058 27908 2186 27966
rect 2058 27862 2107 27908
rect 2153 27862 2186 27908
rect 2058 27846 2186 27862
rect 1929 27758 1964 27795
rect 1659 27745 1705 27754
rect 1848 27665 1964 27758
rect 2058 27794 2096 27846
rect 2148 27804 2186 27846
rect 2058 27758 2107 27794
rect 2153 27758 2186 27804
rect 2058 27754 2186 27758
rect 2290 28535 2418 28540
rect 2520 28539 2636 28594
rect 2779 28640 2825 28653
rect 2779 28540 2825 28594
rect 2968 28640 3084 28939
rect 2968 28594 3003 28640
rect 3049 28594 3084 28640
rect 2968 28540 3084 28594
rect 3227 28640 3273 28653
rect 2290 28500 2331 28535
rect 2377 28500 2418 28535
rect 2290 28448 2328 28500
rect 2380 28448 2418 28500
rect 2290 28430 2418 28448
rect 2290 28384 2331 28430
rect 2377 28384 2418 28430
rect 2290 28325 2418 28384
rect 2290 28282 2331 28325
rect 2377 28282 2418 28325
rect 2290 28230 2328 28282
rect 2380 28230 2418 28282
rect 2290 28220 2418 28230
rect 2290 28174 2331 28220
rect 2377 28174 2418 28220
rect 2290 28116 2418 28174
rect 2290 28070 2331 28116
rect 2377 28070 2418 28116
rect 2290 28064 2418 28070
rect 2290 28012 2328 28064
rect 2380 28012 2418 28064
rect 2290 27966 2331 28012
rect 2377 27966 2418 28012
rect 2290 27908 2418 27966
rect 2290 27862 2331 27908
rect 2377 27862 2418 27908
rect 2290 27846 2418 27862
rect 2290 27794 2328 27846
rect 2380 27794 2418 27846
rect 2290 27758 2331 27794
rect 2377 27758 2418 27794
rect 2290 27754 2418 27758
rect 2555 28535 2601 28539
rect 2555 28430 2601 28489
rect 2555 28325 2601 28384
rect 2555 28220 2601 28279
rect 2555 28116 2601 28174
rect 2555 28012 2601 28070
rect 2555 27908 2601 27966
rect 2555 27804 2601 27862
rect 2107 27745 2153 27754
rect 2296 27665 2412 27754
rect 2555 27745 2601 27758
rect 2738 28535 2866 28540
rect 2968 28539 3098 28540
rect 2738 28500 2779 28535
rect 2825 28500 2866 28535
rect 2738 28448 2776 28500
rect 2828 28448 2866 28500
rect 2738 28430 2866 28448
rect 2738 28384 2779 28430
rect 2825 28384 2866 28430
rect 2738 28325 2866 28384
rect 2738 28282 2779 28325
rect 2825 28282 2866 28325
rect 2738 28230 2776 28282
rect 2828 28230 2866 28282
rect 2738 28220 2866 28230
rect 2738 28174 2779 28220
rect 2825 28174 2866 28220
rect 2738 28116 2866 28174
rect 2738 28070 2779 28116
rect 2825 28070 2866 28116
rect 2738 28064 2866 28070
rect 2738 28012 2776 28064
rect 2828 28012 2866 28064
rect 2738 27966 2779 28012
rect 2825 27966 2866 28012
rect 2738 27908 2866 27966
rect 2738 27862 2779 27908
rect 2825 27862 2866 27908
rect 2738 27846 2866 27862
rect 2738 27794 2776 27846
rect 2828 27794 2866 27846
rect 2738 27758 2779 27794
rect 2825 27758 2866 27794
rect 2738 27754 2866 27758
rect 2970 28535 3098 28539
rect 2970 28489 3003 28535
rect 3049 28500 3098 28535
rect 2970 28448 3008 28489
rect 3060 28448 3098 28500
rect 2970 28430 3098 28448
rect 2970 28384 3003 28430
rect 3049 28384 3098 28430
rect 2970 28325 3098 28384
rect 2970 28279 3003 28325
rect 3049 28282 3098 28325
rect 2970 28230 3008 28279
rect 3060 28230 3098 28282
rect 2970 28220 3098 28230
rect 2970 28174 3003 28220
rect 3049 28174 3098 28220
rect 2970 28116 3098 28174
rect 2970 28070 3003 28116
rect 3049 28070 3098 28116
rect 2970 28064 3098 28070
rect 2970 28012 3008 28064
rect 3060 28012 3098 28064
rect 2970 27966 3003 28012
rect 3049 27966 3098 28012
rect 2970 27908 3098 27966
rect 2970 27862 3003 27908
rect 3049 27862 3098 27908
rect 2970 27846 3098 27862
rect 2970 27804 3008 27846
rect 2970 27758 3003 27804
rect 3060 27794 3098 27846
rect 3227 28535 3273 28594
rect 3416 28640 3532 28939
rect 3416 28594 3451 28640
rect 3497 28594 3532 28640
rect 3416 28540 3532 28594
rect 3675 28640 3721 28653
rect 3227 28430 3273 28489
rect 3227 28325 3273 28384
rect 3227 28220 3273 28279
rect 3227 28116 3273 28174
rect 3227 28012 3273 28070
rect 3227 27908 3273 27966
rect 3227 27804 3273 27862
rect 3049 27758 3098 27794
rect 2970 27754 3098 27758
rect 3192 27758 3227 27795
rect 3410 28535 3538 28540
rect 3410 28500 3451 28535
rect 3497 28500 3538 28535
rect 3410 28448 3448 28500
rect 3500 28448 3538 28500
rect 3410 28430 3538 28448
rect 3410 28384 3451 28430
rect 3497 28384 3538 28430
rect 3410 28325 3538 28384
rect 3410 28282 3451 28325
rect 3497 28282 3538 28325
rect 3410 28230 3448 28282
rect 3500 28230 3538 28282
rect 3410 28220 3538 28230
rect 3410 28174 3451 28220
rect 3497 28174 3538 28220
rect 3410 28116 3538 28174
rect 3410 28070 3451 28116
rect 3497 28070 3538 28116
rect 3410 28064 3538 28070
rect 3410 28012 3448 28064
rect 3500 28012 3538 28064
rect 3410 27966 3451 28012
rect 3497 27966 3538 28012
rect 3410 27908 3538 27966
rect 3410 27862 3451 27908
rect 3497 27862 3538 27908
rect 3410 27846 3538 27862
rect 3273 27758 3308 27795
rect 1848 27546 2412 27665
rect 1659 27452 1705 27465
rect 1659 27392 1705 27406
rect 1848 27452 1964 27546
rect 1848 27406 1883 27452
rect 1929 27406 1964 27452
rect 1848 27396 1964 27406
rect 2107 27452 2153 27465
rect 1618 27353 1746 27392
rect 1618 27301 1656 27353
rect 1708 27301 1746 27353
rect 1618 27242 1746 27301
rect 1618 27196 1659 27242
rect 1705 27196 1746 27242
rect 1618 27137 1746 27196
rect 1618 27135 1659 27137
rect 1705 27135 1746 27137
rect 1618 27083 1656 27135
rect 1708 27083 1746 27135
rect 1618 27032 1746 27083
rect 1618 26986 1659 27032
rect 1705 26986 1746 27032
rect 1618 26927 1746 26986
rect 1618 26917 1659 26927
rect 1705 26917 1746 26927
rect 1618 26865 1656 26917
rect 1708 26865 1746 26917
rect 1618 26825 1746 26865
rect 1883 27347 1929 27396
rect 2107 27392 2153 27406
rect 2296 27452 2412 27546
rect 2744 27665 2860 27754
rect 3003 27745 3049 27754
rect 3192 27665 3308 27758
rect 3410 27794 3448 27846
rect 3500 27794 3538 27846
rect 3675 28535 3721 28594
rect 3864 28640 3980 28939
rect 3864 28594 3899 28640
rect 3945 28594 3980 28640
rect 3864 28540 3980 28594
rect 4123 28640 4169 28653
rect 4123 28540 4169 28594
rect 4312 28640 4428 28939
rect 4312 28594 4347 28640
rect 4393 28594 4428 28640
rect 3675 28430 3721 28489
rect 3675 28325 3721 28384
rect 3675 28220 3721 28279
rect 3675 28116 3721 28174
rect 3675 28012 3721 28070
rect 3675 27908 3721 27966
rect 3675 27804 3721 27862
rect 3410 27758 3451 27794
rect 3497 27758 3538 27794
rect 3410 27754 3538 27758
rect 3640 27758 3675 27795
rect 3850 28539 3980 28540
rect 3850 28535 3978 28539
rect 3850 28500 3899 28535
rect 3850 28448 3888 28500
rect 3945 28489 3978 28535
rect 3940 28448 3978 28489
rect 3850 28430 3978 28448
rect 3850 28384 3899 28430
rect 3945 28384 3978 28430
rect 3850 28325 3978 28384
rect 3850 28282 3899 28325
rect 3850 28230 3888 28282
rect 3945 28279 3978 28325
rect 3940 28230 3978 28279
rect 3850 28220 3978 28230
rect 3850 28174 3899 28220
rect 3945 28174 3978 28220
rect 3850 28116 3978 28174
rect 3850 28070 3899 28116
rect 3945 28070 3978 28116
rect 3850 28064 3978 28070
rect 3850 28012 3888 28064
rect 3940 28012 3978 28064
rect 3850 27966 3899 28012
rect 3945 27966 3978 28012
rect 3850 27908 3978 27966
rect 3850 27862 3899 27908
rect 3945 27862 3978 27908
rect 3850 27846 3978 27862
rect 3721 27758 3756 27795
rect 3451 27745 3497 27754
rect 2744 27546 3308 27665
rect 2296 27406 2331 27452
rect 2377 27406 2412 27452
rect 2296 27396 2412 27406
rect 2555 27452 2601 27465
rect 1883 27242 1929 27301
rect 1883 27137 1929 27196
rect 1883 27032 1929 27091
rect 1883 26927 1929 26986
rect 1659 26822 1705 26825
rect 1659 26717 1705 26776
rect 1659 26612 1705 26671
rect 1659 26507 1705 26566
rect 1659 26402 1705 26461
rect 1659 26297 1705 26356
rect 1659 26192 1705 26251
rect 1659 26088 1705 26146
rect 1659 25984 1705 26042
rect 1659 25880 1705 25938
rect 1659 25776 1705 25834
rect 1659 25672 1705 25730
rect 1659 25568 1705 25626
rect 1659 25464 1705 25522
rect 1659 25360 1705 25418
rect 1659 25256 1705 25314
rect 1659 25197 1705 25210
rect 1883 26822 1929 26881
rect 2066 27353 2194 27392
rect 2066 27301 2104 27353
rect 2156 27301 2194 27353
rect 2066 27242 2194 27301
rect 2066 27196 2107 27242
rect 2153 27196 2194 27242
rect 2066 27137 2194 27196
rect 2066 27135 2107 27137
rect 2153 27135 2194 27137
rect 2066 27083 2104 27135
rect 2156 27083 2194 27135
rect 2066 27032 2194 27083
rect 2066 26986 2107 27032
rect 2153 26986 2194 27032
rect 2066 26927 2194 26986
rect 2066 26917 2107 26927
rect 2153 26917 2194 26927
rect 2066 26865 2104 26917
rect 2156 26865 2194 26917
rect 2066 26825 2194 26865
rect 2331 27347 2377 27396
rect 2555 27392 2601 27406
rect 2744 27452 2860 27546
rect 2744 27406 2779 27452
rect 2825 27406 2860 27452
rect 2744 27396 2860 27406
rect 3003 27452 3049 27465
rect 2331 27242 2377 27301
rect 2331 27137 2377 27196
rect 2331 27032 2377 27091
rect 2331 26927 2377 26986
rect 1883 26717 1929 26776
rect 1883 26612 1929 26671
rect 1883 26507 1929 26566
rect 1883 26402 1929 26461
rect 1883 26297 1929 26356
rect 1883 26192 1929 26251
rect 1883 26088 1929 26146
rect 1883 25984 1929 26042
rect 1883 25880 1929 25938
rect 1883 25776 1929 25834
rect 1883 25672 1929 25730
rect 1883 25568 1929 25626
rect 1883 25464 1929 25522
rect 1883 25360 1929 25418
rect 1883 25256 1929 25314
rect 1883 25197 1929 25210
rect 2107 26822 2153 26825
rect 2107 26717 2153 26776
rect 2107 26612 2153 26671
rect 2107 26507 2153 26566
rect 2107 26402 2153 26461
rect 2107 26297 2153 26356
rect 2107 26192 2153 26251
rect 2107 26088 2153 26146
rect 2107 25984 2153 26042
rect 2107 25880 2153 25938
rect 2107 25776 2153 25834
rect 2107 25672 2153 25730
rect 2107 25568 2153 25626
rect 2107 25464 2153 25522
rect 2107 25360 2153 25418
rect 2107 25256 2153 25314
rect 2107 25197 2153 25210
rect 2331 26822 2377 26881
rect 2514 27353 2642 27392
rect 2514 27301 2552 27353
rect 2604 27301 2642 27353
rect 2514 27242 2642 27301
rect 2514 27196 2555 27242
rect 2601 27196 2642 27242
rect 2514 27137 2642 27196
rect 2514 27135 2555 27137
rect 2601 27135 2642 27137
rect 2514 27083 2552 27135
rect 2604 27083 2642 27135
rect 2514 27032 2642 27083
rect 2514 26986 2555 27032
rect 2601 26986 2642 27032
rect 2514 26927 2642 26986
rect 2514 26917 2555 26927
rect 2601 26917 2642 26927
rect 2514 26865 2552 26917
rect 2604 26865 2642 26917
rect 2514 26825 2642 26865
rect 2779 27347 2825 27396
rect 3003 27392 3049 27406
rect 3192 27452 3308 27546
rect 3640 27665 3756 27758
rect 3850 27794 3888 27846
rect 3940 27804 3978 27846
rect 3850 27758 3899 27794
rect 3945 27758 3978 27804
rect 3850 27754 3978 27758
rect 4082 28535 4210 28540
rect 4312 28539 4428 28594
rect 4571 28640 4617 28653
rect 4571 28540 4617 28594
rect 4760 28640 4876 28939
rect 5208 28934 5401 28939
rect 5447 28934 5559 28980
rect 5605 28934 5717 28980
rect 5763 28934 5875 28980
rect 5921 28934 6033 28980
rect 6079 28934 6191 28980
rect 6237 28934 6349 28980
rect 6395 28934 6507 28980
rect 6553 28934 6666 28980
rect 6712 28934 6824 28980
rect 6870 28934 6982 28980
rect 7028 28934 7140 28980
rect 7186 28934 7298 28980
rect 7344 28934 7456 28980
rect 7502 28934 7614 28980
rect 7660 28934 7773 28980
rect 7819 28934 7931 28980
rect 7977 28934 8089 28980
rect 8135 28934 8247 28980
rect 8293 28934 8405 28980
rect 8451 28934 8563 28980
rect 8609 28934 8721 28980
rect 8767 28934 8879 28980
rect 8925 28934 9037 28980
rect 12562 28950 12780 28980
rect 9083 28939 12780 28950
rect 9083 28934 9119 28939
rect 5208 28897 9119 28934
rect 4760 28594 4795 28640
rect 4841 28594 4876 28640
rect 4760 28540 4876 28594
rect 5019 28640 5065 28653
rect 4082 28500 4123 28535
rect 4169 28500 4210 28535
rect 4082 28448 4120 28500
rect 4172 28448 4210 28500
rect 4082 28430 4210 28448
rect 4082 28384 4123 28430
rect 4169 28384 4210 28430
rect 4082 28325 4210 28384
rect 4082 28282 4123 28325
rect 4169 28282 4210 28325
rect 4082 28230 4120 28282
rect 4172 28230 4210 28282
rect 4082 28220 4210 28230
rect 4082 28174 4123 28220
rect 4169 28174 4210 28220
rect 4082 28116 4210 28174
rect 4082 28070 4123 28116
rect 4169 28070 4210 28116
rect 4082 28064 4210 28070
rect 4082 28012 4120 28064
rect 4172 28012 4210 28064
rect 4082 27966 4123 28012
rect 4169 27966 4210 28012
rect 4082 27908 4210 27966
rect 4082 27862 4123 27908
rect 4169 27862 4210 27908
rect 4082 27846 4210 27862
rect 4082 27794 4120 27846
rect 4172 27794 4210 27846
rect 4082 27758 4123 27794
rect 4169 27758 4210 27794
rect 4082 27754 4210 27758
rect 4347 28535 4393 28539
rect 4347 28430 4393 28489
rect 4347 28325 4393 28384
rect 4347 28220 4393 28279
rect 4347 28116 4393 28174
rect 4347 28012 4393 28070
rect 4347 27908 4393 27966
rect 4347 27804 4393 27862
rect 3899 27745 3945 27754
rect 4088 27665 4204 27754
rect 4347 27745 4393 27758
rect 4530 28535 4658 28540
rect 4760 28539 4890 28540
rect 4530 28500 4571 28535
rect 4617 28500 4658 28535
rect 4530 28448 4568 28500
rect 4620 28448 4658 28500
rect 4530 28430 4658 28448
rect 4530 28384 4571 28430
rect 4617 28384 4658 28430
rect 4530 28325 4658 28384
rect 4530 28282 4571 28325
rect 4617 28282 4658 28325
rect 4530 28230 4568 28282
rect 4620 28230 4658 28282
rect 4530 28220 4658 28230
rect 4530 28174 4571 28220
rect 4617 28174 4658 28220
rect 4530 28116 4658 28174
rect 4530 28070 4571 28116
rect 4617 28070 4658 28116
rect 4530 28064 4658 28070
rect 4530 28012 4568 28064
rect 4620 28012 4658 28064
rect 4530 27966 4571 28012
rect 4617 27966 4658 28012
rect 4530 27908 4658 27966
rect 4530 27862 4571 27908
rect 4617 27862 4658 27908
rect 4530 27846 4658 27862
rect 4530 27794 4568 27846
rect 4620 27794 4658 27846
rect 4530 27758 4571 27794
rect 4617 27758 4658 27794
rect 4530 27754 4658 27758
rect 4762 28535 4890 28539
rect 4762 28489 4795 28535
rect 4841 28500 4890 28535
rect 4762 28448 4800 28489
rect 4852 28448 4890 28500
rect 4762 28430 4890 28448
rect 4762 28384 4795 28430
rect 4841 28384 4890 28430
rect 4762 28325 4890 28384
rect 4762 28279 4795 28325
rect 4841 28282 4890 28325
rect 4762 28230 4800 28279
rect 4852 28230 4890 28282
rect 4762 28220 4890 28230
rect 4762 28174 4795 28220
rect 4841 28174 4890 28220
rect 4762 28116 4890 28174
rect 4762 28070 4795 28116
rect 4841 28070 4890 28116
rect 4762 28064 4890 28070
rect 4762 28012 4800 28064
rect 4852 28012 4890 28064
rect 4762 27966 4795 28012
rect 4841 27966 4890 28012
rect 4762 27908 4890 27966
rect 4762 27862 4795 27908
rect 4841 27862 4890 27908
rect 4762 27846 4890 27862
rect 4762 27804 4800 27846
rect 4762 27758 4795 27804
rect 4852 27794 4890 27846
rect 5019 28535 5065 28594
rect 5208 28640 5324 28897
rect 5208 28594 5243 28640
rect 5289 28594 5324 28640
rect 5208 28540 5324 28594
rect 5897 28896 6014 28897
rect 5019 28430 5065 28489
rect 5019 28325 5065 28384
rect 5019 28220 5065 28279
rect 5019 28116 5065 28174
rect 5019 28012 5065 28070
rect 5019 27908 5065 27966
rect 5019 27804 5065 27862
rect 4841 27758 4890 27794
rect 4762 27754 4890 27758
rect 4984 27758 5019 27795
rect 5202 28535 5330 28540
rect 5202 28500 5243 28535
rect 5289 28500 5330 28535
rect 5202 28448 5240 28500
rect 5292 28448 5330 28500
rect 5202 28430 5330 28448
rect 5897 28440 6013 28896
rect 6345 28440 6461 28897
rect 5202 28384 5243 28430
rect 5289 28384 5330 28430
rect 5202 28325 5330 28384
rect 5202 28282 5243 28325
rect 5289 28282 5330 28325
rect 5202 28230 5240 28282
rect 5292 28230 5330 28282
rect 5202 28220 5330 28230
rect 5202 28174 5243 28220
rect 5289 28174 5330 28220
rect 5202 28116 5330 28174
rect 5202 28070 5243 28116
rect 5289 28070 5330 28116
rect 5202 28064 5330 28070
rect 5202 28012 5240 28064
rect 5292 28012 5330 28064
rect 5202 27966 5243 28012
rect 5289 27966 5330 28012
rect 5202 27908 5330 27966
rect 5202 27862 5243 27908
rect 5289 27862 5330 27908
rect 5885 28401 6013 28440
rect 5885 28349 5923 28401
rect 5975 28349 6013 28401
rect 5885 28183 6013 28349
rect 5885 28131 5923 28183
rect 5975 28131 6013 28183
rect 6324 28401 6461 28440
rect 6324 28349 6362 28401
rect 6414 28349 6461 28401
rect 7716 28896 7832 28897
rect 7716 28384 7831 28896
rect 9003 28640 9119 28897
rect 9003 28594 9038 28640
rect 9084 28594 9119 28640
rect 9003 28540 9119 28594
rect 9262 28640 9308 28653
rect 8997 28535 9125 28540
rect 8997 28500 9038 28535
rect 9084 28500 9125 28535
rect 8997 28448 9035 28500
rect 9087 28448 9125 28500
rect 8997 28430 9125 28448
rect 8997 28384 9038 28430
rect 9084 28384 9125 28430
rect 7716 28383 7832 28384
rect 6324 28183 6461 28349
rect 7708 28344 7836 28383
rect 7708 28292 7746 28344
rect 7798 28292 7836 28344
rect 5885 28082 6013 28131
rect 5885 27965 5933 28082
rect 5885 27913 5923 27965
rect 5885 27873 5933 27913
rect 5202 27846 5330 27862
rect 5065 27758 5100 27795
rect 3640 27546 4204 27665
rect 3192 27406 3227 27452
rect 3273 27406 3308 27452
rect 3192 27396 3308 27406
rect 3451 27452 3497 27465
rect 2779 27242 2825 27301
rect 2779 27137 2825 27196
rect 2779 27032 2825 27091
rect 2779 26927 2825 26986
rect 2331 26717 2377 26776
rect 2331 26612 2377 26671
rect 2331 26507 2377 26566
rect 2331 26402 2377 26461
rect 2331 26297 2377 26356
rect 2331 26192 2377 26251
rect 2331 26088 2377 26146
rect 2331 25984 2377 26042
rect 2331 25880 2377 25938
rect 2331 25776 2377 25834
rect 2331 25672 2377 25730
rect 2331 25568 2377 25626
rect 2331 25464 2377 25522
rect 2331 25360 2377 25418
rect 2331 25256 2377 25314
rect 2331 25197 2377 25210
rect 2555 26822 2601 26825
rect 2555 26717 2601 26776
rect 2555 26612 2601 26671
rect 2555 26507 2601 26566
rect 2555 26402 2601 26461
rect 2555 26297 2601 26356
rect 2555 26192 2601 26251
rect 2555 26088 2601 26146
rect 2555 25984 2601 26042
rect 2555 25880 2601 25938
rect 2555 25776 2601 25834
rect 2555 25672 2601 25730
rect 2555 25568 2601 25626
rect 2555 25464 2601 25522
rect 2555 25360 2601 25418
rect 2555 25256 2601 25314
rect 2555 25197 2601 25210
rect 2779 26822 2825 26881
rect 2962 27353 3090 27392
rect 2962 27301 3000 27353
rect 3052 27301 3090 27353
rect 2962 27242 3090 27301
rect 2962 27196 3003 27242
rect 3049 27196 3090 27242
rect 2962 27137 3090 27196
rect 2962 27135 3003 27137
rect 3049 27135 3090 27137
rect 2962 27083 3000 27135
rect 3052 27083 3090 27135
rect 2962 27032 3090 27083
rect 2962 26986 3003 27032
rect 3049 26986 3090 27032
rect 2962 26927 3090 26986
rect 2962 26917 3003 26927
rect 3049 26917 3090 26927
rect 2962 26865 3000 26917
rect 3052 26865 3090 26917
rect 2962 26825 3090 26865
rect 3227 27347 3273 27396
rect 3451 27392 3497 27406
rect 3640 27452 3756 27546
rect 3640 27406 3675 27452
rect 3721 27406 3756 27452
rect 3640 27396 3756 27406
rect 3899 27452 3945 27465
rect 3227 27242 3273 27301
rect 3227 27137 3273 27196
rect 3227 27032 3273 27091
rect 3227 26927 3273 26986
rect 2779 26717 2825 26776
rect 2779 26612 2825 26671
rect 2779 26507 2825 26566
rect 2779 26402 2825 26461
rect 2779 26297 2825 26356
rect 2779 26192 2825 26251
rect 2779 26088 2825 26146
rect 2779 25984 2825 26042
rect 2779 25880 2825 25938
rect 2779 25776 2825 25834
rect 2779 25672 2825 25730
rect 2779 25568 2825 25626
rect 2779 25464 2825 25522
rect 2779 25360 2825 25418
rect 2779 25256 2825 25314
rect 2779 25197 2825 25210
rect 3003 26822 3049 26825
rect 3003 26717 3049 26776
rect 3003 26612 3049 26671
rect 3003 26507 3049 26566
rect 3003 26402 3049 26461
rect 3003 26297 3049 26356
rect 3003 26192 3049 26251
rect 3003 26088 3049 26146
rect 3003 25984 3049 26042
rect 3003 25880 3049 25938
rect 3003 25776 3049 25834
rect 3003 25672 3049 25730
rect 3003 25568 3049 25626
rect 3003 25464 3049 25522
rect 3003 25360 3049 25418
rect 3003 25256 3049 25314
rect 3003 25197 3049 25210
rect 3227 26822 3273 26881
rect 3410 27353 3538 27392
rect 3410 27301 3448 27353
rect 3500 27301 3538 27353
rect 3410 27242 3538 27301
rect 3410 27196 3451 27242
rect 3497 27196 3538 27242
rect 3410 27137 3538 27196
rect 3410 27135 3451 27137
rect 3497 27135 3538 27137
rect 3410 27083 3448 27135
rect 3500 27083 3538 27135
rect 3410 27032 3538 27083
rect 3410 26986 3451 27032
rect 3497 26986 3538 27032
rect 3410 26927 3538 26986
rect 3410 26917 3451 26927
rect 3497 26917 3538 26927
rect 3410 26865 3448 26917
rect 3500 26865 3538 26917
rect 3410 26825 3538 26865
rect 3675 27347 3721 27396
rect 3899 27392 3945 27406
rect 4088 27452 4204 27546
rect 4536 27665 4652 27754
rect 4795 27745 4841 27754
rect 4984 27665 5100 27758
rect 5202 27794 5240 27846
rect 5292 27794 5330 27846
rect 5897 27834 5933 27873
rect 5979 27834 6013 28082
rect 5897 27821 6013 27834
rect 6121 28082 6237 28135
rect 6121 27834 6157 28082
rect 6203 27834 6237 28082
rect 6324 28131 6362 28183
rect 6414 28131 6461 28183
rect 6324 28082 6461 28131
rect 6324 27965 6381 28082
rect 6324 27913 6362 27965
rect 6324 27873 6381 27913
rect 5202 27758 5243 27794
rect 5289 27758 5330 27794
rect 5202 27754 5330 27758
rect 5243 27745 5289 27754
rect 6121 27733 6237 27834
rect 6345 27834 6381 27873
rect 6427 27834 6461 28082
rect 6546 28185 6670 28225
rect 6546 28133 6582 28185
rect 6634 28133 6670 28185
rect 6546 28026 6670 28133
rect 6546 27967 6587 28026
rect 6633 27967 6670 28026
rect 7708 28126 7836 28292
rect 7708 28074 7746 28126
rect 7798 28074 7836 28126
rect 6546 27915 6582 27967
rect 6634 27915 6670 27967
rect 6546 27886 6587 27915
rect 6633 27886 6670 27915
rect 6546 27875 6670 27886
rect 7527 27996 7573 28009
rect 7527 27876 7573 27950
rect 6345 27821 6461 27834
rect 4536 27546 5100 27665
rect 5825 27683 6005 27695
rect 5825 27631 5837 27683
rect 5994 27637 6005 27683
rect 5993 27631 6005 27637
rect 5825 27619 6005 27631
rect 6121 27614 6461 27733
rect 7527 27702 7573 27830
rect 7708 27996 7836 28074
rect 7708 27950 7751 27996
rect 7797 27950 7836 27996
rect 7708 27908 7836 27950
rect 7708 27856 7746 27908
rect 7798 27856 7836 27908
rect 7708 27830 7751 27856
rect 7797 27830 7836 27856
rect 7708 27816 7836 27830
rect 8997 28325 9125 28384
rect 8997 28282 9038 28325
rect 9084 28282 9125 28325
rect 8997 28230 9035 28282
rect 9087 28230 9125 28282
rect 8997 28220 9125 28230
rect 8997 28174 9038 28220
rect 9084 28174 9125 28220
rect 8997 28116 9125 28174
rect 8997 28070 9038 28116
rect 9084 28070 9125 28116
rect 8997 28064 9125 28070
rect 8997 28012 9035 28064
rect 9087 28012 9125 28064
rect 8997 27966 9038 28012
rect 9084 27966 9125 28012
rect 8997 27908 9125 27966
rect 8997 27862 9038 27908
rect 9084 27862 9125 27908
rect 8997 27846 9125 27862
rect 8997 27794 9035 27846
rect 9087 27794 9125 27846
rect 9262 28535 9308 28594
rect 9451 28640 9567 28939
rect 9451 28594 9486 28640
rect 9532 28594 9567 28640
rect 9451 28540 9567 28594
rect 9710 28640 9756 28653
rect 9710 28540 9756 28594
rect 9899 28640 10015 28939
rect 9899 28594 9934 28640
rect 9980 28594 10015 28640
rect 9262 28430 9308 28489
rect 9262 28325 9308 28384
rect 9262 28220 9308 28279
rect 9262 28116 9308 28174
rect 9262 28012 9308 28070
rect 9262 27908 9308 27966
rect 9262 27804 9308 27862
rect 8997 27758 9038 27794
rect 9084 27758 9125 27794
rect 8997 27754 9125 27758
rect 9227 27758 9262 27795
rect 9437 28539 9567 28540
rect 9437 28535 9565 28539
rect 9437 28500 9486 28535
rect 9437 28448 9475 28500
rect 9532 28489 9565 28535
rect 9527 28448 9565 28489
rect 9437 28430 9565 28448
rect 9437 28384 9486 28430
rect 9532 28384 9565 28430
rect 9437 28325 9565 28384
rect 9437 28282 9486 28325
rect 9437 28230 9475 28282
rect 9532 28279 9565 28325
rect 9527 28230 9565 28279
rect 9437 28220 9565 28230
rect 9437 28174 9486 28220
rect 9532 28174 9565 28220
rect 9437 28116 9565 28174
rect 9437 28070 9486 28116
rect 9532 28070 9565 28116
rect 9437 28064 9565 28070
rect 9437 28012 9475 28064
rect 9527 28012 9565 28064
rect 9437 27966 9486 28012
rect 9532 27966 9565 28012
rect 9437 27908 9565 27966
rect 9437 27862 9486 27908
rect 9532 27862 9565 27908
rect 9437 27846 9565 27862
rect 9308 27758 9343 27795
rect 9038 27745 9084 27754
rect 8742 27702 8866 27735
rect 7527 27695 8868 27702
rect 6753 27683 6933 27695
rect 6753 27631 6765 27683
rect 6921 27631 6933 27683
rect 6753 27619 6933 27631
rect 4088 27406 4123 27452
rect 4169 27406 4204 27452
rect 4088 27396 4204 27406
rect 4347 27452 4393 27465
rect 3675 27242 3721 27301
rect 3675 27137 3721 27196
rect 3675 27032 3721 27091
rect 3675 26927 3721 26986
rect 3227 26717 3273 26776
rect 3227 26612 3273 26671
rect 3227 26507 3273 26566
rect 3227 26402 3273 26461
rect 3227 26297 3273 26356
rect 3227 26192 3273 26251
rect 3227 26088 3273 26146
rect 3227 25984 3273 26042
rect 3227 25880 3273 25938
rect 3227 25776 3273 25834
rect 3227 25672 3273 25730
rect 3227 25568 3273 25626
rect 3227 25464 3273 25522
rect 3227 25360 3273 25418
rect 3227 25256 3273 25314
rect 3227 25197 3273 25210
rect 3451 26822 3497 26825
rect 3451 26717 3497 26776
rect 3451 26612 3497 26671
rect 3451 26507 3497 26566
rect 3451 26402 3497 26461
rect 3451 26297 3497 26356
rect 3451 26192 3497 26251
rect 3451 26088 3497 26146
rect 3451 25984 3497 26042
rect 3451 25880 3497 25938
rect 3451 25776 3497 25834
rect 3451 25672 3497 25730
rect 3451 25568 3497 25626
rect 3451 25464 3497 25522
rect 3451 25360 3497 25418
rect 3451 25256 3497 25314
rect 3451 25197 3497 25210
rect 3675 26822 3721 26881
rect 3858 27353 3986 27392
rect 3858 27301 3896 27353
rect 3948 27301 3986 27353
rect 3858 27242 3986 27301
rect 3858 27196 3899 27242
rect 3945 27196 3986 27242
rect 3858 27137 3986 27196
rect 3858 27135 3899 27137
rect 3945 27135 3986 27137
rect 3858 27083 3896 27135
rect 3948 27083 3986 27135
rect 3858 27032 3986 27083
rect 3858 26986 3899 27032
rect 3945 26986 3986 27032
rect 3858 26927 3986 26986
rect 3858 26917 3899 26927
rect 3945 26917 3986 26927
rect 3858 26865 3896 26917
rect 3948 26865 3986 26917
rect 3858 26825 3986 26865
rect 4123 27347 4169 27396
rect 4347 27392 4393 27406
rect 4536 27452 4652 27546
rect 4536 27406 4571 27452
rect 4617 27406 4652 27452
rect 4536 27396 4652 27406
rect 4795 27452 4841 27465
rect 4123 27242 4169 27301
rect 4123 27137 4169 27196
rect 4123 27032 4169 27091
rect 4123 26927 4169 26986
rect 3675 26717 3721 26776
rect 3675 26612 3721 26671
rect 3675 26507 3721 26566
rect 3675 26402 3721 26461
rect 3675 26297 3721 26356
rect 3675 26192 3721 26251
rect 3675 26088 3721 26146
rect 3675 25984 3721 26042
rect 3675 25880 3721 25938
rect 3675 25776 3721 25834
rect 3675 25672 3721 25730
rect 3675 25568 3721 25626
rect 3675 25464 3721 25522
rect 3675 25360 3721 25418
rect 3675 25256 3721 25314
rect 3675 25197 3721 25210
rect 3899 26822 3945 26825
rect 3899 26717 3945 26776
rect 3899 26612 3945 26671
rect 3899 26507 3945 26566
rect 3899 26402 3945 26461
rect 3899 26297 3945 26356
rect 3899 26192 3945 26251
rect 3899 26088 3945 26146
rect 3899 25984 3945 26042
rect 3899 25880 3945 25938
rect 3899 25776 3945 25834
rect 3899 25672 3945 25730
rect 3899 25568 3945 25626
rect 3899 25464 3945 25522
rect 3899 25360 3945 25418
rect 3899 25256 3945 25314
rect 3899 25197 3945 25210
rect 4123 26822 4169 26881
rect 4306 27353 4434 27392
rect 4306 27301 4344 27353
rect 4396 27301 4434 27353
rect 4306 27242 4434 27301
rect 4306 27196 4347 27242
rect 4393 27196 4434 27242
rect 4306 27137 4434 27196
rect 4306 27135 4347 27137
rect 4393 27135 4434 27137
rect 4306 27083 4344 27135
rect 4396 27083 4434 27135
rect 4306 27032 4434 27083
rect 4306 26986 4347 27032
rect 4393 26986 4434 27032
rect 4306 26927 4434 26986
rect 4306 26917 4347 26927
rect 4393 26917 4434 26927
rect 4306 26865 4344 26917
rect 4396 26865 4434 26917
rect 4306 26825 4434 26865
rect 4571 27347 4617 27396
rect 4795 27392 4841 27406
rect 4984 27452 5100 27546
rect 4984 27406 5019 27452
rect 5065 27406 5100 27452
rect 4984 27396 5100 27406
rect 5243 27452 5289 27465
rect 5897 27418 6013 27432
rect 4571 27242 4617 27301
rect 4571 27137 4617 27196
rect 4571 27032 4617 27091
rect 4571 26927 4617 26986
rect 4123 26717 4169 26776
rect 4123 26612 4169 26671
rect 4123 26507 4169 26566
rect 4123 26402 4169 26461
rect 4123 26297 4169 26356
rect 4123 26192 4169 26251
rect 4123 26088 4169 26146
rect 4123 25984 4169 26042
rect 4123 25880 4169 25938
rect 4123 25776 4169 25834
rect 4123 25672 4169 25730
rect 4123 25568 4169 25626
rect 4123 25464 4169 25522
rect 4123 25360 4169 25418
rect 4123 25256 4169 25314
rect 4123 25197 4169 25210
rect 4347 26822 4393 26825
rect 4347 26717 4393 26776
rect 4347 26612 4393 26671
rect 4347 26507 4393 26566
rect 4347 26402 4393 26461
rect 4347 26297 4393 26356
rect 4347 26192 4393 26251
rect 4347 26088 4393 26146
rect 4347 25984 4393 26042
rect 4347 25880 4393 25938
rect 4347 25776 4393 25834
rect 4347 25672 4393 25730
rect 4347 25568 4393 25626
rect 4347 25464 4393 25522
rect 4347 25360 4393 25418
rect 4347 25256 4393 25314
rect 4347 25197 4393 25210
rect 4571 26822 4617 26881
rect 4754 27353 4882 27392
rect 4754 27301 4792 27353
rect 4844 27301 4882 27353
rect 4754 27242 4882 27301
rect 4754 27196 4795 27242
rect 4841 27196 4882 27242
rect 4754 27137 4882 27196
rect 4754 27135 4795 27137
rect 4841 27135 4882 27137
rect 4754 27083 4792 27135
rect 4844 27083 4882 27135
rect 4754 27032 4882 27083
rect 4754 26986 4795 27032
rect 4841 26986 4882 27032
rect 4754 26927 4882 26986
rect 4754 26917 4795 26927
rect 4841 26917 4882 26927
rect 4754 26865 4792 26917
rect 4844 26865 4882 26917
rect 4754 26825 4882 26865
rect 5019 27347 5065 27396
rect 5243 27392 5289 27406
rect 5019 27242 5065 27301
rect 5019 27137 5065 27196
rect 5019 27032 5065 27091
rect 5019 26927 5065 26986
rect 4571 26717 4617 26776
rect 4571 26612 4617 26671
rect 4571 26507 4617 26566
rect 4571 26402 4617 26461
rect 4571 26297 4617 26356
rect 4571 26192 4617 26251
rect 4571 26088 4617 26146
rect 4571 25984 4617 26042
rect 4571 25880 4617 25938
rect 4571 25776 4617 25834
rect 4571 25672 4617 25730
rect 4571 25568 4617 25626
rect 4571 25464 4617 25522
rect 4571 25360 4617 25418
rect 4571 25256 4617 25314
rect 4571 25197 4617 25210
rect 4795 26822 4841 26825
rect 4795 26717 4841 26776
rect 4795 26612 4841 26671
rect 4795 26507 4841 26566
rect 4795 26402 4841 26461
rect 4795 26297 4841 26356
rect 4795 26192 4841 26251
rect 4795 26088 4841 26146
rect 4795 25984 4841 26042
rect 4795 25880 4841 25938
rect 4795 25776 4841 25834
rect 4795 25672 4841 25730
rect 4795 25568 4841 25626
rect 4795 25464 4841 25522
rect 4795 25360 4841 25418
rect 4795 25256 4841 25314
rect 4795 25197 4841 25210
rect 5019 26822 5065 26881
rect 5202 27353 5330 27392
rect 5202 27301 5240 27353
rect 5292 27301 5330 27353
rect 5202 27242 5330 27301
rect 5202 27196 5243 27242
rect 5289 27196 5330 27242
rect 5202 27137 5330 27196
rect 5202 27135 5243 27137
rect 5289 27135 5330 27137
rect 5202 27083 5240 27135
rect 5292 27083 5330 27135
rect 5202 27032 5330 27083
rect 5611 27378 5735 27418
rect 5611 27326 5647 27378
rect 5699 27326 5735 27378
rect 5611 27160 5649 27326
rect 5695 27160 5735 27326
rect 5611 27108 5647 27160
rect 5699 27108 5735 27160
rect 5611 27068 5735 27108
rect 5887 27382 6013 27418
rect 5887 27378 5933 27382
rect 5887 27326 5923 27378
rect 5979 27336 6013 27382
rect 5975 27326 6013 27336
rect 5887 27178 6013 27326
rect 5887 27160 5933 27178
rect 5887 27108 5923 27160
rect 5979 27132 6013 27178
rect 5975 27108 6013 27132
rect 5887 27095 6013 27108
rect 6345 27382 6461 27614
rect 6771 27574 6933 27619
rect 6771 27528 6782 27574
rect 6922 27528 6933 27574
rect 7527 27643 8778 27695
rect 8830 27643 8868 27695
rect 7527 27568 8868 27643
rect 9227 27665 9343 27758
rect 9437 27794 9475 27846
rect 9527 27804 9565 27846
rect 9437 27758 9486 27794
rect 9532 27758 9565 27804
rect 9437 27754 9565 27758
rect 9669 28535 9797 28540
rect 9899 28539 10015 28594
rect 10158 28640 10204 28653
rect 10158 28540 10204 28594
rect 10347 28640 10463 28939
rect 10347 28594 10382 28640
rect 10428 28594 10463 28640
rect 10347 28540 10463 28594
rect 10606 28640 10652 28653
rect 9669 28500 9710 28535
rect 9756 28500 9797 28535
rect 9669 28448 9707 28500
rect 9759 28448 9797 28500
rect 9669 28430 9797 28448
rect 9669 28384 9710 28430
rect 9756 28384 9797 28430
rect 9669 28325 9797 28384
rect 9669 28282 9710 28325
rect 9756 28282 9797 28325
rect 9669 28230 9707 28282
rect 9759 28230 9797 28282
rect 9669 28220 9797 28230
rect 9669 28174 9710 28220
rect 9756 28174 9797 28220
rect 9669 28116 9797 28174
rect 9669 28070 9710 28116
rect 9756 28070 9797 28116
rect 9669 28064 9797 28070
rect 9669 28012 9707 28064
rect 9759 28012 9797 28064
rect 9669 27966 9710 28012
rect 9756 27966 9797 28012
rect 9669 27908 9797 27966
rect 9669 27862 9710 27908
rect 9756 27862 9797 27908
rect 9669 27846 9797 27862
rect 9669 27794 9707 27846
rect 9759 27794 9797 27846
rect 9669 27758 9710 27794
rect 9756 27758 9797 27794
rect 9669 27754 9797 27758
rect 9934 28535 9980 28539
rect 9934 28430 9980 28489
rect 9934 28325 9980 28384
rect 9934 28220 9980 28279
rect 9934 28116 9980 28174
rect 9934 28012 9980 28070
rect 9934 27908 9980 27966
rect 9934 27804 9980 27862
rect 9486 27745 9532 27754
rect 9675 27665 9791 27754
rect 9934 27745 9980 27758
rect 10117 28535 10245 28540
rect 10347 28539 10477 28540
rect 10117 28500 10158 28535
rect 10204 28500 10245 28535
rect 10117 28448 10155 28500
rect 10207 28448 10245 28500
rect 10117 28430 10245 28448
rect 10117 28384 10158 28430
rect 10204 28384 10245 28430
rect 10117 28325 10245 28384
rect 10117 28282 10158 28325
rect 10204 28282 10245 28325
rect 10117 28230 10155 28282
rect 10207 28230 10245 28282
rect 10117 28220 10245 28230
rect 10117 28174 10158 28220
rect 10204 28174 10245 28220
rect 10117 28116 10245 28174
rect 10117 28070 10158 28116
rect 10204 28070 10245 28116
rect 10117 28064 10245 28070
rect 10117 28012 10155 28064
rect 10207 28012 10245 28064
rect 10117 27966 10158 28012
rect 10204 27966 10245 28012
rect 10117 27908 10245 27966
rect 10117 27862 10158 27908
rect 10204 27862 10245 27908
rect 10117 27846 10245 27862
rect 10117 27794 10155 27846
rect 10207 27794 10245 27846
rect 10117 27758 10158 27794
rect 10204 27758 10245 27794
rect 10117 27754 10245 27758
rect 10349 28535 10477 28539
rect 10349 28489 10382 28535
rect 10428 28500 10477 28535
rect 10349 28448 10387 28489
rect 10439 28448 10477 28500
rect 10349 28430 10477 28448
rect 10349 28384 10382 28430
rect 10428 28384 10477 28430
rect 10349 28325 10477 28384
rect 10349 28279 10382 28325
rect 10428 28282 10477 28325
rect 10349 28230 10387 28279
rect 10439 28230 10477 28282
rect 10349 28220 10477 28230
rect 10349 28174 10382 28220
rect 10428 28174 10477 28220
rect 10349 28116 10477 28174
rect 10349 28070 10382 28116
rect 10428 28070 10477 28116
rect 10349 28064 10477 28070
rect 10349 28012 10387 28064
rect 10439 28012 10477 28064
rect 10349 27966 10382 28012
rect 10428 27966 10477 28012
rect 10349 27908 10477 27966
rect 10349 27862 10382 27908
rect 10428 27862 10477 27908
rect 10349 27846 10477 27862
rect 10349 27804 10387 27846
rect 10349 27758 10382 27804
rect 10439 27794 10477 27846
rect 10606 28535 10652 28594
rect 10795 28640 10911 28939
rect 10795 28594 10830 28640
rect 10876 28594 10911 28640
rect 10795 28540 10911 28594
rect 11054 28640 11100 28653
rect 10606 28430 10652 28489
rect 10606 28325 10652 28384
rect 10606 28220 10652 28279
rect 10606 28116 10652 28174
rect 10606 28012 10652 28070
rect 10606 27908 10652 27966
rect 10606 27804 10652 27862
rect 10428 27758 10477 27794
rect 10349 27754 10477 27758
rect 10571 27758 10606 27795
rect 10789 28535 10917 28540
rect 10789 28500 10830 28535
rect 10876 28500 10917 28535
rect 10789 28448 10827 28500
rect 10879 28448 10917 28500
rect 10789 28430 10917 28448
rect 10789 28384 10830 28430
rect 10876 28384 10917 28430
rect 10789 28325 10917 28384
rect 10789 28282 10830 28325
rect 10876 28282 10917 28325
rect 10789 28230 10827 28282
rect 10879 28230 10917 28282
rect 10789 28220 10917 28230
rect 10789 28174 10830 28220
rect 10876 28174 10917 28220
rect 10789 28116 10917 28174
rect 10789 28070 10830 28116
rect 10876 28070 10917 28116
rect 10789 28064 10917 28070
rect 10789 28012 10827 28064
rect 10879 28012 10917 28064
rect 10789 27966 10830 28012
rect 10876 27966 10917 28012
rect 10789 27908 10917 27966
rect 10789 27862 10830 27908
rect 10876 27862 10917 27908
rect 10789 27846 10917 27862
rect 10652 27758 10687 27795
rect 6771 27517 6933 27528
rect 6345 27336 6381 27382
rect 6427 27336 6461 27382
rect 6345 27178 6461 27336
rect 6345 27132 6381 27178
rect 6427 27132 6461 27178
rect 5887 27068 6011 27095
rect 5202 26986 5243 27032
rect 5289 26986 5330 27032
rect 5202 26927 5330 26986
rect 5202 26917 5243 26927
rect 5289 26917 5330 26927
rect 5202 26865 5240 26917
rect 5292 26865 5330 26917
rect 6345 27015 6461 27132
rect 6793 27382 7455 27432
rect 6793 27336 6829 27382
rect 6875 27336 7455 27382
rect 6793 27315 7455 27336
rect 6793 27269 7409 27315
rect 6793 27210 7455 27269
rect 6793 27178 7007 27210
rect 6793 27132 6829 27178
rect 6875 27158 7007 27178
rect 7059 27158 7219 27210
rect 7271 27159 7455 27210
rect 7271 27158 7409 27159
rect 6875 27132 7409 27158
rect 6793 27113 7409 27132
rect 6793 27100 7455 27113
rect 7633 27315 7679 27568
rect 8742 27477 8866 27568
rect 7633 27159 7679 27269
rect 7633 27100 7679 27113
rect 7857 27392 8227 27432
rect 7857 27340 8136 27392
rect 8188 27340 8227 27392
rect 8742 27425 8778 27477
rect 8830 27425 8866 27477
rect 9227 27546 9791 27665
rect 8742 27385 8866 27425
rect 9038 27452 9084 27465
rect 9038 27392 9084 27406
rect 9227 27452 9343 27546
rect 9227 27406 9262 27452
rect 9308 27406 9343 27452
rect 9227 27396 9343 27406
rect 9486 27452 9532 27465
rect 7857 27315 8141 27340
rect 7903 27269 8141 27315
rect 7857 27174 8141 27269
rect 8187 27174 8227 27340
rect 7857 27159 8136 27174
rect 7903 27122 8136 27159
rect 8188 27122 8227 27174
rect 7903 27113 8227 27122
rect 7857 27108 8227 27113
rect 8997 27353 9125 27392
rect 8997 27301 9035 27353
rect 9087 27301 9125 27353
rect 8997 27242 9125 27301
rect 8997 27196 9038 27242
rect 9084 27196 9125 27242
rect 8997 27137 9125 27196
rect 8997 27135 9038 27137
rect 9084 27135 9125 27137
rect 7857 27100 7903 27108
rect 6793 27095 6909 27100
rect 8100 27082 8224 27108
rect 8997 27083 9035 27135
rect 9087 27083 9125 27135
rect 8997 27032 9125 27083
rect 7539 27021 7795 27032
rect 7539 27015 7550 27021
rect 6345 26975 7550 27015
rect 7784 26975 7795 27021
rect 6345 26974 7795 26975
rect 6345 26922 7005 26974
rect 7057 26922 7217 26974
rect 7269 26922 7795 26974
rect 6345 26895 7795 26922
rect 8997 26986 9038 27032
rect 9084 26986 9125 27032
rect 8997 26927 9125 26986
rect 8997 26917 9038 26927
rect 9084 26917 9125 26927
rect 6967 26882 7307 26895
rect 5202 26825 5330 26865
rect 8997 26865 9035 26917
rect 9087 26865 9125 26917
rect 8997 26825 9125 26865
rect 9262 27347 9308 27396
rect 9486 27392 9532 27406
rect 9675 27452 9791 27546
rect 10123 27665 10239 27754
rect 10382 27745 10428 27754
rect 10571 27665 10687 27758
rect 10789 27794 10827 27846
rect 10879 27794 10917 27846
rect 11054 28535 11100 28594
rect 11243 28640 11359 28939
rect 11243 28594 11278 28640
rect 11324 28594 11359 28640
rect 11243 28540 11359 28594
rect 11502 28640 11548 28653
rect 11502 28540 11548 28594
rect 11691 28640 11807 28939
rect 11691 28594 11726 28640
rect 11772 28594 11807 28640
rect 11054 28430 11100 28489
rect 11054 28325 11100 28384
rect 11054 28220 11100 28279
rect 11054 28116 11100 28174
rect 11054 28012 11100 28070
rect 11054 27908 11100 27966
rect 11054 27804 11100 27862
rect 10789 27758 10830 27794
rect 10876 27758 10917 27794
rect 10789 27754 10917 27758
rect 11019 27758 11054 27795
rect 11229 28539 11359 28540
rect 11229 28535 11357 28539
rect 11229 28500 11278 28535
rect 11229 28448 11267 28500
rect 11324 28489 11357 28535
rect 11319 28448 11357 28489
rect 11229 28430 11357 28448
rect 11229 28384 11278 28430
rect 11324 28384 11357 28430
rect 11229 28325 11357 28384
rect 11229 28282 11278 28325
rect 11229 28230 11267 28282
rect 11324 28279 11357 28325
rect 11319 28230 11357 28279
rect 11229 28220 11357 28230
rect 11229 28174 11278 28220
rect 11324 28174 11357 28220
rect 11229 28116 11357 28174
rect 11229 28070 11278 28116
rect 11324 28070 11357 28116
rect 11229 28064 11357 28070
rect 11229 28012 11267 28064
rect 11319 28012 11357 28064
rect 11229 27966 11278 28012
rect 11324 27966 11357 28012
rect 11229 27908 11357 27966
rect 11229 27862 11278 27908
rect 11324 27862 11357 27908
rect 11229 27846 11357 27862
rect 11100 27758 11135 27795
rect 10830 27745 10876 27754
rect 10123 27546 10687 27665
rect 9675 27406 9710 27452
rect 9756 27406 9791 27452
rect 9675 27396 9791 27406
rect 9934 27452 9980 27465
rect 9262 27242 9308 27301
rect 9262 27137 9308 27196
rect 9262 27032 9308 27091
rect 9262 26927 9308 26986
rect 5019 26717 5065 26776
rect 5019 26612 5065 26671
rect 5019 26507 5065 26566
rect 5019 26402 5065 26461
rect 5019 26297 5065 26356
rect 5019 26192 5065 26251
rect 5019 26088 5065 26146
rect 5019 25984 5065 26042
rect 5019 25880 5065 25938
rect 5019 25776 5065 25834
rect 5019 25672 5065 25730
rect 5019 25568 5065 25626
rect 5019 25464 5065 25522
rect 5019 25360 5065 25418
rect 5019 25256 5065 25314
rect 5019 25197 5065 25210
rect 5243 26822 5289 26825
rect 5243 26717 5289 26776
rect 9038 26822 9084 26825
rect 5243 26612 5289 26671
rect 6091 26731 6137 26744
rect 5243 26507 5289 26566
rect 5243 26402 5289 26461
rect 5243 26297 5289 26356
rect 5243 26192 5289 26251
rect 5243 26088 5289 26146
rect 5243 25984 5289 26042
rect 5243 25880 5289 25938
rect 5243 25776 5289 25834
rect 5243 25672 5289 25730
rect 5243 25568 5289 25626
rect 5243 25464 5289 25522
rect 5243 25360 5289 25418
rect 5739 26545 6091 26643
rect 5739 26499 5787 26545
rect 5833 26514 6091 26545
rect 6315 26731 6361 26744
rect 5833 26499 5874 26514
rect 5739 26462 5874 26499
rect 5926 26462 6081 26514
rect 5739 26382 6091 26462
rect 5739 26336 5787 26382
rect 5833 26379 6091 26382
rect 6137 26379 6171 26643
rect 5833 26336 6171 26379
rect 5739 26322 6171 26336
rect 5739 26296 6091 26322
rect 5739 26244 5874 26296
rect 5926 26244 6081 26296
rect 6137 26276 6171 26322
rect 6133 26244 6171 26276
rect 5739 26219 6171 26244
rect 5739 26218 6091 26219
rect 5739 26172 5787 26218
rect 5833 26173 6091 26218
rect 6137 26173 6171 26219
rect 5833 26172 6171 26173
rect 5739 26116 6171 26172
rect 5739 26078 6091 26116
rect 5739 26055 5874 26078
rect 5739 26009 5787 26055
rect 5833 26026 5874 26055
rect 5926 26026 6081 26078
rect 6137 26070 6171 26116
rect 6133 26026 6171 26070
rect 5833 26013 6171 26026
rect 5833 26009 6091 26013
rect 5739 25967 6091 26009
rect 6137 25967 6171 26013
rect 5739 25910 6171 25967
rect 5739 25892 6091 25910
rect 5739 25846 5787 25892
rect 5833 25864 6091 25892
rect 6137 25864 6171 25910
rect 5833 25860 6171 25864
rect 5833 25846 5874 25860
rect 5739 25808 5874 25846
rect 5926 25808 6081 25860
rect 6133 25808 6171 25860
rect 5739 25807 6171 25808
rect 5739 25761 6091 25807
rect 6137 25761 6171 25807
rect 5739 25728 6171 25761
rect 5739 25682 5787 25728
rect 5833 25704 6171 25728
rect 5833 25682 6091 25704
rect 5739 25658 6091 25682
rect 6137 25658 6171 25704
rect 5739 25601 6171 25658
rect 5739 25565 6091 25601
rect 5739 25519 5787 25565
rect 5833 25555 6091 25565
rect 6137 25555 6171 25601
rect 5833 25519 6171 25555
rect 5739 25498 6171 25519
rect 5739 25452 6091 25498
rect 6137 25452 6171 25498
rect 5739 25395 6171 25452
rect 7782 26731 7828 26744
rect 7430 26545 7782 26643
rect 6315 26322 6361 26379
rect 6315 26219 6361 26276
rect 6315 26116 6361 26173
rect 6315 26013 6361 26070
rect 6315 25910 6361 25967
rect 6315 25807 6361 25864
rect 6315 25704 6361 25761
rect 6563 26491 6691 26531
rect 6563 26439 6601 26491
rect 6653 26439 6691 26491
rect 7430 26499 7478 26545
rect 7524 26514 7782 26545
rect 8006 26731 8052 26744
rect 7524 26499 7565 26514
rect 7430 26462 7565 26499
rect 7617 26462 7772 26514
rect 6563 26400 6605 26439
rect 6651 26400 6691 26439
rect 6563 26338 6691 26400
rect 6563 26292 6605 26338
rect 6651 26292 6691 26338
rect 6563 26273 6691 26292
rect 6563 26221 6601 26273
rect 6653 26221 6691 26273
rect 6563 26184 6605 26221
rect 6651 26184 6691 26221
rect 6563 26122 6691 26184
rect 6563 26076 6605 26122
rect 6651 26076 6691 26122
rect 6563 26055 6691 26076
rect 6563 26003 6601 26055
rect 6653 26003 6691 26055
rect 6563 25968 6605 26003
rect 6651 25968 6691 26003
rect 6563 25906 6691 25968
rect 6563 25860 6605 25906
rect 6651 25860 6691 25906
rect 6563 25837 6691 25860
rect 6563 25785 6601 25837
rect 6653 25785 6691 25837
rect 6563 25752 6605 25785
rect 6651 25752 6691 25785
rect 6563 25745 6691 25752
rect 6829 26446 6875 26459
rect 6829 26338 6875 26400
rect 6829 26230 6875 26292
rect 6829 26122 6875 26184
rect 6829 26014 6875 26076
rect 6829 25906 6875 25968
rect 6829 25798 6875 25860
rect 6315 25601 6361 25658
rect 6315 25498 6361 25555
rect 6315 25405 6361 25452
rect 6605 25690 6651 25745
rect 6605 25582 6651 25644
rect 6605 25474 6651 25536
rect 6605 25415 6651 25428
rect 6829 25690 6875 25752
rect 6829 25582 6875 25644
rect 6829 25474 6875 25536
rect 5739 25349 6091 25395
rect 6137 25349 6171 25395
rect 5739 25344 6171 25349
rect 6280 25395 6395 25405
rect 6280 25349 6315 25395
rect 6361 25349 6395 25395
rect 6091 25336 6137 25344
rect 5243 25256 5289 25314
rect 5243 25197 5289 25210
rect 5836 25255 6176 25262
rect 6280 25255 6395 25349
rect 5836 25221 6193 25255
rect 5836 25169 5874 25221
rect 5926 25218 6086 25221
rect 6138 25218 6193 25221
rect 5926 25172 5954 25218
rect 6000 25172 6086 25218
rect 6158 25172 6193 25218
rect 5926 25169 6086 25172
rect 6138 25169 6193 25172
rect 5836 25135 6193 25169
rect 6280 25218 6703 25255
rect 6280 25172 6464 25218
rect 6510 25172 6622 25218
rect 6668 25172 6703 25218
rect 6280 25135 6703 25172
rect 5836 25129 6176 25135
rect 1736 25088 2524 25126
rect 1736 25042 1895 25088
rect 2317 25042 2524 25088
rect 1736 25007 2524 25042
rect 2632 25088 3420 25126
rect 2632 25042 2839 25088
rect 3261 25042 3420 25088
rect 2632 25007 3420 25042
rect 3528 25088 4316 25126
rect 3528 25042 3687 25088
rect 4109 25042 4316 25088
rect 3528 25007 4316 25042
rect 4424 25088 5212 25126
rect 4424 25042 4631 25088
rect 5053 25042 5212 25088
rect 4424 25007 5212 25042
rect 2006 25006 2123 25007
rect 3033 25006 3150 25007
rect 1484 24854 1898 24890
rect 1484 24808 1659 24854
rect 1705 24808 1818 24854
rect 1864 24813 1898 24854
rect 1864 24808 1907 24813
rect 1484 24773 1907 24808
rect 1484 24771 1817 24773
rect 1779 24721 1817 24771
rect 1869 24721 1907 24773
rect 1779 24556 1907 24721
rect 1779 22722 1817 24556
rect 1869 24504 1907 24556
rect 1863 24338 1907 24504
rect 2006 24550 2122 25006
rect 2006 24456 2041 24550
rect 1869 24286 1907 24338
rect 1863 24121 1907 24286
rect 1869 24069 1907 24121
rect 1863 23903 1907 24069
rect 1869 23851 1907 23903
rect 1863 23685 1907 23851
rect 1869 23633 1907 23685
rect 1863 23467 1907 23633
rect 1869 23415 1907 23467
rect 1863 23250 1907 23415
rect 1869 23198 1907 23250
rect 1863 23032 1907 23198
rect 1869 22980 1907 23032
rect 1863 22815 1907 22980
rect 1869 22763 1907 22815
rect 1863 22722 1907 22763
rect 1817 22509 1863 22566
rect 1817 22406 1863 22463
rect 1817 22303 1863 22360
rect 1817 22200 1863 22257
rect 1817 22097 1863 22154
rect 1817 21994 1863 22051
rect 1817 21891 1863 21948
rect 2087 24456 2122 24550
rect 2230 24854 2926 24890
rect 2230 24808 2266 24854
rect 2312 24808 2424 24854
rect 2470 24808 2686 24854
rect 2732 24808 2844 24854
rect 2890 24808 2926 24854
rect 2230 24773 2926 24808
rect 2230 24721 2269 24773
rect 2321 24721 2552 24773
rect 2604 24721 2835 24773
rect 2887 24721 2926 24773
rect 2230 24556 2926 24721
rect 2230 24550 2269 24556
rect 2041 22509 2087 22566
rect 2041 22406 2087 22463
rect 2041 22303 2087 22360
rect 2041 22200 2087 22257
rect 2041 22097 2087 22154
rect 2041 21994 2087 22051
rect 2041 21891 2087 21948
rect 1817 21788 1863 21845
rect 1817 21685 1863 21742
rect 1817 21582 1863 21639
rect 1817 21523 1863 21536
rect 2003 21845 2041 21882
rect 2230 22566 2265 24550
rect 2321 24504 2552 24556
rect 2604 24504 2835 24556
rect 2887 24550 2926 24556
rect 2311 24338 2845 24504
rect 2321 24286 2552 24338
rect 2604 24286 2835 24338
rect 2311 24121 2845 24286
rect 2321 24069 2552 24121
rect 2604 24069 2835 24121
rect 2311 23903 2845 24069
rect 2321 23851 2552 23903
rect 2604 23851 2835 23903
rect 2311 23685 2845 23851
rect 2321 23633 2552 23685
rect 2604 23633 2835 23685
rect 2311 23467 2845 23633
rect 2321 23415 2552 23467
rect 2604 23415 2835 23467
rect 2311 23250 2845 23415
rect 2321 23198 2552 23250
rect 2604 23198 2835 23250
rect 2311 23032 2845 23198
rect 2321 22980 2552 23032
rect 2604 22980 2835 23032
rect 2311 22815 2845 22980
rect 2321 22763 2552 22815
rect 2604 22763 2835 22815
rect 2311 22566 2845 22763
rect 2891 22566 2926 24550
rect 3034 24550 3150 25006
rect 3798 25006 3915 25007
rect 4825 25006 4942 25007
rect 6091 25006 6137 25015
rect 3258 24854 3690 24890
rect 3258 24813 3292 24854
rect 3034 24456 3069 24550
rect 2230 22509 2926 22566
rect 2230 22463 2265 22509
rect 2311 22463 2845 22509
rect 2891 22463 2926 22509
rect 2230 22406 2926 22463
rect 2230 22360 2265 22406
rect 2311 22360 2845 22406
rect 2891 22360 2926 22406
rect 2230 22303 2926 22360
rect 2230 22257 2265 22303
rect 2311 22257 2845 22303
rect 2891 22257 2926 22303
rect 2230 22200 2926 22257
rect 2230 22154 2265 22200
rect 2311 22154 2845 22200
rect 2891 22154 2926 22200
rect 2230 22097 2926 22154
rect 2230 22051 2265 22097
rect 2311 22051 2845 22097
rect 2891 22051 2926 22097
rect 2230 21994 2926 22051
rect 2230 21948 2265 21994
rect 2311 21989 2845 21994
rect 2311 21948 2555 21989
rect 2230 21891 2555 21948
rect 2087 21845 2127 21882
rect 2003 21842 2127 21845
rect 2003 21790 2039 21842
rect 2091 21790 2127 21842
rect 2003 21788 2127 21790
rect 2003 21742 2041 21788
rect 2087 21742 2127 21788
rect 2003 21685 2127 21742
rect 2003 21639 2041 21685
rect 2087 21639 2127 21685
rect 2003 21624 2127 21639
rect 2003 21572 2039 21624
rect 2091 21572 2127 21624
rect 2003 21536 2041 21572
rect 2087 21536 2127 21572
rect 2003 21532 2127 21536
rect 2230 21845 2265 21891
rect 2311 21845 2555 21891
rect 2230 21788 2555 21845
rect 2230 21742 2265 21788
rect 2311 21742 2555 21788
rect 2230 21685 2555 21742
rect 2230 21639 2265 21685
rect 2311 21661 2555 21685
rect 2601 21948 2845 21989
rect 2891 21948 2926 21994
rect 2601 21891 2926 21948
rect 2601 21845 2845 21891
rect 2891 21845 2926 21891
rect 3115 24456 3150 24550
rect 3249 24808 3292 24813
rect 3338 24808 3451 24854
rect 3497 24808 3610 24854
rect 3656 24813 3690 24854
rect 3656 24808 3699 24813
rect 3249 24773 3699 24808
rect 3249 24721 3287 24773
rect 3339 24771 3609 24773
rect 3339 24721 3377 24771
rect 3249 24556 3377 24721
rect 3249 24504 3287 24556
rect 3249 24338 3293 24504
rect 3249 24286 3287 24338
rect 3249 24121 3293 24286
rect 3249 24069 3287 24121
rect 3249 23903 3293 24069
rect 3249 23851 3287 23903
rect 3249 23685 3293 23851
rect 3249 23633 3287 23685
rect 3249 23467 3293 23633
rect 3249 23415 3287 23467
rect 3249 23250 3293 23415
rect 3249 23198 3287 23250
rect 3249 23032 3293 23198
rect 3249 22980 3287 23032
rect 3249 22815 3293 22980
rect 3249 22763 3287 22815
rect 3249 22722 3293 22763
rect 3069 22509 3115 22566
rect 3069 22406 3115 22463
rect 3069 22303 3115 22360
rect 3069 22200 3115 22257
rect 3069 22097 3115 22154
rect 3069 21994 3115 22051
rect 3069 21891 3115 21948
rect 2601 21788 2926 21845
rect 2601 21742 2845 21788
rect 2891 21742 2926 21788
rect 2601 21685 2926 21742
rect 2601 21661 2845 21685
rect 2311 21639 2845 21661
rect 2891 21639 2926 21685
rect 2230 21582 2926 21639
rect 2230 21536 2265 21582
rect 2311 21536 2845 21582
rect 2891 21536 2926 21582
rect 2041 21523 2087 21532
rect 2230 21531 2926 21536
rect 3029 21845 3069 21882
rect 3339 22722 3377 24556
rect 3571 24721 3609 24771
rect 3661 24721 3699 24773
rect 3571 24556 3699 24721
rect 3571 22722 3609 24556
rect 3661 24504 3699 24556
rect 3655 24338 3699 24504
rect 3798 24550 3914 25006
rect 3798 24456 3833 24550
rect 3661 24286 3699 24338
rect 3655 24121 3699 24286
rect 3661 24069 3699 24121
rect 3655 23903 3699 24069
rect 3661 23851 3699 23903
rect 3655 23685 3699 23851
rect 3661 23633 3699 23685
rect 3655 23467 3699 23633
rect 3661 23415 3699 23467
rect 3655 23250 3699 23415
rect 3661 23198 3699 23250
rect 3655 23032 3699 23198
rect 3661 22980 3699 23032
rect 3655 22815 3699 22980
rect 3661 22763 3699 22815
rect 3293 22509 3339 22566
rect 3293 22406 3339 22463
rect 3293 22303 3339 22360
rect 3293 22200 3339 22257
rect 3293 22097 3339 22154
rect 3293 21994 3339 22051
rect 3293 21891 3339 21948
rect 3115 21845 3153 21882
rect 3029 21842 3153 21845
rect 3029 21790 3065 21842
rect 3117 21790 3153 21842
rect 3029 21788 3153 21790
rect 3029 21742 3069 21788
rect 3115 21742 3153 21788
rect 3029 21685 3153 21742
rect 3029 21639 3069 21685
rect 3115 21639 3153 21685
rect 3029 21624 3153 21639
rect 3029 21572 3065 21624
rect 3117 21572 3153 21624
rect 3029 21536 3069 21572
rect 3115 21536 3153 21572
rect 3029 21532 3153 21536
rect 3293 21788 3339 21845
rect 3293 21685 3339 21742
rect 3293 21582 3339 21639
rect 2265 21523 2311 21531
rect 2845 21523 2891 21531
rect 3069 21523 3115 21532
rect 3293 21523 3339 21536
rect 3655 22722 3699 22763
rect 3609 22509 3655 22566
rect 3609 22406 3655 22463
rect 3609 22303 3655 22360
rect 3609 22200 3655 22257
rect 3609 22097 3655 22154
rect 3609 21994 3655 22051
rect 3609 21891 3655 21948
rect 3879 24456 3914 24550
rect 4022 24854 4718 24890
rect 4022 24808 4058 24854
rect 4104 24808 4216 24854
rect 4262 24808 4478 24854
rect 4524 24808 4636 24854
rect 4682 24808 4718 24854
rect 4022 24773 4718 24808
rect 4022 24721 4061 24773
rect 4113 24721 4344 24773
rect 4396 24721 4627 24773
rect 4679 24721 4718 24773
rect 4022 24556 4718 24721
rect 4022 24550 4061 24556
rect 3833 22509 3879 22566
rect 3833 22406 3879 22463
rect 3833 22303 3879 22360
rect 3833 22200 3879 22257
rect 3833 22097 3879 22154
rect 3833 21994 3879 22051
rect 3833 21891 3879 21948
rect 3609 21788 3655 21845
rect 3609 21685 3655 21742
rect 3609 21582 3655 21639
rect 3609 21523 3655 21536
rect 3795 21845 3833 21882
rect 4022 22566 4057 24550
rect 4113 24504 4344 24556
rect 4396 24504 4627 24556
rect 4679 24550 4718 24556
rect 4103 24338 4637 24504
rect 4113 24286 4344 24338
rect 4396 24286 4627 24338
rect 4103 24121 4637 24286
rect 4113 24069 4344 24121
rect 4396 24069 4627 24121
rect 4103 23903 4637 24069
rect 4113 23851 4344 23903
rect 4396 23851 4627 23903
rect 4103 23685 4637 23851
rect 4113 23633 4344 23685
rect 4396 23633 4627 23685
rect 4103 23467 4637 23633
rect 4113 23415 4344 23467
rect 4396 23415 4627 23467
rect 4103 23250 4637 23415
rect 4113 23198 4344 23250
rect 4396 23198 4627 23250
rect 4103 23032 4637 23198
rect 4113 22980 4344 23032
rect 4396 22980 4627 23032
rect 4103 22815 4637 22980
rect 4113 22763 4344 22815
rect 4396 22763 4627 22815
rect 4103 22566 4637 22763
rect 4683 22566 4718 24550
rect 4826 24550 4942 25006
rect 5691 25002 6171 25006
rect 5691 24890 6091 25002
rect 5050 24854 6091 24890
rect 5050 24813 5084 24854
rect 4826 24456 4861 24550
rect 4022 22509 4718 22566
rect 4022 22463 4057 22509
rect 4103 22463 4637 22509
rect 4683 22463 4718 22509
rect 4022 22406 4718 22463
rect 4022 22360 4057 22406
rect 4103 22360 4637 22406
rect 4683 22360 4718 22406
rect 4022 22303 4718 22360
rect 4022 22257 4057 22303
rect 4103 22257 4637 22303
rect 4683 22257 4718 22303
rect 4022 22200 4718 22257
rect 4022 22154 4057 22200
rect 4103 22154 4637 22200
rect 4683 22154 4718 22200
rect 4022 22097 4718 22154
rect 4022 22051 4057 22097
rect 4103 22051 4637 22097
rect 4683 22051 4718 22097
rect 4022 21994 4718 22051
rect 4022 21948 4057 21994
rect 4103 21989 4637 21994
rect 4103 21948 4347 21989
rect 4022 21891 4347 21948
rect 3879 21845 3919 21882
rect 3795 21842 3919 21845
rect 3795 21790 3831 21842
rect 3883 21790 3919 21842
rect 3795 21788 3919 21790
rect 3795 21742 3833 21788
rect 3879 21742 3919 21788
rect 3795 21685 3919 21742
rect 3795 21639 3833 21685
rect 3879 21639 3919 21685
rect 3795 21624 3919 21639
rect 3795 21572 3831 21624
rect 3883 21572 3919 21624
rect 3795 21536 3833 21572
rect 3879 21536 3919 21572
rect 3795 21532 3919 21536
rect 4022 21845 4057 21891
rect 4103 21845 4347 21891
rect 4022 21788 4347 21845
rect 4022 21742 4057 21788
rect 4103 21742 4347 21788
rect 4022 21685 4347 21742
rect 4022 21639 4057 21685
rect 4103 21661 4347 21685
rect 4393 21948 4637 21989
rect 4683 21948 4718 21994
rect 4393 21891 4718 21948
rect 4393 21845 4637 21891
rect 4683 21845 4718 21891
rect 4907 24456 4942 24550
rect 5041 24808 5084 24813
rect 5130 24808 5243 24854
rect 5289 24808 5726 24854
rect 5772 24808 6091 24854
rect 5041 24773 6091 24808
rect 6137 24843 6171 25002
rect 6280 25002 6395 25135
rect 6137 24842 6175 24843
rect 6137 24802 6184 24842
rect 5041 24721 5079 24773
rect 5131 24771 6091 24773
rect 5131 24721 5169 24771
rect 5041 24556 5169 24721
rect 5041 24504 5079 24556
rect 5041 24338 5085 24504
rect 5041 24286 5079 24338
rect 5041 24121 5085 24286
rect 5041 24069 5079 24121
rect 5041 23903 5085 24069
rect 5041 23851 5079 23903
rect 5041 23685 5085 23851
rect 5041 23633 5079 23685
rect 5041 23467 5085 23633
rect 5041 23415 5079 23467
rect 5041 23250 5085 23415
rect 5041 23198 5079 23250
rect 5041 23032 5085 23198
rect 5041 22980 5079 23032
rect 5041 22815 5085 22980
rect 5041 22763 5079 22815
rect 5041 22722 5085 22763
rect 4861 22509 4907 22566
rect 4861 22406 4907 22463
rect 4861 22303 4907 22360
rect 4861 22200 4907 22257
rect 4861 22097 4907 22154
rect 4861 21994 4907 22051
rect 4861 21891 4907 21948
rect 4393 21788 4718 21845
rect 4393 21742 4637 21788
rect 4683 21742 4718 21788
rect 4393 21685 4718 21742
rect 4393 21661 4637 21685
rect 4103 21639 4637 21661
rect 4683 21639 4718 21685
rect 4022 21582 4718 21639
rect 4022 21536 4057 21582
rect 4103 21536 4637 21582
rect 4683 21536 4718 21582
rect 3833 21523 3879 21532
rect 4022 21531 4718 21536
rect 4821 21845 4861 21882
rect 5131 22722 5169 24556
rect 5691 24690 6091 24771
rect 6146 24750 6184 24802
rect 5691 24644 5726 24690
rect 5772 24644 6091 24690
rect 5691 24527 6091 24644
rect 6137 24585 6184 24750
rect 6280 24668 6315 25002
rect 6146 24533 6184 24585
rect 5691 24481 5726 24527
rect 5772 24481 6091 24527
rect 5691 24364 6091 24481
rect 6137 24367 6184 24533
rect 5691 24318 5726 24364
rect 5772 24318 6091 24364
rect 5691 24201 6091 24318
rect 6146 24315 6184 24367
rect 5691 24155 5726 24201
rect 5772 24155 6091 24201
rect 5691 24037 6091 24155
rect 6137 24150 6184 24315
rect 6146 24098 6184 24150
rect 5691 23991 5726 24037
rect 5772 23991 6091 24037
rect 5691 23874 6091 23991
rect 6137 23932 6184 24098
rect 6146 23880 6184 23932
rect 5691 23828 5726 23874
rect 5772 23828 6091 23874
rect 5691 23711 6091 23828
rect 6137 23714 6184 23880
rect 5691 23665 5726 23711
rect 5772 23665 6091 23711
rect 5691 23548 6091 23665
rect 6146 23662 6184 23714
rect 5691 23502 5726 23548
rect 5772 23502 6091 23548
rect 5691 23384 6091 23502
rect 6137 23496 6184 23662
rect 6146 23444 6184 23496
rect 5691 23338 5726 23384
rect 5772 23338 6091 23384
rect 5691 23221 6091 23338
rect 6137 23279 6184 23444
rect 6146 23227 6184 23279
rect 5691 23175 5726 23221
rect 5772 23175 6091 23221
rect 5691 23058 6091 23175
rect 6137 23061 6184 23227
rect 5691 23012 5726 23058
rect 5772 23012 6091 23058
rect 5691 22894 6091 23012
rect 6146 23009 6184 23061
rect 5691 22848 5726 22894
rect 5772 22848 6091 22894
rect 5691 22731 6091 22848
rect 6137 22844 6184 23009
rect 6146 22792 6184 22844
rect 5085 22509 5131 22566
rect 5085 22406 5131 22463
rect 5085 22303 5131 22360
rect 5085 22200 5131 22257
rect 5085 22097 5131 22154
rect 5085 21994 5131 22051
rect 5085 21891 5131 21948
rect 4907 21845 4945 21882
rect 4821 21842 4945 21845
rect 4821 21790 4857 21842
rect 4909 21790 4945 21842
rect 4821 21788 4945 21790
rect 4821 21742 4861 21788
rect 4907 21742 4945 21788
rect 4821 21685 4945 21742
rect 4821 21639 4861 21685
rect 4907 21639 4945 21685
rect 4821 21624 4945 21639
rect 4821 21572 4857 21624
rect 4909 21572 4945 21624
rect 4821 21536 4861 21572
rect 4907 21536 4945 21572
rect 4821 21532 4945 21536
rect 5085 21788 5131 21845
rect 5085 21685 5131 21742
rect 5085 21582 5131 21639
rect 4057 21523 4103 21531
rect 4637 21523 4683 21531
rect 4861 21523 4907 21532
rect 5085 21523 5131 21536
rect 5691 22685 5726 22731
rect 5772 22685 6091 22731
rect 5691 22568 6091 22685
rect 5691 22522 5726 22568
rect 5772 22522 6091 22568
rect 5691 22405 6091 22522
rect 5691 22359 5726 22405
rect 5772 22359 6091 22405
rect 5691 22241 6091 22359
rect 5691 22195 5726 22241
rect 5772 22195 6091 22241
rect 5691 22078 6091 22195
rect 5691 22032 5726 22078
rect 5772 22032 6091 22078
rect 5691 21915 6091 22032
rect 5691 21869 5726 21915
rect 5772 21869 6091 21915
rect 5691 21752 6091 21869
rect 5691 21706 5726 21752
rect 5772 21706 6091 21752
rect 5691 21588 6091 21706
rect 5691 21542 5726 21588
rect 5772 21542 6091 21588
rect 5691 21490 6091 21542
rect 6137 22751 6184 22792
rect 6137 21490 6171 22751
rect 5691 21486 6171 21490
rect 6273 21796 6315 21837
rect 6361 24668 6395 25002
rect 6605 25003 6651 25016
rect 6571 23427 6605 24851
rect 6829 25003 6875 25428
rect 7430 26382 7782 26462
rect 7430 26336 7478 26382
rect 7524 26379 7782 26382
rect 7828 26379 7862 26643
rect 7524 26336 7862 26379
rect 7430 26322 7862 26336
rect 7430 26296 7782 26322
rect 7430 26244 7565 26296
rect 7617 26244 7772 26296
rect 7828 26276 7862 26322
rect 7824 26244 7862 26276
rect 7430 26219 7862 26244
rect 7430 26218 7782 26219
rect 7430 26172 7478 26218
rect 7524 26173 7782 26218
rect 7828 26173 7862 26219
rect 7524 26172 7862 26173
rect 7430 26116 7862 26172
rect 7430 26078 7782 26116
rect 7430 26055 7565 26078
rect 7430 26009 7478 26055
rect 7524 26026 7565 26055
rect 7617 26026 7772 26078
rect 7828 26070 7862 26116
rect 7824 26026 7862 26070
rect 7524 26013 7862 26026
rect 7524 26009 7782 26013
rect 7430 25967 7782 26009
rect 7828 25967 7862 26013
rect 7430 25910 7862 25967
rect 7430 25892 7782 25910
rect 7430 25846 7478 25892
rect 7524 25864 7782 25892
rect 7828 25864 7862 25910
rect 7524 25860 7862 25864
rect 7524 25846 7565 25860
rect 7430 25808 7565 25846
rect 7617 25808 7772 25860
rect 7824 25808 7862 25860
rect 7430 25807 7862 25808
rect 7430 25761 7782 25807
rect 7828 25761 7862 25807
rect 7430 25728 7862 25761
rect 7430 25682 7478 25728
rect 7524 25704 7862 25728
rect 7524 25682 7782 25704
rect 7430 25658 7782 25682
rect 7828 25658 7862 25704
rect 7430 25601 7862 25658
rect 7430 25565 7782 25601
rect 7430 25519 7478 25565
rect 7524 25555 7782 25565
rect 7828 25555 7862 25601
rect 7524 25519 7862 25555
rect 7430 25498 7862 25519
rect 7430 25452 7782 25498
rect 7828 25452 7862 25498
rect 7430 25395 7862 25452
rect 9038 26717 9084 26776
rect 9038 26612 9084 26671
rect 8006 26322 8052 26379
rect 8006 26219 8052 26276
rect 8006 26116 8052 26173
rect 8006 26013 8052 26070
rect 8006 25910 8052 25967
rect 8006 25807 8052 25864
rect 8006 25704 8052 25761
rect 8254 26491 8382 26531
rect 8254 26439 8292 26491
rect 8344 26439 8382 26491
rect 9038 26507 9084 26566
rect 8254 26400 8296 26439
rect 8342 26400 8382 26439
rect 8254 26338 8382 26400
rect 8254 26292 8296 26338
rect 8342 26292 8382 26338
rect 8254 26273 8382 26292
rect 8254 26221 8292 26273
rect 8344 26221 8382 26273
rect 8254 26184 8296 26221
rect 8342 26184 8382 26221
rect 8254 26122 8382 26184
rect 8254 26076 8296 26122
rect 8342 26076 8382 26122
rect 8254 26055 8382 26076
rect 8254 26003 8292 26055
rect 8344 26003 8382 26055
rect 8254 25968 8296 26003
rect 8342 25968 8382 26003
rect 8254 25906 8382 25968
rect 8254 25860 8296 25906
rect 8342 25860 8382 25906
rect 8254 25837 8382 25860
rect 8254 25785 8292 25837
rect 8344 25785 8382 25837
rect 8254 25752 8296 25785
rect 8342 25752 8382 25785
rect 8254 25745 8382 25752
rect 8520 26446 8566 26459
rect 8520 26338 8566 26400
rect 8520 26230 8566 26292
rect 8520 26122 8566 26184
rect 8520 26014 8566 26076
rect 8520 25906 8566 25968
rect 8520 25798 8566 25860
rect 8006 25601 8052 25658
rect 8006 25498 8052 25555
rect 8006 25405 8052 25452
rect 8296 25690 8342 25745
rect 8296 25582 8342 25644
rect 8296 25474 8342 25536
rect 8296 25415 8342 25428
rect 8520 25690 8566 25752
rect 8520 25582 8566 25644
rect 8520 25474 8566 25536
rect 7430 25349 7782 25395
rect 7828 25349 7862 25395
rect 7430 25344 7862 25349
rect 7971 25395 8086 25405
rect 7971 25349 8006 25395
rect 8052 25349 8086 25395
rect 7782 25336 7828 25344
rect 7527 25255 7867 25262
rect 7971 25255 8086 25349
rect 7527 25221 7884 25255
rect 7527 25169 7565 25221
rect 7617 25218 7777 25221
rect 7829 25218 7884 25221
rect 7617 25172 7645 25218
rect 7691 25172 7777 25218
rect 7849 25172 7884 25218
rect 7617 25169 7777 25172
rect 7829 25169 7884 25172
rect 7527 25135 7884 25169
rect 7971 25218 8394 25255
rect 7971 25172 8155 25218
rect 8201 25172 8313 25218
rect 8359 25172 8394 25218
rect 7971 25135 8394 25172
rect 7527 25129 7867 25135
rect 7782 25006 7828 25015
rect 6651 24811 6698 24851
rect 6660 24759 6698 24811
rect 6651 24593 6698 24759
rect 6660 24541 6698 24593
rect 6651 24376 6698 24541
rect 6660 24324 6698 24376
rect 6651 24158 6698 24324
rect 6660 24106 6698 24158
rect 6651 23940 6698 24106
rect 6660 23888 6698 23940
rect 6651 23722 6698 23888
rect 6660 23670 6698 23722
rect 6651 23505 6698 23670
rect 6660 23453 6698 23505
rect 6651 23427 6698 23453
rect 6571 23370 6698 23427
rect 6571 23324 6605 23370
rect 6651 23324 6698 23370
rect 6571 23287 6698 23324
rect 6571 23267 6608 23287
rect 6571 23221 6605 23267
rect 6660 23235 6698 23287
rect 6651 23221 6698 23235
rect 6571 23195 6698 23221
rect 6829 23370 6875 23427
rect 6829 23267 6875 23324
rect 6605 23164 6651 23195
rect 6605 23061 6651 23118
rect 6605 22958 6651 23015
rect 6605 22855 6651 22912
rect 6605 22752 6651 22809
rect 6829 23164 6875 23221
rect 6829 23061 6875 23118
rect 6829 22958 6875 23015
rect 6829 22855 6875 22912
rect 6829 22752 6875 22809
rect 6605 22649 6651 22706
rect 6605 22546 6651 22603
rect 6605 22443 6651 22500
rect 6605 22384 6651 22397
rect 6789 22706 6829 22743
rect 7382 25002 7862 25006
rect 7382 24854 7782 25002
rect 7382 24808 7417 24854
rect 7463 24808 7782 24854
rect 7382 24690 7782 24808
rect 7828 24843 7862 25002
rect 7971 25002 8086 25135
rect 7828 24842 7866 24843
rect 7828 24802 7875 24842
rect 7837 24750 7875 24802
rect 7382 24644 7417 24690
rect 7463 24644 7782 24690
rect 7382 24527 7782 24644
rect 7828 24585 7875 24750
rect 7971 24668 8006 25002
rect 7837 24533 7875 24585
rect 7382 24481 7417 24527
rect 7463 24481 7782 24527
rect 7382 24364 7782 24481
rect 7828 24367 7875 24533
rect 7382 24318 7417 24364
rect 7463 24318 7782 24364
rect 7382 24201 7782 24318
rect 7837 24315 7875 24367
rect 7382 24155 7417 24201
rect 7463 24155 7782 24201
rect 7382 24037 7782 24155
rect 7828 24150 7875 24315
rect 7837 24098 7875 24150
rect 7382 23991 7417 24037
rect 7463 23991 7782 24037
rect 7382 23874 7782 23991
rect 7828 23932 7875 24098
rect 7837 23880 7875 23932
rect 7382 23828 7417 23874
rect 7463 23828 7782 23874
rect 7382 23711 7782 23828
rect 7828 23714 7875 23880
rect 7382 23665 7417 23711
rect 7463 23665 7782 23711
rect 7382 23548 7782 23665
rect 7837 23662 7875 23714
rect 7382 23502 7417 23548
rect 7463 23502 7782 23548
rect 7382 23384 7782 23502
rect 7828 23496 7875 23662
rect 7837 23444 7875 23496
rect 7382 23338 7417 23384
rect 7463 23338 7782 23384
rect 7382 23221 7782 23338
rect 7828 23279 7875 23444
rect 7837 23227 7875 23279
rect 7382 23175 7417 23221
rect 7463 23175 7782 23221
rect 7382 23058 7782 23175
rect 7828 23061 7875 23227
rect 7382 23012 7417 23058
rect 7463 23012 7782 23058
rect 7382 22894 7782 23012
rect 7837 23009 7875 23061
rect 7382 22848 7417 22894
rect 7463 22848 7782 22894
rect 6875 22706 6913 22743
rect 6789 22703 6913 22706
rect 6789 22651 6825 22703
rect 6877 22651 6913 22703
rect 6789 22649 6913 22651
rect 6789 22603 6829 22649
rect 6875 22603 6913 22649
rect 6789 22546 6913 22603
rect 6789 22500 6829 22546
rect 6875 22500 6913 22546
rect 6789 22485 6913 22500
rect 6789 22433 6825 22485
rect 6877 22433 6913 22485
rect 6789 22397 6829 22433
rect 6875 22397 6913 22433
rect 6789 22393 6913 22397
rect 7382 22731 7782 22848
rect 7828 22844 7875 23009
rect 7837 22792 7875 22844
rect 7382 22685 7417 22731
rect 7463 22685 7782 22731
rect 7382 22568 7782 22685
rect 7382 22522 7417 22568
rect 7463 22522 7782 22568
rect 7382 22405 7782 22522
rect 6829 22384 6875 22393
rect 7382 22359 7417 22405
rect 7463 22359 7782 22405
rect 7382 22241 7782 22359
rect 7382 22195 7417 22241
rect 7463 22195 7782 22241
rect 7382 22078 7782 22195
rect 7382 22032 7417 22078
rect 7463 22032 7782 22078
rect 7382 21915 7782 22032
rect 7382 21869 7417 21915
rect 7463 21869 7782 21915
rect 6361 21796 6402 21837
rect 6273 21744 6311 21796
rect 6363 21744 6402 21796
rect 6273 21578 6315 21744
rect 6361 21578 6402 21744
rect 6273 21526 6311 21578
rect 6363 21526 6402 21578
rect 6273 21490 6315 21526
rect 6361 21490 6402 21526
rect 6091 21477 6137 21486
rect 1894 21383 2009 21399
rect 3146 21383 3261 21399
rect 6273 21383 6402 21490
rect 7382 21752 7782 21869
rect 7382 21706 7417 21752
rect 7463 21706 7782 21752
rect 7382 21588 7782 21706
rect 7382 21542 7417 21588
rect 7463 21542 7782 21588
rect 7382 21490 7782 21542
rect 7828 22751 7875 22792
rect 7828 21490 7862 22751
rect 7382 21486 7862 21490
rect 7966 21796 8006 21836
rect 8052 24668 8086 25002
rect 8296 25003 8342 25016
rect 8262 23427 8296 24851
rect 8520 25003 8566 25428
rect 9038 26402 9084 26461
rect 9038 26297 9084 26356
rect 9038 26192 9084 26251
rect 9038 26088 9084 26146
rect 9038 25984 9084 26042
rect 9038 25880 9084 25938
rect 9038 25776 9084 25834
rect 9038 25672 9084 25730
rect 9038 25568 9084 25626
rect 9038 25464 9084 25522
rect 9038 25360 9084 25418
rect 9038 25256 9084 25314
rect 9038 25197 9084 25210
rect 9262 26822 9308 26881
rect 9445 27353 9573 27392
rect 9445 27301 9483 27353
rect 9535 27301 9573 27353
rect 9445 27242 9573 27301
rect 9445 27196 9486 27242
rect 9532 27196 9573 27242
rect 9445 27137 9573 27196
rect 9445 27135 9486 27137
rect 9532 27135 9573 27137
rect 9445 27083 9483 27135
rect 9535 27083 9573 27135
rect 9445 27032 9573 27083
rect 9445 26986 9486 27032
rect 9532 26986 9573 27032
rect 9445 26927 9573 26986
rect 9445 26917 9486 26927
rect 9532 26917 9573 26927
rect 9445 26865 9483 26917
rect 9535 26865 9573 26917
rect 9445 26825 9573 26865
rect 9710 27347 9756 27396
rect 9934 27392 9980 27406
rect 10123 27452 10239 27546
rect 10123 27406 10158 27452
rect 10204 27406 10239 27452
rect 10123 27396 10239 27406
rect 10382 27452 10428 27465
rect 9710 27242 9756 27301
rect 9710 27137 9756 27196
rect 9710 27032 9756 27091
rect 9710 26927 9756 26986
rect 9262 26717 9308 26776
rect 9262 26612 9308 26671
rect 9262 26507 9308 26566
rect 9262 26402 9308 26461
rect 9262 26297 9308 26356
rect 9262 26192 9308 26251
rect 9262 26088 9308 26146
rect 9262 25984 9308 26042
rect 9262 25880 9308 25938
rect 9262 25776 9308 25834
rect 9262 25672 9308 25730
rect 9262 25568 9308 25626
rect 9262 25464 9308 25522
rect 9262 25360 9308 25418
rect 9262 25256 9308 25314
rect 9262 25197 9308 25210
rect 9486 26822 9532 26825
rect 9486 26717 9532 26776
rect 9486 26612 9532 26671
rect 9486 26507 9532 26566
rect 9486 26402 9532 26461
rect 9486 26297 9532 26356
rect 9486 26192 9532 26251
rect 9486 26088 9532 26146
rect 9486 25984 9532 26042
rect 9486 25880 9532 25938
rect 9486 25776 9532 25834
rect 9486 25672 9532 25730
rect 9486 25568 9532 25626
rect 9486 25464 9532 25522
rect 9486 25360 9532 25418
rect 9486 25256 9532 25314
rect 9486 25197 9532 25210
rect 9710 26822 9756 26881
rect 9893 27353 10021 27392
rect 9893 27301 9931 27353
rect 9983 27301 10021 27353
rect 9893 27242 10021 27301
rect 9893 27196 9934 27242
rect 9980 27196 10021 27242
rect 9893 27137 10021 27196
rect 9893 27135 9934 27137
rect 9980 27135 10021 27137
rect 9893 27083 9931 27135
rect 9983 27083 10021 27135
rect 9893 27032 10021 27083
rect 9893 26986 9934 27032
rect 9980 26986 10021 27032
rect 9893 26927 10021 26986
rect 9893 26917 9934 26927
rect 9980 26917 10021 26927
rect 9893 26865 9931 26917
rect 9983 26865 10021 26917
rect 9893 26825 10021 26865
rect 10158 27347 10204 27396
rect 10382 27392 10428 27406
rect 10571 27452 10687 27546
rect 11019 27665 11135 27758
rect 11229 27794 11267 27846
rect 11319 27804 11357 27846
rect 11229 27758 11278 27794
rect 11324 27758 11357 27804
rect 11229 27754 11357 27758
rect 11461 28535 11589 28540
rect 11691 28539 11807 28594
rect 11950 28640 11996 28653
rect 11950 28540 11996 28594
rect 12139 28640 12255 28939
rect 12587 28934 12780 28939
rect 12826 28934 12938 28980
rect 12984 28934 13096 28980
rect 13142 28934 13254 28980
rect 13300 28934 13412 28980
rect 13458 28934 13570 28980
rect 13616 28934 13728 28980
rect 13774 28934 13886 28980
rect 13932 28934 14045 28980
rect 14091 28934 14203 28980
rect 14249 28934 14361 28980
rect 14407 28934 14519 28980
rect 14565 28934 14677 28980
rect 14723 28934 14835 28980
rect 14881 28934 14993 28980
rect 15039 28934 15152 28980
rect 15198 28934 15310 28980
rect 15356 28934 15468 28980
rect 15514 28934 15626 28980
rect 15672 28934 15784 28980
rect 15830 28934 15942 28980
rect 15988 28934 16100 28980
rect 16146 28934 16258 28980
rect 16304 28934 16416 28980
rect 16462 28934 16497 28980
rect 12587 28897 16497 28934
rect 29520 28996 29654 29037
rect 29520 28944 29561 28996
rect 29613 28944 29654 28996
rect 12139 28594 12174 28640
rect 12220 28594 12255 28640
rect 12139 28540 12255 28594
rect 12398 28640 12444 28653
rect 11461 28500 11502 28535
rect 11548 28500 11589 28535
rect 11461 28448 11499 28500
rect 11551 28448 11589 28500
rect 11461 28430 11589 28448
rect 11461 28384 11502 28430
rect 11548 28384 11589 28430
rect 11461 28325 11589 28384
rect 11461 28282 11502 28325
rect 11548 28282 11589 28325
rect 11461 28230 11499 28282
rect 11551 28230 11589 28282
rect 11461 28220 11589 28230
rect 11461 28174 11502 28220
rect 11548 28174 11589 28220
rect 11461 28116 11589 28174
rect 11461 28070 11502 28116
rect 11548 28070 11589 28116
rect 11461 28064 11589 28070
rect 11461 28012 11499 28064
rect 11551 28012 11589 28064
rect 11461 27966 11502 28012
rect 11548 27966 11589 28012
rect 11461 27908 11589 27966
rect 11461 27862 11502 27908
rect 11548 27862 11589 27908
rect 11461 27846 11589 27862
rect 11461 27794 11499 27846
rect 11551 27794 11589 27846
rect 11461 27758 11502 27794
rect 11548 27758 11589 27794
rect 11461 27754 11589 27758
rect 11726 28535 11772 28539
rect 11726 28430 11772 28489
rect 11726 28325 11772 28384
rect 11726 28220 11772 28279
rect 11726 28116 11772 28174
rect 11726 28012 11772 28070
rect 11726 27908 11772 27966
rect 11726 27804 11772 27862
rect 11278 27745 11324 27754
rect 11467 27665 11583 27754
rect 11726 27745 11772 27758
rect 11909 28535 12037 28540
rect 12139 28539 12269 28540
rect 11909 28500 11950 28535
rect 11996 28500 12037 28535
rect 11909 28448 11947 28500
rect 11999 28448 12037 28500
rect 11909 28430 12037 28448
rect 11909 28384 11950 28430
rect 11996 28384 12037 28430
rect 11909 28325 12037 28384
rect 11909 28282 11950 28325
rect 11996 28282 12037 28325
rect 11909 28230 11947 28282
rect 11999 28230 12037 28282
rect 11909 28220 12037 28230
rect 11909 28174 11950 28220
rect 11996 28174 12037 28220
rect 11909 28116 12037 28174
rect 11909 28070 11950 28116
rect 11996 28070 12037 28116
rect 11909 28064 12037 28070
rect 11909 28012 11947 28064
rect 11999 28012 12037 28064
rect 11909 27966 11950 28012
rect 11996 27966 12037 28012
rect 11909 27908 12037 27966
rect 11909 27862 11950 27908
rect 11996 27862 12037 27908
rect 11909 27846 12037 27862
rect 11909 27794 11947 27846
rect 11999 27794 12037 27846
rect 11909 27758 11950 27794
rect 11996 27758 12037 27794
rect 11909 27754 12037 27758
rect 12141 28535 12269 28539
rect 12141 28489 12174 28535
rect 12220 28500 12269 28535
rect 12141 28448 12179 28489
rect 12231 28448 12269 28500
rect 12141 28430 12269 28448
rect 12141 28384 12174 28430
rect 12220 28384 12269 28430
rect 12141 28325 12269 28384
rect 12141 28279 12174 28325
rect 12220 28282 12269 28325
rect 12141 28230 12179 28279
rect 12231 28230 12269 28282
rect 12141 28220 12269 28230
rect 12141 28174 12174 28220
rect 12220 28174 12269 28220
rect 12141 28116 12269 28174
rect 12141 28070 12174 28116
rect 12220 28070 12269 28116
rect 12141 28064 12269 28070
rect 12141 28012 12179 28064
rect 12231 28012 12269 28064
rect 12141 27966 12174 28012
rect 12220 27966 12269 28012
rect 12141 27908 12269 27966
rect 12141 27862 12174 27908
rect 12220 27862 12269 27908
rect 12141 27846 12269 27862
rect 12141 27804 12179 27846
rect 12141 27758 12174 27804
rect 12231 27794 12269 27846
rect 12398 28535 12444 28594
rect 12587 28640 12703 28897
rect 12587 28594 12622 28640
rect 12668 28594 12703 28640
rect 12587 28540 12703 28594
rect 13276 28896 13393 28897
rect 12398 28430 12444 28489
rect 12398 28325 12444 28384
rect 12398 28220 12444 28279
rect 12398 28116 12444 28174
rect 12398 28012 12444 28070
rect 12398 27908 12444 27966
rect 12398 27804 12444 27862
rect 12220 27758 12269 27794
rect 12141 27754 12269 27758
rect 12363 27758 12398 27795
rect 12581 28535 12709 28540
rect 12581 28500 12622 28535
rect 12668 28500 12709 28535
rect 12581 28448 12619 28500
rect 12671 28448 12709 28500
rect 12581 28430 12709 28448
rect 13276 28440 13392 28896
rect 13724 28440 13840 28897
rect 12581 28384 12622 28430
rect 12668 28384 12709 28430
rect 12581 28325 12709 28384
rect 12581 28282 12622 28325
rect 12668 28282 12709 28325
rect 12581 28230 12619 28282
rect 12671 28230 12709 28282
rect 12581 28220 12709 28230
rect 12581 28174 12622 28220
rect 12668 28174 12709 28220
rect 12581 28116 12709 28174
rect 12581 28070 12622 28116
rect 12668 28070 12709 28116
rect 12581 28064 12709 28070
rect 12581 28012 12619 28064
rect 12671 28012 12709 28064
rect 12581 27966 12622 28012
rect 12668 27966 12709 28012
rect 12581 27908 12709 27966
rect 12581 27862 12622 27908
rect 12668 27862 12709 27908
rect 13264 28401 13392 28440
rect 13264 28349 13302 28401
rect 13354 28349 13392 28401
rect 13264 28183 13392 28349
rect 13264 28131 13302 28183
rect 13354 28131 13392 28183
rect 13703 28401 13840 28440
rect 13703 28349 13741 28401
rect 13793 28349 13840 28401
rect 15095 28896 15211 28897
rect 15095 28384 15210 28896
rect 29520 28778 29654 28944
rect 29520 28726 29561 28778
rect 29613 28726 29654 28778
rect 16581 28411 28525 28461
rect 15095 28383 15211 28384
rect 13703 28183 13840 28349
rect 15087 28344 15215 28383
rect 15087 28292 15125 28344
rect 15177 28292 15215 28344
rect 13264 28082 13392 28131
rect 13264 27965 13312 28082
rect 13264 27913 13302 27965
rect 13264 27873 13312 27913
rect 12581 27846 12709 27862
rect 12444 27758 12479 27795
rect 11019 27546 11583 27665
rect 10571 27406 10606 27452
rect 10652 27406 10687 27452
rect 10571 27396 10687 27406
rect 10830 27452 10876 27465
rect 10158 27242 10204 27301
rect 10158 27137 10204 27196
rect 10158 27032 10204 27091
rect 10158 26927 10204 26986
rect 9710 26717 9756 26776
rect 9710 26612 9756 26671
rect 9710 26507 9756 26566
rect 9710 26402 9756 26461
rect 9710 26297 9756 26356
rect 9710 26192 9756 26251
rect 9710 26088 9756 26146
rect 9710 25984 9756 26042
rect 9710 25880 9756 25938
rect 9710 25776 9756 25834
rect 9710 25672 9756 25730
rect 9710 25568 9756 25626
rect 9710 25464 9756 25522
rect 9710 25360 9756 25418
rect 9710 25256 9756 25314
rect 9710 25197 9756 25210
rect 9934 26822 9980 26825
rect 9934 26717 9980 26776
rect 9934 26612 9980 26671
rect 9934 26507 9980 26566
rect 9934 26402 9980 26461
rect 9934 26297 9980 26356
rect 9934 26192 9980 26251
rect 9934 26088 9980 26146
rect 9934 25984 9980 26042
rect 9934 25880 9980 25938
rect 9934 25776 9980 25834
rect 9934 25672 9980 25730
rect 9934 25568 9980 25626
rect 9934 25464 9980 25522
rect 9934 25360 9980 25418
rect 9934 25256 9980 25314
rect 9934 25197 9980 25210
rect 10158 26822 10204 26881
rect 10341 27353 10469 27392
rect 10341 27301 10379 27353
rect 10431 27301 10469 27353
rect 10341 27242 10469 27301
rect 10341 27196 10382 27242
rect 10428 27196 10469 27242
rect 10341 27137 10469 27196
rect 10341 27135 10382 27137
rect 10428 27135 10469 27137
rect 10341 27083 10379 27135
rect 10431 27083 10469 27135
rect 10341 27032 10469 27083
rect 10341 26986 10382 27032
rect 10428 26986 10469 27032
rect 10341 26927 10469 26986
rect 10341 26917 10382 26927
rect 10428 26917 10469 26927
rect 10341 26865 10379 26917
rect 10431 26865 10469 26917
rect 10341 26825 10469 26865
rect 10606 27347 10652 27396
rect 10830 27392 10876 27406
rect 11019 27452 11135 27546
rect 11019 27406 11054 27452
rect 11100 27406 11135 27452
rect 11019 27396 11135 27406
rect 11278 27452 11324 27465
rect 10606 27242 10652 27301
rect 10606 27137 10652 27196
rect 10606 27032 10652 27091
rect 10606 26927 10652 26986
rect 10158 26717 10204 26776
rect 10158 26612 10204 26671
rect 10158 26507 10204 26566
rect 10158 26402 10204 26461
rect 10158 26297 10204 26356
rect 10158 26192 10204 26251
rect 10158 26088 10204 26146
rect 10158 25984 10204 26042
rect 10158 25880 10204 25938
rect 10158 25776 10204 25834
rect 10158 25672 10204 25730
rect 10158 25568 10204 25626
rect 10158 25464 10204 25522
rect 10158 25360 10204 25418
rect 10158 25256 10204 25314
rect 10158 25197 10204 25210
rect 10382 26822 10428 26825
rect 10382 26717 10428 26776
rect 10382 26612 10428 26671
rect 10382 26507 10428 26566
rect 10382 26402 10428 26461
rect 10382 26297 10428 26356
rect 10382 26192 10428 26251
rect 10382 26088 10428 26146
rect 10382 25984 10428 26042
rect 10382 25880 10428 25938
rect 10382 25776 10428 25834
rect 10382 25672 10428 25730
rect 10382 25568 10428 25626
rect 10382 25464 10428 25522
rect 10382 25360 10428 25418
rect 10382 25256 10428 25314
rect 10382 25197 10428 25210
rect 10606 26822 10652 26881
rect 10789 27353 10917 27392
rect 10789 27301 10827 27353
rect 10879 27301 10917 27353
rect 10789 27242 10917 27301
rect 10789 27196 10830 27242
rect 10876 27196 10917 27242
rect 10789 27137 10917 27196
rect 10789 27135 10830 27137
rect 10876 27135 10917 27137
rect 10789 27083 10827 27135
rect 10879 27083 10917 27135
rect 10789 27032 10917 27083
rect 10789 26986 10830 27032
rect 10876 26986 10917 27032
rect 10789 26927 10917 26986
rect 10789 26917 10830 26927
rect 10876 26917 10917 26927
rect 10789 26865 10827 26917
rect 10879 26865 10917 26917
rect 10789 26825 10917 26865
rect 11054 27347 11100 27396
rect 11278 27392 11324 27406
rect 11467 27452 11583 27546
rect 11915 27665 12031 27754
rect 12174 27745 12220 27754
rect 12363 27665 12479 27758
rect 12581 27794 12619 27846
rect 12671 27794 12709 27846
rect 13276 27834 13312 27873
rect 13358 27834 13392 28082
rect 13276 27821 13392 27834
rect 13500 28082 13616 28135
rect 13500 27834 13536 28082
rect 13582 27834 13616 28082
rect 13703 28131 13741 28183
rect 13793 28131 13840 28183
rect 13703 28082 13840 28131
rect 13703 27965 13760 28082
rect 13703 27913 13741 27965
rect 13703 27873 13760 27913
rect 12581 27758 12622 27794
rect 12668 27758 12709 27794
rect 12581 27754 12709 27758
rect 12622 27745 12668 27754
rect 13500 27733 13616 27834
rect 13724 27834 13760 27873
rect 13806 27834 13840 28082
rect 13925 28185 14049 28225
rect 13925 28133 13961 28185
rect 14013 28133 14049 28185
rect 13925 28026 14049 28133
rect 13925 27967 13966 28026
rect 14012 27967 14049 28026
rect 15087 28126 15215 28292
rect 16581 28365 16812 28411
rect 16858 28392 16970 28411
rect 16858 28365 16918 28392
rect 16581 28340 16918 28365
rect 17016 28365 17128 28411
rect 17174 28365 17286 28411
rect 17332 28365 17466 28411
rect 17512 28365 17624 28411
rect 17670 28365 17782 28411
rect 17828 28392 17940 28411
rect 16970 28340 17828 28365
rect 17880 28365 17940 28392
rect 17986 28365 18446 28411
rect 18492 28392 18604 28411
rect 18492 28365 18552 28392
rect 17880 28340 18552 28365
rect 18650 28365 18762 28411
rect 18808 28365 18920 28411
rect 18966 28365 19100 28411
rect 19146 28365 19258 28411
rect 19304 28365 19416 28411
rect 19462 28392 19574 28411
rect 18604 28340 19462 28365
rect 19514 28365 19574 28392
rect 19620 28365 20079 28411
rect 20125 28392 20237 28411
rect 20125 28365 20185 28392
rect 19514 28340 20185 28365
rect 20283 28365 20395 28411
rect 20441 28365 20553 28411
rect 20599 28365 20733 28411
rect 20779 28365 20891 28411
rect 20937 28365 21049 28411
rect 21095 28392 21207 28411
rect 20237 28340 21095 28365
rect 21147 28365 21207 28392
rect 21253 28365 21713 28411
rect 21759 28392 21871 28411
rect 21759 28365 21819 28392
rect 21147 28340 21819 28365
rect 21917 28365 22029 28411
rect 22075 28365 22187 28411
rect 22233 28365 22367 28411
rect 22413 28365 22525 28411
rect 22571 28365 22683 28411
rect 22729 28392 22841 28411
rect 21871 28340 22729 28365
rect 22781 28365 22841 28392
rect 22887 28407 24726 28411
rect 22887 28365 23231 28407
rect 22781 28361 23231 28365
rect 24499 28365 24726 28407
rect 24772 28365 24884 28411
rect 24930 28365 25042 28411
rect 25088 28365 25200 28411
rect 25246 28365 25358 28411
rect 25404 28365 25516 28411
rect 25562 28365 25674 28411
rect 25720 28365 25833 28411
rect 25879 28365 25991 28411
rect 26037 28365 26149 28411
rect 26195 28365 26307 28411
rect 26353 28365 26465 28411
rect 26511 28365 26623 28411
rect 26669 28365 26781 28411
rect 26827 28365 26939 28411
rect 26985 28365 27097 28411
rect 27143 28365 27256 28411
rect 27302 28365 27414 28411
rect 27460 28365 27572 28411
rect 27618 28365 27730 28411
rect 27776 28365 27888 28411
rect 27934 28365 28046 28411
rect 28092 28365 28204 28411
rect 28250 28365 28362 28411
rect 28408 28365 28525 28411
rect 24499 28361 28525 28365
rect 22781 28349 23787 28361
rect 23839 28349 24226 28361
rect 24278 28349 28525 28361
rect 22781 28344 28525 28349
rect 22781 28340 25610 28344
rect 16581 28314 25610 28340
rect 16581 28174 23118 28314
rect 16581 28170 16918 28174
rect 15087 28074 15125 28126
rect 15177 28074 15215 28126
rect 16880 28122 16918 28170
rect 16970 28170 17828 28174
rect 16970 28122 17009 28170
rect 13925 27915 13961 27967
rect 14013 27915 14049 27967
rect 13925 27886 13966 27915
rect 14012 27886 14049 27915
rect 13925 27875 14049 27886
rect 14906 27996 14952 28009
rect 14906 27876 14952 27950
rect 13724 27821 13840 27834
rect 11915 27546 12479 27665
rect 13204 27683 13384 27695
rect 13204 27631 13216 27683
rect 13373 27637 13384 27683
rect 13372 27631 13384 27637
rect 13204 27619 13384 27631
rect 13500 27614 13840 27733
rect 14906 27702 14952 27830
rect 15087 27996 15215 28074
rect 15087 27950 15130 27996
rect 15176 27950 15215 27996
rect 15087 27908 15215 27950
rect 15087 27856 15125 27908
rect 15177 27856 15215 27908
rect 15087 27830 15130 27856
rect 15176 27830 15215 27856
rect 15087 27816 15215 27830
rect 16704 28076 16750 28089
rect 16704 27971 16750 28030
rect 16704 27866 16750 27925
rect 16704 27761 16750 27820
rect 16121 27702 16245 27735
rect 14906 27695 16247 27702
rect 14132 27683 14312 27695
rect 14132 27631 14144 27683
rect 14300 27631 14312 27683
rect 14132 27619 14312 27631
rect 11467 27406 11502 27452
rect 11548 27406 11583 27452
rect 11467 27396 11583 27406
rect 11726 27452 11772 27465
rect 11054 27242 11100 27301
rect 11054 27137 11100 27196
rect 11054 27032 11100 27091
rect 11054 26927 11100 26986
rect 10606 26717 10652 26776
rect 10606 26612 10652 26671
rect 10606 26507 10652 26566
rect 10606 26402 10652 26461
rect 10606 26297 10652 26356
rect 10606 26192 10652 26251
rect 10606 26088 10652 26146
rect 10606 25984 10652 26042
rect 10606 25880 10652 25938
rect 10606 25776 10652 25834
rect 10606 25672 10652 25730
rect 10606 25568 10652 25626
rect 10606 25464 10652 25522
rect 10606 25360 10652 25418
rect 10606 25256 10652 25314
rect 10606 25197 10652 25210
rect 10830 26822 10876 26825
rect 10830 26717 10876 26776
rect 10830 26612 10876 26671
rect 10830 26507 10876 26566
rect 10830 26402 10876 26461
rect 10830 26297 10876 26356
rect 10830 26192 10876 26251
rect 10830 26088 10876 26146
rect 10830 25984 10876 26042
rect 10830 25880 10876 25938
rect 10830 25776 10876 25834
rect 10830 25672 10876 25730
rect 10830 25568 10876 25626
rect 10830 25464 10876 25522
rect 10830 25360 10876 25418
rect 10830 25256 10876 25314
rect 10830 25197 10876 25210
rect 11054 26822 11100 26881
rect 11237 27353 11365 27392
rect 11237 27301 11275 27353
rect 11327 27301 11365 27353
rect 11237 27242 11365 27301
rect 11237 27196 11278 27242
rect 11324 27196 11365 27242
rect 11237 27137 11365 27196
rect 11237 27135 11278 27137
rect 11324 27135 11365 27137
rect 11237 27083 11275 27135
rect 11327 27083 11365 27135
rect 11237 27032 11365 27083
rect 11237 26986 11278 27032
rect 11324 26986 11365 27032
rect 11237 26927 11365 26986
rect 11237 26917 11278 26927
rect 11324 26917 11365 26927
rect 11237 26865 11275 26917
rect 11327 26865 11365 26917
rect 11237 26825 11365 26865
rect 11502 27347 11548 27396
rect 11726 27392 11772 27406
rect 11915 27452 12031 27546
rect 11915 27406 11950 27452
rect 11996 27406 12031 27452
rect 11915 27396 12031 27406
rect 12174 27452 12220 27465
rect 11502 27242 11548 27301
rect 11502 27137 11548 27196
rect 11502 27032 11548 27091
rect 11502 26927 11548 26986
rect 11054 26717 11100 26776
rect 11054 26612 11100 26671
rect 11054 26507 11100 26566
rect 11054 26402 11100 26461
rect 11054 26297 11100 26356
rect 11054 26192 11100 26251
rect 11054 26088 11100 26146
rect 11054 25984 11100 26042
rect 11054 25880 11100 25938
rect 11054 25776 11100 25834
rect 11054 25672 11100 25730
rect 11054 25568 11100 25626
rect 11054 25464 11100 25522
rect 11054 25360 11100 25418
rect 11054 25256 11100 25314
rect 11054 25197 11100 25210
rect 11278 26822 11324 26825
rect 11278 26717 11324 26776
rect 11278 26612 11324 26671
rect 11278 26507 11324 26566
rect 11278 26402 11324 26461
rect 11278 26297 11324 26356
rect 11278 26192 11324 26251
rect 11278 26088 11324 26146
rect 11278 25984 11324 26042
rect 11278 25880 11324 25938
rect 11278 25776 11324 25834
rect 11278 25672 11324 25730
rect 11278 25568 11324 25626
rect 11278 25464 11324 25522
rect 11278 25360 11324 25418
rect 11278 25256 11324 25314
rect 11278 25197 11324 25210
rect 11502 26822 11548 26881
rect 11685 27353 11813 27392
rect 11685 27301 11723 27353
rect 11775 27301 11813 27353
rect 11685 27242 11813 27301
rect 11685 27196 11726 27242
rect 11772 27196 11813 27242
rect 11685 27137 11813 27196
rect 11685 27135 11726 27137
rect 11772 27135 11813 27137
rect 11685 27083 11723 27135
rect 11775 27083 11813 27135
rect 11685 27032 11813 27083
rect 11685 26986 11726 27032
rect 11772 26986 11813 27032
rect 11685 26927 11813 26986
rect 11685 26917 11726 26927
rect 11772 26917 11813 26927
rect 11685 26865 11723 26917
rect 11775 26865 11813 26917
rect 11685 26825 11813 26865
rect 11950 27347 11996 27396
rect 12174 27392 12220 27406
rect 12363 27452 12479 27546
rect 12363 27406 12398 27452
rect 12444 27406 12479 27452
rect 12363 27396 12479 27406
rect 12622 27452 12668 27465
rect 13276 27418 13392 27432
rect 11950 27242 11996 27301
rect 11950 27137 11996 27196
rect 11950 27032 11996 27091
rect 11950 26927 11996 26986
rect 11502 26717 11548 26776
rect 11502 26612 11548 26671
rect 11502 26507 11548 26566
rect 11502 26402 11548 26461
rect 11502 26297 11548 26356
rect 11502 26192 11548 26251
rect 11502 26088 11548 26146
rect 11502 25984 11548 26042
rect 11502 25880 11548 25938
rect 11502 25776 11548 25834
rect 11502 25672 11548 25730
rect 11502 25568 11548 25626
rect 11502 25464 11548 25522
rect 11502 25360 11548 25418
rect 11502 25256 11548 25314
rect 11502 25197 11548 25210
rect 11726 26822 11772 26825
rect 11726 26717 11772 26776
rect 11726 26612 11772 26671
rect 11726 26507 11772 26566
rect 11726 26402 11772 26461
rect 11726 26297 11772 26356
rect 11726 26192 11772 26251
rect 11726 26088 11772 26146
rect 11726 25984 11772 26042
rect 11726 25880 11772 25938
rect 11726 25776 11772 25834
rect 11726 25672 11772 25730
rect 11726 25568 11772 25626
rect 11726 25464 11772 25522
rect 11726 25360 11772 25418
rect 11726 25256 11772 25314
rect 11726 25197 11772 25210
rect 11950 26822 11996 26881
rect 12133 27353 12261 27392
rect 12133 27301 12171 27353
rect 12223 27301 12261 27353
rect 12133 27242 12261 27301
rect 12133 27196 12174 27242
rect 12220 27196 12261 27242
rect 12133 27137 12261 27196
rect 12133 27135 12174 27137
rect 12220 27135 12261 27137
rect 12133 27083 12171 27135
rect 12223 27083 12261 27135
rect 12133 27032 12261 27083
rect 12133 26986 12174 27032
rect 12220 26986 12261 27032
rect 12133 26927 12261 26986
rect 12133 26917 12174 26927
rect 12220 26917 12261 26927
rect 12133 26865 12171 26917
rect 12223 26865 12261 26917
rect 12133 26825 12261 26865
rect 12398 27347 12444 27396
rect 12622 27392 12668 27406
rect 12398 27242 12444 27301
rect 12398 27137 12444 27196
rect 12398 27032 12444 27091
rect 12398 26927 12444 26986
rect 11950 26717 11996 26776
rect 11950 26612 11996 26671
rect 11950 26507 11996 26566
rect 11950 26402 11996 26461
rect 11950 26297 11996 26356
rect 11950 26192 11996 26251
rect 11950 26088 11996 26146
rect 11950 25984 11996 26042
rect 11950 25880 11996 25938
rect 11950 25776 11996 25834
rect 11950 25672 11996 25730
rect 11950 25568 11996 25626
rect 11950 25464 11996 25522
rect 11950 25360 11996 25418
rect 11950 25256 11996 25314
rect 11950 25197 11996 25210
rect 12174 26822 12220 26825
rect 12174 26717 12220 26776
rect 12174 26612 12220 26671
rect 12174 26507 12220 26566
rect 12174 26402 12220 26461
rect 12174 26297 12220 26356
rect 12174 26192 12220 26251
rect 12174 26088 12220 26146
rect 12174 25984 12220 26042
rect 12174 25880 12220 25938
rect 12174 25776 12220 25834
rect 12174 25672 12220 25730
rect 12174 25568 12220 25626
rect 12174 25464 12220 25522
rect 12174 25360 12220 25418
rect 12174 25256 12220 25314
rect 12174 25197 12220 25210
rect 12398 26822 12444 26881
rect 12581 27353 12709 27392
rect 12581 27301 12619 27353
rect 12671 27301 12709 27353
rect 12581 27242 12709 27301
rect 12581 27196 12622 27242
rect 12668 27196 12709 27242
rect 12581 27137 12709 27196
rect 12581 27135 12622 27137
rect 12668 27135 12709 27137
rect 12581 27083 12619 27135
rect 12671 27083 12709 27135
rect 12581 27032 12709 27083
rect 12990 27378 13114 27418
rect 12990 27326 13026 27378
rect 13078 27326 13114 27378
rect 12990 27160 13028 27326
rect 13074 27160 13114 27326
rect 12990 27108 13026 27160
rect 13078 27108 13114 27160
rect 12990 27068 13114 27108
rect 13266 27382 13392 27418
rect 13266 27378 13312 27382
rect 13266 27326 13302 27378
rect 13358 27336 13392 27382
rect 13354 27326 13392 27336
rect 13266 27178 13392 27326
rect 13266 27160 13312 27178
rect 13266 27108 13302 27160
rect 13358 27132 13392 27178
rect 13354 27108 13392 27132
rect 13266 27095 13392 27108
rect 13724 27382 13840 27614
rect 14150 27574 14312 27619
rect 14150 27528 14161 27574
rect 14301 27528 14312 27574
rect 14906 27643 16157 27695
rect 16209 27643 16247 27695
rect 14906 27568 16247 27643
rect 16704 27656 16750 27715
rect 16880 28076 17009 28122
rect 17152 28080 17198 28089
rect 16880 28030 16928 28076
rect 16974 28030 17009 28076
rect 16880 27975 17009 28030
rect 17113 28076 17241 28080
rect 17113 28041 17152 28076
rect 17198 28041 17241 28076
rect 17113 27989 17151 28041
rect 17203 27989 17241 28041
rect 16880 27971 17008 27975
rect 16880 27956 16928 27971
rect 16880 27904 16918 27956
rect 16974 27925 17008 27971
rect 16970 27904 17008 27925
rect 16880 27866 17008 27904
rect 16880 27820 16928 27866
rect 16974 27820 17008 27866
rect 16880 27761 17008 27820
rect 16880 27738 16928 27761
rect 16880 27686 16918 27738
rect 16974 27715 17008 27761
rect 16970 27686 17008 27715
rect 16880 27656 17008 27686
rect 16880 27646 16928 27656
rect 14150 27517 14312 27528
rect 13724 27336 13760 27382
rect 13806 27336 13840 27382
rect 13724 27178 13840 27336
rect 13724 27132 13760 27178
rect 13806 27132 13840 27178
rect 13266 27068 13390 27095
rect 12581 26986 12622 27032
rect 12668 26986 12709 27032
rect 12581 26927 12709 26986
rect 12581 26917 12622 26927
rect 12668 26917 12709 26927
rect 12581 26865 12619 26917
rect 12671 26865 12709 26917
rect 13724 27015 13840 27132
rect 14172 27382 14834 27432
rect 14172 27336 14208 27382
rect 14254 27336 14834 27382
rect 14172 27315 14834 27336
rect 14172 27269 14788 27315
rect 14172 27210 14834 27269
rect 14172 27178 14386 27210
rect 14172 27132 14208 27178
rect 14254 27158 14386 27178
rect 14438 27158 14598 27210
rect 14650 27159 14834 27210
rect 14650 27158 14788 27159
rect 14254 27132 14788 27158
rect 14172 27113 14788 27132
rect 14172 27100 14834 27113
rect 15012 27315 15058 27568
rect 16121 27477 16245 27568
rect 15012 27159 15058 27269
rect 15012 27100 15058 27113
rect 15236 27392 15606 27432
rect 15236 27340 15515 27392
rect 15567 27340 15606 27392
rect 16121 27425 16157 27477
rect 16209 27425 16245 27477
rect 16121 27385 16245 27425
rect 16704 27552 16750 27610
rect 16704 27448 16750 27506
rect 15236 27315 15520 27340
rect 15282 27269 15520 27315
rect 15236 27174 15520 27269
rect 15566 27174 15606 27340
rect 16704 27344 16750 27402
rect 16704 27265 16750 27298
rect 16974 27646 17008 27656
rect 17113 27971 17241 27989
rect 17341 28076 17457 28170
rect 17789 28122 17828 28170
rect 17880 28170 18552 28174
rect 17880 28122 17918 28170
rect 17600 28080 17646 28089
rect 17341 28030 17376 28076
rect 17422 28030 17457 28076
rect 17341 27975 17457 28030
rect 17557 28076 17685 28080
rect 17557 28041 17600 28076
rect 17646 28041 17685 28076
rect 17557 27989 17595 28041
rect 17647 27989 17685 28041
rect 17113 27925 17152 27971
rect 17198 27925 17241 27971
rect 17113 27866 17241 27925
rect 17113 27823 17152 27866
rect 17198 27823 17241 27866
rect 17113 27771 17151 27823
rect 17203 27771 17241 27823
rect 17113 27761 17241 27771
rect 17113 27715 17152 27761
rect 17198 27715 17241 27761
rect 17113 27656 17241 27715
rect 16928 27552 16974 27610
rect 17113 27610 17152 27656
rect 17198 27610 17241 27656
rect 17113 27605 17241 27610
rect 17113 27553 17151 27605
rect 17203 27553 17241 27605
rect 17113 27552 17241 27553
rect 17113 27513 17152 27552
rect 16928 27448 16974 27506
rect 16928 27344 16974 27402
rect 15236 27159 15515 27174
rect 15282 27122 15515 27159
rect 15567 27122 15606 27174
rect 15282 27113 15606 27122
rect 15236 27108 15606 27113
rect 16670 27240 16785 27265
rect 16670 27194 16704 27240
rect 16750 27194 16785 27240
rect 15236 27100 15282 27108
rect 14172 27095 14288 27100
rect 15479 27082 15603 27108
rect 16670 27105 16785 27194
rect 16928 27240 16974 27298
rect 17198 27513 17241 27552
rect 17376 27971 17422 27975
rect 17376 27866 17422 27925
rect 17376 27761 17422 27820
rect 17376 27656 17422 27715
rect 17376 27552 17422 27610
rect 17152 27448 17198 27506
rect 17152 27344 17198 27402
rect 17152 27265 17198 27298
rect 17557 27971 17685 27989
rect 17789 28076 17918 28122
rect 18514 28122 18552 28170
rect 18604 28170 19462 28174
rect 18604 28122 18643 28170
rect 17789 28030 17824 28076
rect 17870 28030 17918 28076
rect 17789 27975 17918 28030
rect 17557 27925 17600 27971
rect 17646 27925 17685 27971
rect 17557 27866 17685 27925
rect 17557 27823 17600 27866
rect 17646 27823 17685 27866
rect 17557 27771 17595 27823
rect 17647 27771 17685 27823
rect 17557 27761 17685 27771
rect 17557 27715 17600 27761
rect 17646 27715 17685 27761
rect 17557 27656 17685 27715
rect 17557 27610 17600 27656
rect 17646 27610 17685 27656
rect 17790 27971 17918 27975
rect 17790 27925 17824 27971
rect 17870 27956 17918 27971
rect 17790 27904 17828 27925
rect 17880 27904 17918 27956
rect 17790 27866 17918 27904
rect 17790 27820 17824 27866
rect 17870 27820 17918 27866
rect 17790 27761 17918 27820
rect 17790 27715 17824 27761
rect 17870 27738 17918 27761
rect 17790 27686 17828 27715
rect 17880 27686 17918 27738
rect 17790 27656 17918 27686
rect 17790 27646 17824 27656
rect 17557 27605 17685 27610
rect 17557 27553 17595 27605
rect 17647 27553 17685 27605
rect 17557 27552 17685 27553
rect 17557 27513 17600 27552
rect 17376 27448 17422 27506
rect 17376 27344 17422 27402
rect 16928 27181 16974 27194
rect 17118 27240 17233 27265
rect 17118 27194 17152 27240
rect 17198 27194 17233 27240
rect 17118 27105 17233 27194
rect 17376 27240 17422 27298
rect 17646 27513 17685 27552
rect 17870 27646 17918 27656
rect 18048 28076 18094 28089
rect 18048 27971 18094 28030
rect 18048 27866 18094 27925
rect 18048 27761 18094 27820
rect 18048 27656 18094 27715
rect 17824 27552 17870 27610
rect 17600 27448 17646 27506
rect 17600 27344 17646 27402
rect 17600 27265 17646 27298
rect 17824 27448 17870 27506
rect 17824 27344 17870 27402
rect 17376 27181 17422 27194
rect 17565 27240 17680 27265
rect 17565 27194 17600 27240
rect 17646 27194 17680 27240
rect 14918 27021 15174 27032
rect 14918 27015 14929 27021
rect 13724 26975 14929 27015
rect 15163 26975 15174 27021
rect 13724 26974 15174 26975
rect 13724 26922 14384 26974
rect 14436 26922 14596 26974
rect 14648 26922 15174 26974
rect 13724 26895 15174 26922
rect 16670 26986 17233 27105
rect 14346 26882 14686 26895
rect 16670 26888 16785 26986
rect 17117 26985 17233 26986
rect 12581 26825 12709 26865
rect 16670 26842 16704 26888
rect 16750 26842 16785 26888
rect 16670 26841 16785 26842
rect 16928 26888 16974 26901
rect 12398 26717 12444 26776
rect 12398 26612 12444 26671
rect 12398 26507 12444 26566
rect 12398 26402 12444 26461
rect 12398 26297 12444 26356
rect 12398 26192 12444 26251
rect 12398 26088 12444 26146
rect 12398 25984 12444 26042
rect 12398 25880 12444 25938
rect 12398 25776 12444 25834
rect 12398 25672 12444 25730
rect 12398 25568 12444 25626
rect 12398 25464 12444 25522
rect 12398 25360 12444 25418
rect 12398 25256 12444 25314
rect 12398 25197 12444 25210
rect 12622 26822 12668 26825
rect 12622 26717 12668 26776
rect 16704 26783 16750 26841
rect 12622 26612 12668 26671
rect 13470 26731 13516 26744
rect 12622 26507 12668 26566
rect 12622 26402 12668 26461
rect 12622 26297 12668 26356
rect 12622 26192 12668 26251
rect 12622 26088 12668 26146
rect 12622 25984 12668 26042
rect 12622 25880 12668 25938
rect 12622 25776 12668 25834
rect 12622 25672 12668 25730
rect 12622 25568 12668 25626
rect 12622 25464 12668 25522
rect 12622 25360 12668 25418
rect 13118 26545 13470 26643
rect 13118 26499 13166 26545
rect 13212 26514 13470 26545
rect 13694 26731 13740 26744
rect 13212 26499 13253 26514
rect 13118 26462 13253 26499
rect 13305 26462 13460 26514
rect 13118 26382 13470 26462
rect 13118 26336 13166 26382
rect 13212 26379 13470 26382
rect 13516 26379 13550 26643
rect 13212 26336 13550 26379
rect 13118 26322 13550 26336
rect 13118 26296 13470 26322
rect 13118 26244 13253 26296
rect 13305 26244 13460 26296
rect 13516 26276 13550 26322
rect 13512 26244 13550 26276
rect 13118 26219 13550 26244
rect 13118 26218 13470 26219
rect 13118 26172 13166 26218
rect 13212 26173 13470 26218
rect 13516 26173 13550 26219
rect 13212 26172 13550 26173
rect 13118 26116 13550 26172
rect 13118 26078 13470 26116
rect 13118 26055 13253 26078
rect 13118 26009 13166 26055
rect 13212 26026 13253 26055
rect 13305 26026 13460 26078
rect 13516 26070 13550 26116
rect 13512 26026 13550 26070
rect 13212 26013 13550 26026
rect 13212 26009 13470 26013
rect 13118 25967 13470 26009
rect 13516 25967 13550 26013
rect 13118 25910 13550 25967
rect 13118 25892 13470 25910
rect 13118 25846 13166 25892
rect 13212 25864 13470 25892
rect 13516 25864 13550 25910
rect 13212 25860 13550 25864
rect 13212 25846 13253 25860
rect 13118 25808 13253 25846
rect 13305 25808 13460 25860
rect 13512 25808 13550 25860
rect 13118 25807 13550 25808
rect 13118 25761 13470 25807
rect 13516 25761 13550 25807
rect 13118 25728 13550 25761
rect 13118 25682 13166 25728
rect 13212 25704 13550 25728
rect 13212 25682 13470 25704
rect 13118 25658 13470 25682
rect 13516 25658 13550 25704
rect 13118 25601 13550 25658
rect 13118 25565 13470 25601
rect 13118 25519 13166 25565
rect 13212 25555 13470 25565
rect 13516 25555 13550 25601
rect 13212 25519 13550 25555
rect 13118 25498 13550 25519
rect 13118 25452 13470 25498
rect 13516 25452 13550 25498
rect 13118 25395 13550 25452
rect 15161 26731 15207 26744
rect 14809 26545 15161 26643
rect 13694 26322 13740 26379
rect 13694 26219 13740 26276
rect 13694 26116 13740 26173
rect 13694 26013 13740 26070
rect 13694 25910 13740 25967
rect 13694 25807 13740 25864
rect 13694 25704 13740 25761
rect 13942 26491 14070 26531
rect 13942 26439 13980 26491
rect 14032 26439 14070 26491
rect 14809 26499 14857 26545
rect 14903 26514 15161 26545
rect 15385 26731 15431 26744
rect 14903 26499 14944 26514
rect 14809 26462 14944 26499
rect 14996 26462 15151 26514
rect 13942 26400 13984 26439
rect 14030 26400 14070 26439
rect 13942 26338 14070 26400
rect 13942 26292 13984 26338
rect 14030 26292 14070 26338
rect 13942 26273 14070 26292
rect 13942 26221 13980 26273
rect 14032 26221 14070 26273
rect 13942 26184 13984 26221
rect 14030 26184 14070 26221
rect 13942 26122 14070 26184
rect 13942 26076 13984 26122
rect 14030 26076 14070 26122
rect 13942 26055 14070 26076
rect 13942 26003 13980 26055
rect 14032 26003 14070 26055
rect 13942 25968 13984 26003
rect 14030 25968 14070 26003
rect 13942 25906 14070 25968
rect 13942 25860 13984 25906
rect 14030 25860 14070 25906
rect 13942 25837 14070 25860
rect 13942 25785 13980 25837
rect 14032 25785 14070 25837
rect 13942 25752 13984 25785
rect 14030 25752 14070 25785
rect 13942 25745 14070 25752
rect 14208 26446 14254 26459
rect 14208 26338 14254 26400
rect 14208 26230 14254 26292
rect 14208 26122 14254 26184
rect 14208 26014 14254 26076
rect 14208 25906 14254 25968
rect 14208 25798 14254 25860
rect 13694 25601 13740 25658
rect 13694 25498 13740 25555
rect 13694 25405 13740 25452
rect 13984 25690 14030 25745
rect 13984 25582 14030 25644
rect 13984 25474 14030 25536
rect 13984 25415 14030 25428
rect 14208 25690 14254 25752
rect 14208 25582 14254 25644
rect 14208 25474 14254 25536
rect 13118 25349 13470 25395
rect 13516 25349 13550 25395
rect 13118 25344 13550 25349
rect 13659 25395 13774 25405
rect 13659 25349 13694 25395
rect 13740 25349 13774 25395
rect 13470 25336 13516 25344
rect 12622 25256 12668 25314
rect 12622 25197 12668 25210
rect 13215 25255 13555 25262
rect 13659 25255 13774 25349
rect 13215 25221 13572 25255
rect 13215 25169 13253 25221
rect 13305 25218 13465 25221
rect 13517 25218 13572 25221
rect 13305 25172 13333 25218
rect 13379 25172 13465 25218
rect 13537 25172 13572 25218
rect 13305 25169 13465 25172
rect 13517 25169 13572 25172
rect 13215 25135 13572 25169
rect 13659 25218 14082 25255
rect 13659 25172 13843 25218
rect 13889 25172 14001 25218
rect 14047 25172 14082 25218
rect 13659 25135 14082 25172
rect 13215 25129 13555 25135
rect 9115 25088 9903 25126
rect 9115 25042 9274 25088
rect 9696 25042 9903 25088
rect 9115 25007 9903 25042
rect 10011 25088 10799 25126
rect 10011 25042 10218 25088
rect 10640 25042 10799 25088
rect 10011 25007 10799 25042
rect 10907 25088 11695 25126
rect 10907 25042 11066 25088
rect 11488 25042 11695 25088
rect 10907 25007 11695 25042
rect 11803 25088 12591 25126
rect 11803 25042 12010 25088
rect 12432 25042 12591 25088
rect 11803 25007 12591 25042
rect 8342 24811 8389 24851
rect 8351 24759 8389 24811
rect 8342 24593 8389 24759
rect 8351 24541 8389 24593
rect 8342 24376 8389 24541
rect 8351 24324 8389 24376
rect 8342 24158 8389 24324
rect 8351 24106 8389 24158
rect 8342 23940 8389 24106
rect 8351 23888 8389 23940
rect 8342 23722 8389 23888
rect 8351 23670 8389 23722
rect 8342 23505 8389 23670
rect 8351 23453 8389 23505
rect 8342 23427 8389 23453
rect 8262 23370 8389 23427
rect 8262 23324 8296 23370
rect 8342 23324 8389 23370
rect 8262 23287 8389 23324
rect 8262 23267 8299 23287
rect 8262 23221 8296 23267
rect 8351 23235 8389 23287
rect 8342 23221 8389 23235
rect 8262 23195 8389 23221
rect 9385 25006 9502 25007
rect 10412 25006 10529 25007
rect 8863 24854 9277 24890
rect 8863 24808 9038 24854
rect 9084 24808 9197 24854
rect 9243 24813 9277 24854
rect 9243 24808 9286 24813
rect 8863 24773 9286 24808
rect 8863 24771 9196 24773
rect 8520 23370 8566 23427
rect 8520 23267 8566 23324
rect 8296 23164 8342 23195
rect 8296 23061 8342 23118
rect 8296 22958 8342 23015
rect 8296 22855 8342 22912
rect 8296 22752 8342 22809
rect 8520 23164 8566 23221
rect 8520 23061 8566 23118
rect 8520 22958 8566 23015
rect 8520 22855 8566 22912
rect 8520 22752 8566 22809
rect 8296 22649 8342 22706
rect 8296 22546 8342 22603
rect 8296 22443 8342 22500
rect 8296 22384 8342 22397
rect 8480 22706 8520 22743
rect 9158 24721 9196 24771
rect 9248 24721 9286 24773
rect 9158 24556 9286 24721
rect 8566 22706 8604 22743
rect 9158 22722 9196 24556
rect 9248 24504 9286 24556
rect 9242 24338 9286 24504
rect 9385 24550 9501 25006
rect 9385 24456 9420 24550
rect 9248 24286 9286 24338
rect 9242 24121 9286 24286
rect 9248 24069 9286 24121
rect 9242 23903 9286 24069
rect 9248 23851 9286 23903
rect 9242 23685 9286 23851
rect 9248 23633 9286 23685
rect 9242 23467 9286 23633
rect 9248 23415 9286 23467
rect 9242 23250 9286 23415
rect 9248 23198 9286 23250
rect 9242 23032 9286 23198
rect 9248 22980 9286 23032
rect 9242 22815 9286 22980
rect 9248 22763 9286 22815
rect 8480 22703 8604 22706
rect 8480 22651 8516 22703
rect 8568 22651 8604 22703
rect 8480 22649 8604 22651
rect 8480 22603 8520 22649
rect 8566 22603 8604 22649
rect 8480 22546 8604 22603
rect 8480 22500 8520 22546
rect 8566 22500 8604 22546
rect 8480 22485 8604 22500
rect 8480 22433 8516 22485
rect 8568 22433 8604 22485
rect 8480 22397 8520 22433
rect 8566 22397 8604 22433
rect 8480 22393 8604 22397
rect 9242 22722 9286 22763
rect 9196 22509 9242 22566
rect 9196 22406 9242 22463
rect 8520 22384 8566 22393
rect 9196 22303 9242 22360
rect 9196 22200 9242 22257
rect 9196 22097 9242 22154
rect 9196 21994 9242 22051
rect 9196 21891 9242 21948
rect 9466 24456 9501 24550
rect 9609 24854 10305 24890
rect 9609 24808 9645 24854
rect 9691 24808 9803 24854
rect 9849 24808 10065 24854
rect 10111 24808 10223 24854
rect 10269 24808 10305 24854
rect 9609 24773 10305 24808
rect 9609 24721 9648 24773
rect 9700 24721 9931 24773
rect 9983 24721 10214 24773
rect 10266 24721 10305 24773
rect 9609 24556 10305 24721
rect 9609 24550 9648 24556
rect 9420 22509 9466 22566
rect 9420 22406 9466 22463
rect 9420 22303 9466 22360
rect 9420 22200 9466 22257
rect 9420 22097 9466 22154
rect 9420 21994 9466 22051
rect 9420 21891 9466 21948
rect 8052 21796 8090 21836
rect 7966 21744 8002 21796
rect 8054 21744 8090 21796
rect 7966 21578 8006 21744
rect 8052 21578 8090 21744
rect 7966 21526 8002 21578
rect 8054 21526 8090 21578
rect 7966 21490 8006 21526
rect 8052 21490 8090 21526
rect 9196 21788 9242 21845
rect 9196 21685 9242 21742
rect 9196 21582 9242 21639
rect 9196 21523 9242 21536
rect 9382 21845 9420 21882
rect 9609 22566 9644 24550
rect 9700 24504 9931 24556
rect 9983 24504 10214 24556
rect 10266 24550 10305 24556
rect 9690 24338 10224 24504
rect 9700 24286 9931 24338
rect 9983 24286 10214 24338
rect 9690 24121 10224 24286
rect 9700 24069 9931 24121
rect 9983 24069 10214 24121
rect 9690 23903 10224 24069
rect 9700 23851 9931 23903
rect 9983 23851 10214 23903
rect 9690 23685 10224 23851
rect 9700 23633 9931 23685
rect 9983 23633 10214 23685
rect 9690 23467 10224 23633
rect 9700 23415 9931 23467
rect 9983 23415 10214 23467
rect 9690 23250 10224 23415
rect 9700 23198 9931 23250
rect 9983 23198 10214 23250
rect 9690 23032 10224 23198
rect 9700 22980 9931 23032
rect 9983 22980 10214 23032
rect 9690 22815 10224 22980
rect 9700 22763 9931 22815
rect 9983 22763 10214 22815
rect 9690 22566 10224 22763
rect 10270 22566 10305 24550
rect 10413 24550 10529 25006
rect 11177 25006 11294 25007
rect 12204 25006 12321 25007
rect 13470 25006 13516 25015
rect 10637 24854 11069 24890
rect 10637 24813 10671 24854
rect 10413 24456 10448 24550
rect 9609 22509 10305 22566
rect 9609 22463 9644 22509
rect 9690 22463 10224 22509
rect 10270 22463 10305 22509
rect 9609 22406 10305 22463
rect 9609 22360 9644 22406
rect 9690 22360 10224 22406
rect 10270 22360 10305 22406
rect 9609 22303 10305 22360
rect 9609 22257 9644 22303
rect 9690 22257 10224 22303
rect 10270 22257 10305 22303
rect 9609 22200 10305 22257
rect 9609 22154 9644 22200
rect 9690 22154 10224 22200
rect 10270 22154 10305 22200
rect 9609 22097 10305 22154
rect 9609 22051 9644 22097
rect 9690 22051 10224 22097
rect 10270 22051 10305 22097
rect 9609 21994 10305 22051
rect 9609 21948 9644 21994
rect 9690 21989 10224 21994
rect 9690 21948 9934 21989
rect 9609 21891 9934 21948
rect 9466 21845 9506 21882
rect 9382 21842 9506 21845
rect 9382 21790 9418 21842
rect 9470 21790 9506 21842
rect 9382 21788 9506 21790
rect 9382 21742 9420 21788
rect 9466 21742 9506 21788
rect 9382 21685 9506 21742
rect 9382 21639 9420 21685
rect 9466 21639 9506 21685
rect 9382 21624 9506 21639
rect 9382 21572 9418 21624
rect 9470 21572 9506 21624
rect 9382 21536 9420 21572
rect 9466 21536 9506 21572
rect 9382 21532 9506 21536
rect 9609 21845 9644 21891
rect 9690 21845 9934 21891
rect 9609 21788 9934 21845
rect 9609 21742 9644 21788
rect 9690 21742 9934 21788
rect 9609 21685 9934 21742
rect 9609 21639 9644 21685
rect 9690 21661 9934 21685
rect 9980 21948 10224 21989
rect 10270 21948 10305 21994
rect 9980 21891 10305 21948
rect 9980 21845 10224 21891
rect 10270 21845 10305 21891
rect 10494 24456 10529 24550
rect 10628 24808 10671 24813
rect 10717 24808 10830 24854
rect 10876 24808 10989 24854
rect 11035 24813 11069 24854
rect 11035 24808 11078 24813
rect 10628 24773 11078 24808
rect 10628 24721 10666 24773
rect 10718 24771 10988 24773
rect 10718 24721 10756 24771
rect 10628 24556 10756 24721
rect 10628 24504 10666 24556
rect 10628 24338 10672 24504
rect 10628 24286 10666 24338
rect 10628 24121 10672 24286
rect 10628 24069 10666 24121
rect 10628 23903 10672 24069
rect 10628 23851 10666 23903
rect 10628 23685 10672 23851
rect 10628 23633 10666 23685
rect 10628 23467 10672 23633
rect 10628 23415 10666 23467
rect 10628 23250 10672 23415
rect 10628 23198 10666 23250
rect 10628 23032 10672 23198
rect 10628 22980 10666 23032
rect 10628 22815 10672 22980
rect 10628 22763 10666 22815
rect 10628 22722 10672 22763
rect 10448 22509 10494 22566
rect 10448 22406 10494 22463
rect 10448 22303 10494 22360
rect 10448 22200 10494 22257
rect 10448 22097 10494 22154
rect 10448 21994 10494 22051
rect 10448 21891 10494 21948
rect 9980 21788 10305 21845
rect 9980 21742 10224 21788
rect 10270 21742 10305 21788
rect 9980 21685 10305 21742
rect 9980 21661 10224 21685
rect 9690 21639 10224 21661
rect 10270 21639 10305 21685
rect 9609 21582 10305 21639
rect 9609 21536 9644 21582
rect 9690 21536 10224 21582
rect 10270 21536 10305 21582
rect 9420 21523 9466 21532
rect 9609 21531 10305 21536
rect 10408 21845 10448 21882
rect 10718 22722 10756 24556
rect 10950 24721 10988 24771
rect 11040 24721 11078 24773
rect 10950 24556 11078 24721
rect 10950 22722 10988 24556
rect 11040 24504 11078 24556
rect 11034 24338 11078 24504
rect 11177 24550 11293 25006
rect 11177 24456 11212 24550
rect 11040 24286 11078 24338
rect 11034 24121 11078 24286
rect 11040 24069 11078 24121
rect 11034 23903 11078 24069
rect 11040 23851 11078 23903
rect 11034 23685 11078 23851
rect 11040 23633 11078 23685
rect 11034 23467 11078 23633
rect 11040 23415 11078 23467
rect 11034 23250 11078 23415
rect 11040 23198 11078 23250
rect 11034 23032 11078 23198
rect 11040 22980 11078 23032
rect 11034 22815 11078 22980
rect 11040 22763 11078 22815
rect 10672 22509 10718 22566
rect 10672 22406 10718 22463
rect 10672 22303 10718 22360
rect 10672 22200 10718 22257
rect 10672 22097 10718 22154
rect 10672 21994 10718 22051
rect 10672 21891 10718 21948
rect 10494 21845 10532 21882
rect 10408 21842 10532 21845
rect 10408 21790 10444 21842
rect 10496 21790 10532 21842
rect 10408 21788 10532 21790
rect 10408 21742 10448 21788
rect 10494 21742 10532 21788
rect 10408 21685 10532 21742
rect 10408 21639 10448 21685
rect 10494 21639 10532 21685
rect 10408 21624 10532 21639
rect 10408 21572 10444 21624
rect 10496 21572 10532 21624
rect 10408 21536 10448 21572
rect 10494 21536 10532 21572
rect 10408 21532 10532 21536
rect 10672 21788 10718 21845
rect 10672 21685 10718 21742
rect 10672 21582 10718 21639
rect 9644 21523 9690 21531
rect 10224 21523 10270 21531
rect 10448 21523 10494 21532
rect 10672 21523 10718 21536
rect 11034 22722 11078 22763
rect 10988 22509 11034 22566
rect 10988 22406 11034 22463
rect 10988 22303 11034 22360
rect 10988 22200 11034 22257
rect 10988 22097 11034 22154
rect 10988 21994 11034 22051
rect 10988 21891 11034 21948
rect 11258 24456 11293 24550
rect 11401 24854 12097 24890
rect 11401 24808 11437 24854
rect 11483 24808 11595 24854
rect 11641 24808 11857 24854
rect 11903 24808 12015 24854
rect 12061 24808 12097 24854
rect 11401 24773 12097 24808
rect 11401 24721 11440 24773
rect 11492 24721 11723 24773
rect 11775 24721 12006 24773
rect 12058 24721 12097 24773
rect 11401 24556 12097 24721
rect 11401 24550 11440 24556
rect 11212 22509 11258 22566
rect 11212 22406 11258 22463
rect 11212 22303 11258 22360
rect 11212 22200 11258 22257
rect 11212 22097 11258 22154
rect 11212 21994 11258 22051
rect 11212 21891 11258 21948
rect 10988 21788 11034 21845
rect 10988 21685 11034 21742
rect 10988 21582 11034 21639
rect 10988 21523 11034 21536
rect 11174 21845 11212 21882
rect 11401 22566 11436 24550
rect 11492 24504 11723 24556
rect 11775 24504 12006 24556
rect 12058 24550 12097 24556
rect 11482 24338 12016 24504
rect 11492 24286 11723 24338
rect 11775 24286 12006 24338
rect 11482 24121 12016 24286
rect 11492 24069 11723 24121
rect 11775 24069 12006 24121
rect 11482 23903 12016 24069
rect 11492 23851 11723 23903
rect 11775 23851 12006 23903
rect 11482 23685 12016 23851
rect 11492 23633 11723 23685
rect 11775 23633 12006 23685
rect 11482 23467 12016 23633
rect 11492 23415 11723 23467
rect 11775 23415 12006 23467
rect 11482 23250 12016 23415
rect 11492 23198 11723 23250
rect 11775 23198 12006 23250
rect 11482 23032 12016 23198
rect 11492 22980 11723 23032
rect 11775 22980 12006 23032
rect 11482 22815 12016 22980
rect 11492 22763 11723 22815
rect 11775 22763 12006 22815
rect 11482 22566 12016 22763
rect 12062 22566 12097 24550
rect 12205 24550 12321 25006
rect 13070 25002 13550 25006
rect 13070 24890 13470 25002
rect 12429 24854 13470 24890
rect 12429 24813 12463 24854
rect 12205 24456 12240 24550
rect 11401 22509 12097 22566
rect 11401 22463 11436 22509
rect 11482 22463 12016 22509
rect 12062 22463 12097 22509
rect 11401 22406 12097 22463
rect 11401 22360 11436 22406
rect 11482 22360 12016 22406
rect 12062 22360 12097 22406
rect 11401 22303 12097 22360
rect 11401 22257 11436 22303
rect 11482 22257 12016 22303
rect 12062 22257 12097 22303
rect 11401 22200 12097 22257
rect 11401 22154 11436 22200
rect 11482 22154 12016 22200
rect 12062 22154 12097 22200
rect 11401 22097 12097 22154
rect 11401 22051 11436 22097
rect 11482 22051 12016 22097
rect 12062 22051 12097 22097
rect 11401 21994 12097 22051
rect 11401 21948 11436 21994
rect 11482 21989 12016 21994
rect 11482 21948 11726 21989
rect 11401 21891 11726 21948
rect 11258 21845 11298 21882
rect 11174 21842 11298 21845
rect 11174 21790 11210 21842
rect 11262 21790 11298 21842
rect 11174 21788 11298 21790
rect 11174 21742 11212 21788
rect 11258 21742 11298 21788
rect 11174 21685 11298 21742
rect 11174 21639 11212 21685
rect 11258 21639 11298 21685
rect 11174 21624 11298 21639
rect 11174 21572 11210 21624
rect 11262 21572 11298 21624
rect 11174 21536 11212 21572
rect 11258 21536 11298 21572
rect 11174 21532 11298 21536
rect 11401 21845 11436 21891
rect 11482 21845 11726 21891
rect 11401 21788 11726 21845
rect 11401 21742 11436 21788
rect 11482 21742 11726 21788
rect 11401 21685 11726 21742
rect 11401 21639 11436 21685
rect 11482 21661 11726 21685
rect 11772 21948 12016 21989
rect 12062 21948 12097 21994
rect 11772 21891 12097 21948
rect 11772 21845 12016 21891
rect 12062 21845 12097 21891
rect 12286 24456 12321 24550
rect 12420 24808 12463 24813
rect 12509 24808 12622 24854
rect 12668 24808 13105 24854
rect 13151 24808 13470 24854
rect 12420 24773 13470 24808
rect 13516 24843 13550 25002
rect 13659 25002 13774 25135
rect 13516 24842 13554 24843
rect 13516 24802 13563 24842
rect 12420 24721 12458 24773
rect 12510 24771 13470 24773
rect 12510 24721 12548 24771
rect 12420 24556 12548 24721
rect 12420 24504 12458 24556
rect 12420 24338 12464 24504
rect 12420 24286 12458 24338
rect 12420 24121 12464 24286
rect 12420 24069 12458 24121
rect 12420 23903 12464 24069
rect 12420 23851 12458 23903
rect 12420 23685 12464 23851
rect 12420 23633 12458 23685
rect 12420 23467 12464 23633
rect 12420 23415 12458 23467
rect 12420 23250 12464 23415
rect 12420 23198 12458 23250
rect 12420 23032 12464 23198
rect 12420 22980 12458 23032
rect 12420 22815 12464 22980
rect 12420 22763 12458 22815
rect 12420 22722 12464 22763
rect 12240 22509 12286 22566
rect 12240 22406 12286 22463
rect 12240 22303 12286 22360
rect 12240 22200 12286 22257
rect 12240 22097 12286 22154
rect 12240 21994 12286 22051
rect 12240 21891 12286 21948
rect 11772 21788 12097 21845
rect 11772 21742 12016 21788
rect 12062 21742 12097 21788
rect 11772 21685 12097 21742
rect 11772 21661 12016 21685
rect 11482 21639 12016 21661
rect 12062 21639 12097 21685
rect 11401 21582 12097 21639
rect 11401 21536 11436 21582
rect 11482 21536 12016 21582
rect 12062 21536 12097 21582
rect 11212 21523 11258 21532
rect 11401 21531 12097 21536
rect 12200 21845 12240 21882
rect 12510 22722 12548 24556
rect 13070 24690 13470 24771
rect 13525 24750 13563 24802
rect 13070 24644 13105 24690
rect 13151 24644 13470 24690
rect 13070 24527 13470 24644
rect 13516 24585 13563 24750
rect 13659 24668 13694 25002
rect 13525 24533 13563 24585
rect 13070 24481 13105 24527
rect 13151 24481 13470 24527
rect 13070 24364 13470 24481
rect 13516 24367 13563 24533
rect 13070 24318 13105 24364
rect 13151 24318 13470 24364
rect 13070 24201 13470 24318
rect 13525 24315 13563 24367
rect 13070 24155 13105 24201
rect 13151 24155 13470 24201
rect 13070 24037 13470 24155
rect 13516 24150 13563 24315
rect 13525 24098 13563 24150
rect 13070 23991 13105 24037
rect 13151 23991 13470 24037
rect 13070 23874 13470 23991
rect 13516 23932 13563 24098
rect 13525 23880 13563 23932
rect 13070 23828 13105 23874
rect 13151 23828 13470 23874
rect 13070 23711 13470 23828
rect 13516 23714 13563 23880
rect 13070 23665 13105 23711
rect 13151 23665 13470 23711
rect 13070 23548 13470 23665
rect 13525 23662 13563 23714
rect 13070 23502 13105 23548
rect 13151 23502 13470 23548
rect 13070 23384 13470 23502
rect 13516 23496 13563 23662
rect 13525 23444 13563 23496
rect 13070 23338 13105 23384
rect 13151 23338 13470 23384
rect 13070 23221 13470 23338
rect 13516 23279 13563 23444
rect 13525 23227 13563 23279
rect 13070 23175 13105 23221
rect 13151 23175 13470 23221
rect 13070 23058 13470 23175
rect 13516 23061 13563 23227
rect 13070 23012 13105 23058
rect 13151 23012 13470 23058
rect 13070 22894 13470 23012
rect 13525 23009 13563 23061
rect 13070 22848 13105 22894
rect 13151 22848 13470 22894
rect 13070 22731 13470 22848
rect 13516 22844 13563 23009
rect 13525 22792 13563 22844
rect 12464 22509 12510 22566
rect 12464 22406 12510 22463
rect 12464 22303 12510 22360
rect 12464 22200 12510 22257
rect 12464 22097 12510 22154
rect 12464 21994 12510 22051
rect 12464 21891 12510 21948
rect 12286 21845 12324 21882
rect 12200 21842 12324 21845
rect 12200 21790 12236 21842
rect 12288 21790 12324 21842
rect 12200 21788 12324 21790
rect 12200 21742 12240 21788
rect 12286 21742 12324 21788
rect 12200 21685 12324 21742
rect 12200 21639 12240 21685
rect 12286 21639 12324 21685
rect 12200 21624 12324 21639
rect 12200 21572 12236 21624
rect 12288 21572 12324 21624
rect 12200 21536 12240 21572
rect 12286 21536 12324 21572
rect 12200 21532 12324 21536
rect 12464 21788 12510 21845
rect 12464 21685 12510 21742
rect 12464 21582 12510 21639
rect 11436 21523 11482 21531
rect 12016 21523 12062 21531
rect 12240 21523 12286 21532
rect 12464 21523 12510 21536
rect 13070 22685 13105 22731
rect 13151 22685 13470 22731
rect 13070 22568 13470 22685
rect 13070 22522 13105 22568
rect 13151 22522 13470 22568
rect 13070 22405 13470 22522
rect 13070 22359 13105 22405
rect 13151 22359 13470 22405
rect 13070 22241 13470 22359
rect 13070 22195 13105 22241
rect 13151 22195 13470 22241
rect 13070 22078 13470 22195
rect 13070 22032 13105 22078
rect 13151 22032 13470 22078
rect 13070 21915 13470 22032
rect 13070 21869 13105 21915
rect 13151 21869 13470 21915
rect 13070 21752 13470 21869
rect 13070 21706 13105 21752
rect 13151 21706 13470 21752
rect 13070 21588 13470 21706
rect 13070 21542 13105 21588
rect 13151 21542 13470 21588
rect 7966 21486 8090 21490
rect 13070 21490 13470 21542
rect 13516 22751 13563 22792
rect 13516 21490 13550 22751
rect 13070 21486 13550 21490
rect 13652 21796 13694 21837
rect 13740 24668 13774 25002
rect 13984 25003 14030 25016
rect 13950 23427 13984 24851
rect 14208 25003 14254 25428
rect 14809 26382 15161 26462
rect 14809 26336 14857 26382
rect 14903 26379 15161 26382
rect 15207 26379 15241 26643
rect 14903 26336 15241 26379
rect 14809 26322 15241 26336
rect 14809 26296 15161 26322
rect 14809 26244 14944 26296
rect 14996 26244 15151 26296
rect 15207 26276 15241 26322
rect 15203 26244 15241 26276
rect 14809 26219 15241 26244
rect 14809 26218 15161 26219
rect 14809 26172 14857 26218
rect 14903 26173 15161 26218
rect 15207 26173 15241 26219
rect 14903 26172 15241 26173
rect 14809 26116 15241 26172
rect 14809 26078 15161 26116
rect 14809 26055 14944 26078
rect 14809 26009 14857 26055
rect 14903 26026 14944 26055
rect 14996 26026 15151 26078
rect 15207 26070 15241 26116
rect 15203 26026 15241 26070
rect 14903 26013 15241 26026
rect 14903 26009 15161 26013
rect 14809 25967 15161 26009
rect 15207 25967 15241 26013
rect 14809 25910 15241 25967
rect 14809 25892 15161 25910
rect 14809 25846 14857 25892
rect 14903 25864 15161 25892
rect 15207 25864 15241 25910
rect 14903 25860 15241 25864
rect 14903 25846 14944 25860
rect 14809 25808 14944 25846
rect 14996 25808 15151 25860
rect 15203 25808 15241 25860
rect 14809 25807 15241 25808
rect 14809 25761 15161 25807
rect 15207 25761 15241 25807
rect 14809 25728 15241 25761
rect 14809 25682 14857 25728
rect 14903 25704 15241 25728
rect 14903 25682 15161 25704
rect 14809 25658 15161 25682
rect 15207 25658 15241 25704
rect 14809 25601 15241 25658
rect 14809 25565 15161 25601
rect 14809 25519 14857 25565
rect 14903 25555 15161 25565
rect 15207 25555 15241 25601
rect 14903 25519 15241 25555
rect 14809 25498 15241 25519
rect 14809 25452 15161 25498
rect 15207 25452 15241 25498
rect 14809 25395 15241 25452
rect 16704 26678 16750 26737
rect 16704 26573 16750 26632
rect 15385 26322 15431 26379
rect 15385 26219 15431 26276
rect 15385 26116 15431 26173
rect 15385 26013 15431 26070
rect 15385 25910 15431 25967
rect 15385 25807 15431 25864
rect 15385 25704 15431 25761
rect 15633 26491 15761 26531
rect 15633 26439 15671 26491
rect 15723 26439 15761 26491
rect 16704 26468 16750 26527
rect 15633 26400 15675 26439
rect 15721 26400 15761 26439
rect 15633 26338 15761 26400
rect 15633 26292 15675 26338
rect 15721 26292 15761 26338
rect 15633 26273 15761 26292
rect 15633 26221 15671 26273
rect 15723 26221 15761 26273
rect 15633 26184 15675 26221
rect 15721 26184 15761 26221
rect 15633 26122 15761 26184
rect 15633 26076 15675 26122
rect 15721 26076 15761 26122
rect 15633 26055 15761 26076
rect 15633 26003 15671 26055
rect 15723 26003 15761 26055
rect 15633 25968 15675 26003
rect 15721 25968 15761 26003
rect 15633 25906 15761 25968
rect 15633 25860 15675 25906
rect 15721 25860 15761 25906
rect 15633 25837 15761 25860
rect 15633 25785 15671 25837
rect 15723 25785 15761 25837
rect 15633 25752 15675 25785
rect 15721 25752 15761 25785
rect 15633 25745 15761 25752
rect 15899 26446 15945 26459
rect 15899 26338 15945 26400
rect 15899 26230 15945 26292
rect 15899 26122 15945 26184
rect 15899 26014 15945 26076
rect 15899 25906 15945 25968
rect 15899 25798 15945 25860
rect 15385 25601 15431 25658
rect 15385 25498 15431 25555
rect 15385 25405 15431 25452
rect 15675 25690 15721 25745
rect 15675 25582 15721 25644
rect 15675 25474 15721 25536
rect 15675 25415 15721 25428
rect 15899 25690 15945 25752
rect 15899 25582 15945 25644
rect 15899 25474 15945 25536
rect 14809 25349 15161 25395
rect 15207 25349 15241 25395
rect 14809 25344 15241 25349
rect 15350 25395 15465 25405
rect 15350 25349 15385 25395
rect 15431 25349 15465 25395
rect 15161 25336 15207 25344
rect 14906 25255 15246 25262
rect 15350 25255 15465 25349
rect 14906 25221 15263 25255
rect 14906 25169 14944 25221
rect 14996 25218 15156 25221
rect 15208 25218 15263 25221
rect 14996 25172 15024 25218
rect 15070 25172 15156 25218
rect 15228 25172 15263 25218
rect 14996 25169 15156 25172
rect 15208 25169 15263 25172
rect 14906 25135 15263 25169
rect 15350 25218 15773 25255
rect 15350 25172 15534 25218
rect 15580 25172 15692 25218
rect 15738 25172 15773 25218
rect 15350 25135 15773 25172
rect 14906 25129 15246 25135
rect 15161 25006 15207 25015
rect 14030 24811 14077 24851
rect 14039 24759 14077 24811
rect 14030 24593 14077 24759
rect 14039 24541 14077 24593
rect 14030 24376 14077 24541
rect 14039 24324 14077 24376
rect 14030 24158 14077 24324
rect 14039 24106 14077 24158
rect 14030 23940 14077 24106
rect 14039 23888 14077 23940
rect 14030 23722 14077 23888
rect 14039 23670 14077 23722
rect 14030 23505 14077 23670
rect 14039 23453 14077 23505
rect 14030 23427 14077 23453
rect 13950 23370 14077 23427
rect 13950 23324 13984 23370
rect 14030 23324 14077 23370
rect 13950 23287 14077 23324
rect 13950 23267 13987 23287
rect 13950 23221 13984 23267
rect 14039 23235 14077 23287
rect 14030 23221 14077 23235
rect 13950 23195 14077 23221
rect 14208 23370 14254 23427
rect 14208 23267 14254 23324
rect 13984 23164 14030 23195
rect 13984 23061 14030 23118
rect 13984 22958 14030 23015
rect 13984 22855 14030 22912
rect 13984 22752 14030 22809
rect 14208 23164 14254 23221
rect 14208 23061 14254 23118
rect 14208 22958 14254 23015
rect 14208 22855 14254 22912
rect 14208 22752 14254 22809
rect 13984 22649 14030 22706
rect 13984 22546 14030 22603
rect 13984 22443 14030 22500
rect 13984 22384 14030 22397
rect 14168 22706 14208 22743
rect 14761 25002 15241 25006
rect 14761 24854 15161 25002
rect 14761 24808 14796 24854
rect 14842 24808 15161 24854
rect 14761 24690 15161 24808
rect 15207 24843 15241 25002
rect 15350 25002 15465 25135
rect 15207 24842 15245 24843
rect 15207 24802 15254 24842
rect 15216 24750 15254 24802
rect 14761 24644 14796 24690
rect 14842 24644 15161 24690
rect 14761 24527 15161 24644
rect 15207 24585 15254 24750
rect 15350 24668 15385 25002
rect 15216 24533 15254 24585
rect 14761 24481 14796 24527
rect 14842 24481 15161 24527
rect 14761 24364 15161 24481
rect 15207 24367 15254 24533
rect 14761 24318 14796 24364
rect 14842 24318 15161 24364
rect 14761 24201 15161 24318
rect 15216 24315 15254 24367
rect 14761 24155 14796 24201
rect 14842 24155 15161 24201
rect 14761 24037 15161 24155
rect 15207 24150 15254 24315
rect 15216 24098 15254 24150
rect 14761 23991 14796 24037
rect 14842 23991 15161 24037
rect 14761 23874 15161 23991
rect 15207 23932 15254 24098
rect 15216 23880 15254 23932
rect 14761 23828 14796 23874
rect 14842 23828 15161 23874
rect 14761 23711 15161 23828
rect 15207 23714 15254 23880
rect 14761 23665 14796 23711
rect 14842 23665 15161 23711
rect 14761 23548 15161 23665
rect 15216 23662 15254 23714
rect 14761 23502 14796 23548
rect 14842 23502 15161 23548
rect 14761 23384 15161 23502
rect 15207 23496 15254 23662
rect 15216 23444 15254 23496
rect 14761 23338 14796 23384
rect 14842 23338 15161 23384
rect 14761 23221 15161 23338
rect 15207 23279 15254 23444
rect 15216 23227 15254 23279
rect 14761 23175 14796 23221
rect 14842 23175 15161 23221
rect 14761 23058 15161 23175
rect 15207 23061 15254 23227
rect 14761 23012 14796 23058
rect 14842 23012 15161 23058
rect 14761 22894 15161 23012
rect 15216 23009 15254 23061
rect 14761 22848 14796 22894
rect 14842 22848 15161 22894
rect 14254 22706 14292 22743
rect 14168 22703 14292 22706
rect 14168 22651 14204 22703
rect 14256 22651 14292 22703
rect 14168 22649 14292 22651
rect 14168 22603 14208 22649
rect 14254 22603 14292 22649
rect 14168 22546 14292 22603
rect 14168 22500 14208 22546
rect 14254 22500 14292 22546
rect 14168 22485 14292 22500
rect 14168 22433 14204 22485
rect 14256 22433 14292 22485
rect 14168 22397 14208 22433
rect 14254 22397 14292 22433
rect 14168 22393 14292 22397
rect 14761 22731 15161 22848
rect 15207 22844 15254 23009
rect 15216 22792 15254 22844
rect 14761 22685 14796 22731
rect 14842 22685 15161 22731
rect 14761 22568 15161 22685
rect 14761 22522 14796 22568
rect 14842 22522 15161 22568
rect 14761 22405 15161 22522
rect 14208 22384 14254 22393
rect 14761 22359 14796 22405
rect 14842 22359 15161 22405
rect 14761 22241 15161 22359
rect 14761 22195 14796 22241
rect 14842 22195 15161 22241
rect 14761 22078 15161 22195
rect 14761 22032 14796 22078
rect 14842 22032 15161 22078
rect 14761 21915 15161 22032
rect 14761 21869 14796 21915
rect 14842 21869 15161 21915
rect 13740 21796 13781 21837
rect 13652 21744 13690 21796
rect 13742 21744 13781 21796
rect 13652 21578 13694 21744
rect 13740 21578 13781 21744
rect 13652 21526 13690 21578
rect 13742 21526 13781 21578
rect 13652 21490 13694 21526
rect 13740 21490 13781 21526
rect 7782 21477 7828 21486
rect 8006 21477 8052 21486
rect 13470 21477 13516 21486
rect 9273 21383 9388 21399
rect 10525 21383 10640 21399
rect 13652 21383 13781 21490
rect 14761 21752 15161 21869
rect 14761 21706 14796 21752
rect 14842 21706 15161 21752
rect 14761 21588 15161 21706
rect 14761 21542 14796 21588
rect 14842 21542 15161 21588
rect 14761 21490 15161 21542
rect 15207 22751 15254 22792
rect 15207 21490 15241 22751
rect 14761 21486 15241 21490
rect 15345 21796 15385 21836
rect 15431 24668 15465 25002
rect 15675 25003 15721 25016
rect 15641 23427 15675 24851
rect 15899 25003 15945 25428
rect 15721 24811 15768 24851
rect 15730 24759 15768 24811
rect 15721 24593 15768 24759
rect 15730 24541 15768 24593
rect 15721 24376 15768 24541
rect 15730 24324 15768 24376
rect 15721 24158 15768 24324
rect 15730 24106 15768 24158
rect 15721 23940 15768 24106
rect 15730 23888 15768 23940
rect 15721 23722 15768 23888
rect 15730 23670 15768 23722
rect 15721 23505 15768 23670
rect 15730 23453 15768 23505
rect 15721 23427 15768 23453
rect 15641 23370 15768 23427
rect 15641 23324 15675 23370
rect 15721 23324 15768 23370
rect 15641 23287 15768 23324
rect 15641 23267 15678 23287
rect 15641 23221 15675 23267
rect 15730 23235 15768 23287
rect 15721 23221 15768 23235
rect 15641 23195 15768 23221
rect 16704 26363 16750 26422
rect 16704 26258 16750 26317
rect 16704 26153 16750 26212
rect 16704 26048 16750 26107
rect 16704 25943 16750 26002
rect 16704 25838 16750 25897
rect 16704 25733 16750 25792
rect 16704 25628 16750 25687
rect 16704 25524 16750 25582
rect 16704 25420 16750 25478
rect 16704 25316 16750 25374
rect 16928 26783 16974 26842
rect 17118 26888 17233 26985
rect 17565 27105 17680 27194
rect 17824 27240 17870 27298
rect 18048 27552 18094 27610
rect 18048 27448 18094 27506
rect 18048 27344 18094 27402
rect 18048 27265 18094 27298
rect 18338 28076 18384 28089
rect 18338 27971 18384 28030
rect 18338 27866 18384 27925
rect 18338 27761 18384 27820
rect 18338 27656 18384 27715
rect 18514 28076 18643 28122
rect 18786 28080 18832 28089
rect 18514 28030 18562 28076
rect 18608 28030 18643 28076
rect 18514 27975 18643 28030
rect 18747 28076 18875 28080
rect 18747 28041 18786 28076
rect 18832 28041 18875 28076
rect 18747 27989 18785 28041
rect 18837 27989 18875 28041
rect 18514 27971 18642 27975
rect 18514 27956 18562 27971
rect 18514 27904 18552 27956
rect 18608 27925 18642 27971
rect 18604 27904 18642 27925
rect 18514 27866 18642 27904
rect 18514 27820 18562 27866
rect 18608 27820 18642 27866
rect 18514 27761 18642 27820
rect 18514 27738 18562 27761
rect 18514 27686 18552 27738
rect 18608 27715 18642 27761
rect 18604 27686 18642 27715
rect 18514 27656 18642 27686
rect 18514 27646 18562 27656
rect 18338 27552 18384 27610
rect 18338 27448 18384 27506
rect 18338 27344 18384 27402
rect 18338 27265 18384 27298
rect 18608 27646 18642 27656
rect 18747 27971 18875 27989
rect 18975 28076 19091 28170
rect 19423 28122 19462 28170
rect 19514 28170 20185 28174
rect 19514 28122 19552 28170
rect 19234 28080 19280 28089
rect 18975 28030 19010 28076
rect 19056 28030 19091 28076
rect 18975 27975 19091 28030
rect 19191 28076 19319 28080
rect 19191 28041 19234 28076
rect 19280 28041 19319 28076
rect 19191 27989 19229 28041
rect 19281 27989 19319 28041
rect 18747 27925 18786 27971
rect 18832 27925 18875 27971
rect 18747 27866 18875 27925
rect 18747 27823 18786 27866
rect 18832 27823 18875 27866
rect 18747 27771 18785 27823
rect 18837 27771 18875 27823
rect 18747 27761 18875 27771
rect 18747 27715 18786 27761
rect 18832 27715 18875 27761
rect 18747 27656 18875 27715
rect 18562 27552 18608 27610
rect 18747 27610 18786 27656
rect 18832 27610 18875 27656
rect 18747 27605 18875 27610
rect 18747 27553 18785 27605
rect 18837 27553 18875 27605
rect 18747 27552 18875 27553
rect 18747 27513 18786 27552
rect 18562 27448 18608 27506
rect 18562 27344 18608 27402
rect 17824 27181 17870 27194
rect 18013 27240 18128 27265
rect 18013 27194 18048 27240
rect 18094 27194 18128 27240
rect 18013 27105 18128 27194
rect 17565 26986 18128 27105
rect 17565 26985 17681 26986
rect 17118 26842 17152 26888
rect 17198 26842 17233 26888
rect 17118 26841 17233 26842
rect 17376 26888 17422 26901
rect 16928 26678 16974 26737
rect 16928 26573 16974 26632
rect 16928 26468 16974 26527
rect 16928 26363 16974 26422
rect 16928 26258 16974 26317
rect 16928 26153 16974 26212
rect 16928 26048 16974 26107
rect 16928 25943 16974 26002
rect 16928 25838 16974 25897
rect 16928 25733 16974 25792
rect 16928 25628 16974 25687
rect 16928 25524 16974 25582
rect 16928 25420 16974 25478
rect 16928 25339 16974 25374
rect 17152 26783 17198 26841
rect 17152 26678 17198 26737
rect 17152 26573 17198 26632
rect 17152 26468 17198 26527
rect 17152 26363 17198 26422
rect 17152 26258 17198 26317
rect 17152 26153 17198 26212
rect 17152 26048 17198 26107
rect 17152 25943 17198 26002
rect 17152 25838 17198 25897
rect 17152 25733 17198 25792
rect 17152 25628 17198 25687
rect 17152 25524 17198 25582
rect 17152 25420 17198 25478
rect 16704 25212 16750 25270
rect 16704 25108 16750 25166
rect 16704 25004 16750 25062
rect 16704 24900 16750 24958
rect 16704 24796 16750 24854
rect 16887 25316 17015 25339
rect 16887 25300 16928 25316
rect 16974 25300 17015 25316
rect 16887 25248 16925 25300
rect 16977 25248 17015 25300
rect 16887 25212 17015 25248
rect 16887 25166 16928 25212
rect 16974 25166 17015 25212
rect 16887 25108 17015 25166
rect 16887 25082 16928 25108
rect 16974 25082 17015 25108
rect 16887 25030 16925 25082
rect 16977 25030 17015 25082
rect 16887 25004 17015 25030
rect 16887 24958 16928 25004
rect 16974 24958 17015 25004
rect 16887 24900 17015 24958
rect 16887 24864 16928 24900
rect 16974 24864 17015 24900
rect 16887 24812 16925 24864
rect 16977 24812 17015 24864
rect 16887 24796 17015 24812
rect 16887 24772 16928 24796
rect 16704 24692 16750 24750
rect 16704 24633 16750 24646
rect 16974 24772 17015 24796
rect 17152 25316 17198 25374
rect 17376 26783 17422 26842
rect 17565 26888 17680 26985
rect 17565 26842 17600 26888
rect 17646 26842 17680 26888
rect 17565 26841 17680 26842
rect 17824 26888 17870 26901
rect 17376 26678 17422 26737
rect 17376 26573 17422 26632
rect 17376 26468 17422 26527
rect 17376 26363 17422 26422
rect 17376 26258 17422 26317
rect 17376 26153 17422 26212
rect 17376 26048 17422 26107
rect 17376 25943 17422 26002
rect 17376 25838 17422 25897
rect 17376 25733 17422 25792
rect 17376 25628 17422 25687
rect 17376 25524 17422 25582
rect 17376 25420 17422 25478
rect 17376 25339 17422 25374
rect 17600 26783 17646 26841
rect 17600 26678 17646 26737
rect 17600 26573 17646 26632
rect 17600 26468 17646 26527
rect 17600 26363 17646 26422
rect 17600 26258 17646 26317
rect 17600 26153 17646 26212
rect 17600 26048 17646 26107
rect 17600 25943 17646 26002
rect 17600 25838 17646 25897
rect 17600 25733 17646 25792
rect 17600 25628 17646 25687
rect 17600 25524 17646 25582
rect 17600 25420 17646 25478
rect 17152 25212 17198 25270
rect 17152 25108 17198 25166
rect 17152 25004 17198 25062
rect 17152 24900 17198 24958
rect 17152 24796 17198 24854
rect 16928 24692 16974 24750
rect 16928 24633 16974 24646
rect 17335 25316 17463 25339
rect 17335 25300 17376 25316
rect 17422 25300 17463 25316
rect 17335 25248 17373 25300
rect 17425 25248 17463 25300
rect 17335 25212 17463 25248
rect 17335 25166 17376 25212
rect 17422 25166 17463 25212
rect 17335 25108 17463 25166
rect 17335 25082 17376 25108
rect 17422 25082 17463 25108
rect 17335 25030 17373 25082
rect 17425 25030 17463 25082
rect 17335 25004 17463 25030
rect 17335 24958 17376 25004
rect 17422 24958 17463 25004
rect 17335 24900 17463 24958
rect 17335 24864 17376 24900
rect 17422 24864 17463 24900
rect 17335 24812 17373 24864
rect 17425 24812 17463 24864
rect 17335 24796 17463 24812
rect 17335 24772 17376 24796
rect 17152 24692 17198 24750
rect 17152 24633 17198 24646
rect 17422 24772 17463 24796
rect 17600 25316 17646 25374
rect 17824 26783 17870 26842
rect 18013 26888 18128 26986
rect 18013 26842 18048 26888
rect 18094 26842 18128 26888
rect 18013 26841 18128 26842
rect 18304 27240 18419 27265
rect 18304 27194 18338 27240
rect 18384 27194 18419 27240
rect 18304 27105 18419 27194
rect 18562 27240 18608 27298
rect 18832 27513 18875 27552
rect 19010 27971 19056 27975
rect 19010 27866 19056 27925
rect 19010 27761 19056 27820
rect 19010 27656 19056 27715
rect 19010 27552 19056 27610
rect 18786 27448 18832 27506
rect 18786 27344 18832 27402
rect 18786 27265 18832 27298
rect 19191 27971 19319 27989
rect 19423 28076 19552 28122
rect 20147 28122 20185 28170
rect 20237 28170 21095 28174
rect 20237 28122 20276 28170
rect 19423 28030 19458 28076
rect 19504 28030 19552 28076
rect 19423 27975 19552 28030
rect 19191 27925 19234 27971
rect 19280 27925 19319 27971
rect 19191 27866 19319 27925
rect 19191 27823 19234 27866
rect 19280 27823 19319 27866
rect 19191 27771 19229 27823
rect 19281 27771 19319 27823
rect 19191 27761 19319 27771
rect 19191 27715 19234 27761
rect 19280 27715 19319 27761
rect 19191 27656 19319 27715
rect 19191 27610 19234 27656
rect 19280 27610 19319 27656
rect 19424 27971 19552 27975
rect 19424 27925 19458 27971
rect 19504 27956 19552 27971
rect 19424 27904 19462 27925
rect 19514 27904 19552 27956
rect 19424 27866 19552 27904
rect 19424 27820 19458 27866
rect 19504 27820 19552 27866
rect 19424 27761 19552 27820
rect 19424 27715 19458 27761
rect 19504 27738 19552 27761
rect 19424 27686 19462 27715
rect 19514 27686 19552 27738
rect 19424 27656 19552 27686
rect 19424 27646 19458 27656
rect 19191 27605 19319 27610
rect 19191 27553 19229 27605
rect 19281 27553 19319 27605
rect 19191 27552 19319 27553
rect 19191 27513 19234 27552
rect 19010 27448 19056 27506
rect 19010 27344 19056 27402
rect 18562 27181 18608 27194
rect 18752 27240 18867 27265
rect 18752 27194 18786 27240
rect 18832 27194 18867 27240
rect 18752 27105 18867 27194
rect 19010 27240 19056 27298
rect 19280 27513 19319 27552
rect 19504 27646 19552 27656
rect 19682 28076 19728 28089
rect 19682 27971 19728 28030
rect 19682 27866 19728 27925
rect 19682 27761 19728 27820
rect 19682 27656 19728 27715
rect 19458 27552 19504 27610
rect 19234 27448 19280 27506
rect 19234 27344 19280 27402
rect 19234 27265 19280 27298
rect 19458 27448 19504 27506
rect 19458 27344 19504 27402
rect 19010 27181 19056 27194
rect 19199 27240 19314 27265
rect 19199 27194 19234 27240
rect 19280 27194 19314 27240
rect 18304 26986 18867 27105
rect 18304 26888 18419 26986
rect 18751 26985 18867 26986
rect 18304 26842 18338 26888
rect 18384 26842 18419 26888
rect 18304 26841 18419 26842
rect 18562 26888 18608 26901
rect 17824 26678 17870 26737
rect 17824 26573 17870 26632
rect 17824 26468 17870 26527
rect 17824 26363 17870 26422
rect 17824 26258 17870 26317
rect 17824 26153 17870 26212
rect 17824 26048 17870 26107
rect 17824 25943 17870 26002
rect 17824 25838 17870 25897
rect 17824 25733 17870 25792
rect 17824 25628 17870 25687
rect 17824 25524 17870 25582
rect 17824 25420 17870 25478
rect 17824 25339 17870 25374
rect 18048 26783 18094 26841
rect 18048 26678 18094 26737
rect 18048 26573 18094 26632
rect 18048 26468 18094 26527
rect 18048 26363 18094 26422
rect 18048 26258 18094 26317
rect 18048 26153 18094 26212
rect 18048 26048 18094 26107
rect 18048 25943 18094 26002
rect 18048 25838 18094 25897
rect 18048 25733 18094 25792
rect 18048 25628 18094 25687
rect 18048 25524 18094 25582
rect 18048 25420 18094 25478
rect 17600 25212 17646 25270
rect 17600 25108 17646 25166
rect 17600 25004 17646 25062
rect 17600 24900 17646 24958
rect 17600 24796 17646 24854
rect 17376 24692 17422 24750
rect 17376 24633 17422 24646
rect 17783 25316 17911 25339
rect 17783 25300 17824 25316
rect 17870 25300 17911 25316
rect 17783 25248 17821 25300
rect 17873 25248 17911 25300
rect 17783 25212 17911 25248
rect 17783 25166 17824 25212
rect 17870 25166 17911 25212
rect 17783 25108 17911 25166
rect 17783 25082 17824 25108
rect 17870 25082 17911 25108
rect 17783 25030 17821 25082
rect 17873 25030 17911 25082
rect 17783 25004 17911 25030
rect 17783 24958 17824 25004
rect 17870 24958 17911 25004
rect 17783 24900 17911 24958
rect 17783 24864 17824 24900
rect 17870 24864 17911 24900
rect 17783 24812 17821 24864
rect 17873 24812 17911 24864
rect 17783 24796 17911 24812
rect 17783 24772 17824 24796
rect 17600 24692 17646 24750
rect 17600 24633 17646 24646
rect 17870 24772 17911 24796
rect 18048 25316 18094 25374
rect 18048 25212 18094 25270
rect 18048 25108 18094 25166
rect 18048 25004 18094 25062
rect 18048 24900 18094 24958
rect 18048 24796 18094 24854
rect 17824 24692 17870 24750
rect 17824 24633 17870 24646
rect 18048 24692 18094 24750
rect 18048 24633 18094 24646
rect 18338 26783 18384 26841
rect 18338 26678 18384 26737
rect 18338 26573 18384 26632
rect 18338 26468 18384 26527
rect 18338 26363 18384 26422
rect 18338 26258 18384 26317
rect 18338 26153 18384 26212
rect 18338 26048 18384 26107
rect 18338 25943 18384 26002
rect 18338 25838 18384 25897
rect 18338 25733 18384 25792
rect 18338 25628 18384 25687
rect 18338 25524 18384 25582
rect 18338 25420 18384 25478
rect 18338 25316 18384 25374
rect 18562 26783 18608 26842
rect 18752 26888 18867 26985
rect 19199 27105 19314 27194
rect 19458 27240 19504 27298
rect 19682 27552 19728 27610
rect 19682 27448 19728 27506
rect 19682 27344 19728 27402
rect 19682 27265 19728 27298
rect 19971 28076 20017 28089
rect 19971 27971 20017 28030
rect 19971 27866 20017 27925
rect 19971 27761 20017 27820
rect 19971 27656 20017 27715
rect 20147 28076 20276 28122
rect 20419 28080 20465 28089
rect 20147 28030 20195 28076
rect 20241 28030 20276 28076
rect 20147 27975 20276 28030
rect 20380 28076 20508 28080
rect 20380 28041 20419 28076
rect 20465 28041 20508 28076
rect 20380 27989 20418 28041
rect 20470 27989 20508 28041
rect 20147 27971 20275 27975
rect 20147 27956 20195 27971
rect 20147 27904 20185 27956
rect 20241 27925 20275 27971
rect 20237 27904 20275 27925
rect 20147 27866 20275 27904
rect 20147 27820 20195 27866
rect 20241 27820 20275 27866
rect 20147 27761 20275 27820
rect 20147 27738 20195 27761
rect 20147 27686 20185 27738
rect 20241 27715 20275 27761
rect 20237 27686 20275 27715
rect 20147 27656 20275 27686
rect 20147 27646 20195 27656
rect 19971 27552 20017 27610
rect 19971 27448 20017 27506
rect 19971 27344 20017 27402
rect 19971 27265 20017 27298
rect 20241 27646 20275 27656
rect 20380 27971 20508 27989
rect 20608 28076 20724 28170
rect 21056 28122 21095 28170
rect 21147 28170 21819 28174
rect 21147 28122 21185 28170
rect 20867 28080 20913 28089
rect 20608 28030 20643 28076
rect 20689 28030 20724 28076
rect 20608 27975 20724 28030
rect 20824 28076 20952 28080
rect 20824 28041 20867 28076
rect 20913 28041 20952 28076
rect 20824 27989 20862 28041
rect 20914 27989 20952 28041
rect 20380 27925 20419 27971
rect 20465 27925 20508 27971
rect 20380 27866 20508 27925
rect 20380 27823 20419 27866
rect 20465 27823 20508 27866
rect 20380 27771 20418 27823
rect 20470 27771 20508 27823
rect 20380 27761 20508 27771
rect 20380 27715 20419 27761
rect 20465 27715 20508 27761
rect 20380 27656 20508 27715
rect 20195 27552 20241 27610
rect 20380 27610 20419 27656
rect 20465 27610 20508 27656
rect 20380 27605 20508 27610
rect 20380 27553 20418 27605
rect 20470 27553 20508 27605
rect 20380 27552 20508 27553
rect 20380 27513 20419 27552
rect 20195 27448 20241 27506
rect 20195 27344 20241 27402
rect 19458 27181 19504 27194
rect 19647 27240 19762 27265
rect 19647 27194 19682 27240
rect 19728 27194 19762 27240
rect 19647 27105 19762 27194
rect 19199 26986 19762 27105
rect 19199 26985 19315 26986
rect 18752 26842 18786 26888
rect 18832 26842 18867 26888
rect 18752 26841 18867 26842
rect 19010 26888 19056 26901
rect 18562 26678 18608 26737
rect 18562 26573 18608 26632
rect 18562 26468 18608 26527
rect 18562 26363 18608 26422
rect 18562 26258 18608 26317
rect 18562 26153 18608 26212
rect 18562 26048 18608 26107
rect 18562 25943 18608 26002
rect 18562 25838 18608 25897
rect 18562 25733 18608 25792
rect 18562 25628 18608 25687
rect 18562 25524 18608 25582
rect 18562 25420 18608 25478
rect 18562 25339 18608 25374
rect 18786 26783 18832 26841
rect 18786 26678 18832 26737
rect 18786 26573 18832 26632
rect 18786 26468 18832 26527
rect 18786 26363 18832 26422
rect 18786 26258 18832 26317
rect 18786 26153 18832 26212
rect 18786 26048 18832 26107
rect 18786 25943 18832 26002
rect 18786 25838 18832 25897
rect 18786 25733 18832 25792
rect 18786 25628 18832 25687
rect 18786 25524 18832 25582
rect 18786 25420 18832 25478
rect 18338 25212 18384 25270
rect 18338 25108 18384 25166
rect 18338 25004 18384 25062
rect 18338 24900 18384 24958
rect 18338 24796 18384 24854
rect 18521 25316 18649 25339
rect 18521 25300 18562 25316
rect 18608 25300 18649 25316
rect 18521 25248 18559 25300
rect 18611 25248 18649 25300
rect 18521 25212 18649 25248
rect 18521 25166 18562 25212
rect 18608 25166 18649 25212
rect 18521 25108 18649 25166
rect 18521 25082 18562 25108
rect 18608 25082 18649 25108
rect 18521 25030 18559 25082
rect 18611 25030 18649 25082
rect 18521 25004 18649 25030
rect 18521 24958 18562 25004
rect 18608 24958 18649 25004
rect 18521 24900 18649 24958
rect 18521 24864 18562 24900
rect 18608 24864 18649 24900
rect 18521 24812 18559 24864
rect 18611 24812 18649 24864
rect 18521 24796 18649 24812
rect 18521 24772 18562 24796
rect 18338 24692 18384 24750
rect 18338 24633 18384 24646
rect 18608 24772 18649 24796
rect 18786 25316 18832 25374
rect 19010 26783 19056 26842
rect 19199 26888 19314 26985
rect 19199 26842 19234 26888
rect 19280 26842 19314 26888
rect 19199 26841 19314 26842
rect 19458 26888 19504 26901
rect 19010 26678 19056 26737
rect 19010 26573 19056 26632
rect 19010 26468 19056 26527
rect 19010 26363 19056 26422
rect 19010 26258 19056 26317
rect 19010 26153 19056 26212
rect 19010 26048 19056 26107
rect 19010 25943 19056 26002
rect 19010 25838 19056 25897
rect 19010 25733 19056 25792
rect 19010 25628 19056 25687
rect 19010 25524 19056 25582
rect 19010 25420 19056 25478
rect 19010 25339 19056 25374
rect 19234 26783 19280 26841
rect 19234 26678 19280 26737
rect 19234 26573 19280 26632
rect 19234 26468 19280 26527
rect 19234 26363 19280 26422
rect 19234 26258 19280 26317
rect 19234 26153 19280 26212
rect 19234 26048 19280 26107
rect 19234 25943 19280 26002
rect 19234 25838 19280 25897
rect 19234 25733 19280 25792
rect 19234 25628 19280 25687
rect 19234 25524 19280 25582
rect 19234 25420 19280 25478
rect 18786 25212 18832 25270
rect 18786 25108 18832 25166
rect 18786 25004 18832 25062
rect 18786 24900 18832 24958
rect 18786 24796 18832 24854
rect 18562 24692 18608 24750
rect 18562 24633 18608 24646
rect 18969 25316 19097 25339
rect 18969 25300 19010 25316
rect 19056 25300 19097 25316
rect 18969 25248 19007 25300
rect 19059 25248 19097 25300
rect 18969 25212 19097 25248
rect 18969 25166 19010 25212
rect 19056 25166 19097 25212
rect 18969 25108 19097 25166
rect 18969 25082 19010 25108
rect 19056 25082 19097 25108
rect 18969 25030 19007 25082
rect 19059 25030 19097 25082
rect 18969 25004 19097 25030
rect 18969 24958 19010 25004
rect 19056 24958 19097 25004
rect 18969 24900 19097 24958
rect 18969 24864 19010 24900
rect 19056 24864 19097 24900
rect 18969 24812 19007 24864
rect 19059 24812 19097 24864
rect 18969 24796 19097 24812
rect 18969 24772 19010 24796
rect 18786 24692 18832 24750
rect 18786 24633 18832 24646
rect 19056 24772 19097 24796
rect 19234 25316 19280 25374
rect 19458 26783 19504 26842
rect 19647 26888 19762 26986
rect 19647 26842 19682 26888
rect 19728 26842 19762 26888
rect 19647 26841 19762 26842
rect 19937 27240 20052 27265
rect 19937 27194 19971 27240
rect 20017 27194 20052 27240
rect 19937 27105 20052 27194
rect 20195 27240 20241 27298
rect 20465 27513 20508 27552
rect 20643 27971 20689 27975
rect 20643 27866 20689 27925
rect 20643 27761 20689 27820
rect 20643 27656 20689 27715
rect 20643 27552 20689 27610
rect 20419 27448 20465 27506
rect 20419 27344 20465 27402
rect 20419 27265 20465 27298
rect 20824 27971 20952 27989
rect 21056 28076 21185 28122
rect 21781 28122 21819 28170
rect 21871 28170 22729 28174
rect 21871 28122 21910 28170
rect 21056 28030 21091 28076
rect 21137 28030 21185 28076
rect 21056 27975 21185 28030
rect 20824 27925 20867 27971
rect 20913 27925 20952 27971
rect 20824 27866 20952 27925
rect 20824 27823 20867 27866
rect 20913 27823 20952 27866
rect 20824 27771 20862 27823
rect 20914 27771 20952 27823
rect 20824 27761 20952 27771
rect 20824 27715 20867 27761
rect 20913 27715 20952 27761
rect 20824 27656 20952 27715
rect 20824 27610 20867 27656
rect 20913 27610 20952 27656
rect 21057 27971 21185 27975
rect 21057 27925 21091 27971
rect 21137 27956 21185 27971
rect 21057 27904 21095 27925
rect 21147 27904 21185 27956
rect 21057 27866 21185 27904
rect 21057 27820 21091 27866
rect 21137 27820 21185 27866
rect 21057 27761 21185 27820
rect 21057 27715 21091 27761
rect 21137 27738 21185 27761
rect 21057 27686 21095 27715
rect 21147 27686 21185 27738
rect 21057 27656 21185 27686
rect 21057 27646 21091 27656
rect 20824 27605 20952 27610
rect 20824 27553 20862 27605
rect 20914 27553 20952 27605
rect 20824 27552 20952 27553
rect 20824 27513 20867 27552
rect 20643 27448 20689 27506
rect 20643 27344 20689 27402
rect 20195 27181 20241 27194
rect 20385 27240 20500 27265
rect 20385 27194 20419 27240
rect 20465 27194 20500 27240
rect 20385 27105 20500 27194
rect 20643 27240 20689 27298
rect 20913 27513 20952 27552
rect 21137 27646 21185 27656
rect 21315 28076 21361 28089
rect 21315 27971 21361 28030
rect 21315 27866 21361 27925
rect 21315 27761 21361 27820
rect 21315 27656 21361 27715
rect 21091 27552 21137 27610
rect 20867 27448 20913 27506
rect 20867 27344 20913 27402
rect 20867 27265 20913 27298
rect 21091 27448 21137 27506
rect 21091 27344 21137 27402
rect 20643 27181 20689 27194
rect 20832 27240 20947 27265
rect 20832 27194 20867 27240
rect 20913 27194 20947 27240
rect 19937 26986 20500 27105
rect 19937 26888 20052 26986
rect 20384 26985 20500 26986
rect 19937 26842 19971 26888
rect 20017 26842 20052 26888
rect 19937 26841 20052 26842
rect 20195 26888 20241 26901
rect 19458 26678 19504 26737
rect 19458 26573 19504 26632
rect 19458 26468 19504 26527
rect 19458 26363 19504 26422
rect 19458 26258 19504 26317
rect 19458 26153 19504 26212
rect 19458 26048 19504 26107
rect 19458 25943 19504 26002
rect 19458 25838 19504 25897
rect 19458 25733 19504 25792
rect 19458 25628 19504 25687
rect 19458 25524 19504 25582
rect 19458 25420 19504 25478
rect 19458 25339 19504 25374
rect 19682 26783 19728 26841
rect 19682 26678 19728 26737
rect 19682 26573 19728 26632
rect 19682 26468 19728 26527
rect 19682 26363 19728 26422
rect 19682 26258 19728 26317
rect 19682 26153 19728 26212
rect 19682 26048 19728 26107
rect 19682 25943 19728 26002
rect 19682 25838 19728 25897
rect 19682 25733 19728 25792
rect 19682 25628 19728 25687
rect 19682 25524 19728 25582
rect 19682 25420 19728 25478
rect 19234 25212 19280 25270
rect 19234 25108 19280 25166
rect 19234 25004 19280 25062
rect 19234 24900 19280 24958
rect 19234 24796 19280 24854
rect 19010 24692 19056 24750
rect 19010 24633 19056 24646
rect 19417 25316 19545 25339
rect 19417 25300 19458 25316
rect 19504 25300 19545 25316
rect 19417 25248 19455 25300
rect 19507 25248 19545 25300
rect 19417 25212 19545 25248
rect 19417 25166 19458 25212
rect 19504 25166 19545 25212
rect 19417 25108 19545 25166
rect 19417 25082 19458 25108
rect 19504 25082 19545 25108
rect 19417 25030 19455 25082
rect 19507 25030 19545 25082
rect 19417 25004 19545 25030
rect 19417 24958 19458 25004
rect 19504 24958 19545 25004
rect 19417 24900 19545 24958
rect 19417 24864 19458 24900
rect 19504 24864 19545 24900
rect 19417 24812 19455 24864
rect 19507 24812 19545 24864
rect 19417 24796 19545 24812
rect 19417 24772 19458 24796
rect 19234 24692 19280 24750
rect 19234 24633 19280 24646
rect 19504 24772 19545 24796
rect 19682 25316 19728 25374
rect 19682 25212 19728 25270
rect 19682 25108 19728 25166
rect 19682 25004 19728 25062
rect 19682 24900 19728 24958
rect 19682 24796 19728 24854
rect 19458 24692 19504 24750
rect 19458 24633 19504 24646
rect 19682 24692 19728 24750
rect 19682 24633 19728 24646
rect 19971 26783 20017 26841
rect 19971 26678 20017 26737
rect 19971 26573 20017 26632
rect 19971 26468 20017 26527
rect 19971 26363 20017 26422
rect 19971 26258 20017 26317
rect 19971 26153 20017 26212
rect 19971 26048 20017 26107
rect 19971 25943 20017 26002
rect 19971 25838 20017 25897
rect 19971 25733 20017 25792
rect 19971 25628 20017 25687
rect 19971 25524 20017 25582
rect 19971 25420 20017 25478
rect 19971 25316 20017 25374
rect 20195 26783 20241 26842
rect 20385 26888 20500 26985
rect 20832 27105 20947 27194
rect 21091 27240 21137 27298
rect 21315 27552 21361 27610
rect 21315 27448 21361 27506
rect 21315 27344 21361 27402
rect 21315 27265 21361 27298
rect 21605 28076 21651 28089
rect 21605 27971 21651 28030
rect 21605 27866 21651 27925
rect 21605 27761 21651 27820
rect 21605 27656 21651 27715
rect 21781 28076 21910 28122
rect 22053 28080 22099 28089
rect 21781 28030 21829 28076
rect 21875 28030 21910 28076
rect 21781 27975 21910 28030
rect 22014 28076 22142 28080
rect 22014 28041 22053 28076
rect 22099 28041 22142 28076
rect 22014 27989 22052 28041
rect 22104 27989 22142 28041
rect 21781 27971 21909 27975
rect 21781 27956 21829 27971
rect 21781 27904 21819 27956
rect 21875 27925 21909 27971
rect 21871 27904 21909 27925
rect 21781 27866 21909 27904
rect 21781 27820 21829 27866
rect 21875 27820 21909 27866
rect 21781 27761 21909 27820
rect 21781 27738 21829 27761
rect 21781 27686 21819 27738
rect 21875 27715 21909 27761
rect 21871 27686 21909 27715
rect 21781 27656 21909 27686
rect 21781 27646 21829 27656
rect 21605 27552 21651 27610
rect 21605 27448 21651 27506
rect 21605 27344 21651 27402
rect 21605 27265 21651 27298
rect 21875 27646 21909 27656
rect 22014 27971 22142 27989
rect 22242 28076 22358 28170
rect 22690 28122 22729 28170
rect 22781 28170 23118 28174
rect 23749 28190 23878 28314
rect 23749 28183 23797 28190
rect 22781 28122 22819 28170
rect 22501 28080 22547 28089
rect 22242 28030 22277 28076
rect 22323 28030 22358 28076
rect 22242 27975 22358 28030
rect 22458 28076 22586 28080
rect 22458 28041 22501 28076
rect 22547 28041 22586 28076
rect 22458 27989 22496 28041
rect 22548 27989 22586 28041
rect 22014 27925 22053 27971
rect 22099 27925 22142 27971
rect 22014 27866 22142 27925
rect 22014 27823 22053 27866
rect 22099 27823 22142 27866
rect 22014 27771 22052 27823
rect 22104 27771 22142 27823
rect 22014 27761 22142 27771
rect 22014 27715 22053 27761
rect 22099 27715 22142 27761
rect 22014 27656 22142 27715
rect 21829 27552 21875 27610
rect 22014 27610 22053 27656
rect 22099 27610 22142 27656
rect 22014 27605 22142 27610
rect 22014 27553 22052 27605
rect 22104 27553 22142 27605
rect 22014 27552 22142 27553
rect 22014 27513 22053 27552
rect 21829 27448 21875 27506
rect 21829 27344 21875 27402
rect 21091 27181 21137 27194
rect 21280 27240 21395 27265
rect 21280 27194 21315 27240
rect 21361 27194 21395 27240
rect 21280 27105 21395 27194
rect 20832 26986 21395 27105
rect 20832 26985 20948 26986
rect 20385 26842 20419 26888
rect 20465 26842 20500 26888
rect 20385 26841 20500 26842
rect 20643 26888 20689 26901
rect 20195 26678 20241 26737
rect 20195 26573 20241 26632
rect 20195 26468 20241 26527
rect 20195 26363 20241 26422
rect 20195 26258 20241 26317
rect 20195 26153 20241 26212
rect 20195 26048 20241 26107
rect 20195 25943 20241 26002
rect 20195 25838 20241 25897
rect 20195 25733 20241 25792
rect 20195 25628 20241 25687
rect 20195 25524 20241 25582
rect 20195 25420 20241 25478
rect 20195 25339 20241 25374
rect 20419 26783 20465 26841
rect 20419 26678 20465 26737
rect 20419 26573 20465 26632
rect 20419 26468 20465 26527
rect 20419 26363 20465 26422
rect 20419 26258 20465 26317
rect 20419 26153 20465 26212
rect 20419 26048 20465 26107
rect 20419 25943 20465 26002
rect 20419 25838 20465 25897
rect 20419 25733 20465 25792
rect 20419 25628 20465 25687
rect 20419 25524 20465 25582
rect 20419 25420 20465 25478
rect 19971 25212 20017 25270
rect 19971 25108 20017 25166
rect 19971 25004 20017 25062
rect 19971 24900 20017 24958
rect 19971 24796 20017 24854
rect 20154 25316 20282 25339
rect 20154 25300 20195 25316
rect 20241 25300 20282 25316
rect 20154 25248 20192 25300
rect 20244 25248 20282 25300
rect 20154 25212 20282 25248
rect 20154 25166 20195 25212
rect 20241 25166 20282 25212
rect 20154 25108 20282 25166
rect 20154 25082 20195 25108
rect 20241 25082 20282 25108
rect 20154 25030 20192 25082
rect 20244 25030 20282 25082
rect 20154 25004 20282 25030
rect 20154 24958 20195 25004
rect 20241 24958 20282 25004
rect 20154 24900 20282 24958
rect 20154 24864 20195 24900
rect 20241 24864 20282 24900
rect 20154 24812 20192 24864
rect 20244 24812 20282 24864
rect 20154 24796 20282 24812
rect 20154 24772 20195 24796
rect 19971 24692 20017 24750
rect 19971 24633 20017 24646
rect 20241 24772 20282 24796
rect 20419 25316 20465 25374
rect 20643 26783 20689 26842
rect 20832 26888 20947 26985
rect 20832 26842 20867 26888
rect 20913 26842 20947 26888
rect 20832 26841 20947 26842
rect 21091 26888 21137 26901
rect 20643 26678 20689 26737
rect 20643 26573 20689 26632
rect 20643 26468 20689 26527
rect 20643 26363 20689 26422
rect 20643 26258 20689 26317
rect 20643 26153 20689 26212
rect 20643 26048 20689 26107
rect 20643 25943 20689 26002
rect 20643 25838 20689 25897
rect 20643 25733 20689 25792
rect 20643 25628 20689 25687
rect 20643 25524 20689 25582
rect 20643 25420 20689 25478
rect 20643 25339 20689 25374
rect 20867 26783 20913 26841
rect 20867 26678 20913 26737
rect 20867 26573 20913 26632
rect 20867 26468 20913 26527
rect 20867 26363 20913 26422
rect 20867 26258 20913 26317
rect 20867 26153 20913 26212
rect 20867 26048 20913 26107
rect 20867 25943 20913 26002
rect 20867 25838 20913 25897
rect 20867 25733 20913 25792
rect 20867 25628 20913 25687
rect 20867 25524 20913 25582
rect 20867 25420 20913 25478
rect 20419 25212 20465 25270
rect 20419 25108 20465 25166
rect 20419 25004 20465 25062
rect 20419 24900 20465 24958
rect 20419 24796 20465 24854
rect 20195 24692 20241 24750
rect 20195 24633 20241 24646
rect 20602 25316 20730 25339
rect 20602 25300 20643 25316
rect 20689 25300 20730 25316
rect 20602 25248 20640 25300
rect 20692 25248 20730 25300
rect 20602 25212 20730 25248
rect 20602 25166 20643 25212
rect 20689 25166 20730 25212
rect 20602 25108 20730 25166
rect 20602 25082 20643 25108
rect 20689 25082 20730 25108
rect 20602 25030 20640 25082
rect 20692 25030 20730 25082
rect 20602 25004 20730 25030
rect 20602 24958 20643 25004
rect 20689 24958 20730 25004
rect 20602 24900 20730 24958
rect 20602 24864 20643 24900
rect 20689 24864 20730 24900
rect 20602 24812 20640 24864
rect 20692 24812 20730 24864
rect 20602 24796 20730 24812
rect 20602 24772 20643 24796
rect 20419 24692 20465 24750
rect 20419 24633 20465 24646
rect 20689 24772 20730 24796
rect 20867 25316 20913 25374
rect 21091 26783 21137 26842
rect 21280 26888 21395 26986
rect 21280 26842 21315 26888
rect 21361 26842 21395 26888
rect 21280 26841 21395 26842
rect 21571 27240 21686 27265
rect 21571 27194 21605 27240
rect 21651 27194 21686 27240
rect 21571 27105 21686 27194
rect 21829 27240 21875 27298
rect 22099 27513 22142 27552
rect 22277 27971 22323 27975
rect 22277 27866 22323 27925
rect 22277 27761 22323 27820
rect 22277 27656 22323 27715
rect 22277 27552 22323 27610
rect 22053 27448 22099 27506
rect 22053 27344 22099 27402
rect 22053 27265 22099 27298
rect 22458 27971 22586 27989
rect 22690 28076 22819 28122
rect 23749 28131 23787 28183
rect 23843 28144 23878 28190
rect 23839 28131 23878 28144
rect 24021 28190 24067 28203
rect 24021 28135 24067 28144
rect 24188 28190 24326 28314
rect 25572 28292 25610 28314
rect 25662 28314 28525 28344
rect 25662 28292 25700 28314
rect 24188 28183 24245 28190
rect 22690 28030 22725 28076
rect 22771 28030 22819 28076
rect 22690 27975 22819 28030
rect 22458 27925 22501 27971
rect 22547 27925 22586 27971
rect 22458 27866 22586 27925
rect 22458 27823 22501 27866
rect 22547 27823 22586 27866
rect 22458 27771 22496 27823
rect 22548 27771 22586 27823
rect 22458 27761 22586 27771
rect 22458 27715 22501 27761
rect 22547 27715 22586 27761
rect 22458 27656 22586 27715
rect 22458 27610 22501 27656
rect 22547 27610 22586 27656
rect 22691 27971 22819 27975
rect 22691 27925 22725 27971
rect 22771 27956 22819 27971
rect 22691 27904 22729 27925
rect 22781 27904 22819 27956
rect 22691 27866 22819 27904
rect 22691 27820 22725 27866
rect 22771 27820 22819 27866
rect 22691 27761 22819 27820
rect 22691 27715 22725 27761
rect 22771 27738 22819 27761
rect 22691 27686 22729 27715
rect 22781 27686 22819 27738
rect 22691 27656 22819 27686
rect 22691 27646 22725 27656
rect 22458 27605 22586 27610
rect 22458 27553 22496 27605
rect 22548 27553 22586 27605
rect 22458 27552 22586 27553
rect 22458 27513 22501 27552
rect 22277 27448 22323 27506
rect 22277 27344 22323 27402
rect 21829 27181 21875 27194
rect 22019 27240 22134 27265
rect 22019 27194 22053 27240
rect 22099 27194 22134 27240
rect 22019 27105 22134 27194
rect 22277 27240 22323 27298
rect 22547 27513 22586 27552
rect 22771 27646 22819 27656
rect 22949 28076 22995 28089
rect 22949 27971 22995 28030
rect 22949 27866 22995 27925
rect 23749 28087 23878 28131
rect 23749 28041 23797 28087
rect 23843 28041 23878 28087
rect 23749 27984 23878 28041
rect 23749 27965 23797 27984
rect 23749 27913 23787 27965
rect 23843 27938 23878 27984
rect 23839 27913 23878 27938
rect 23749 27880 23878 27913
rect 23749 27873 23797 27880
rect 23762 27834 23797 27873
rect 23843 27834 23878 27880
rect 23762 27829 23878 27834
rect 23986 28087 24102 28135
rect 23986 28041 24021 28087
rect 24067 28041 24102 28087
rect 23986 27984 24102 28041
rect 23986 27938 24021 27984
rect 24067 27938 24102 27984
rect 23986 27880 24102 27938
rect 23986 27834 24021 27880
rect 24067 27834 24102 27880
rect 24188 28131 24226 28183
rect 24291 28144 24326 28190
rect 24278 28131 24326 28144
rect 24188 28087 24326 28131
rect 24188 28041 24245 28087
rect 24291 28041 24326 28087
rect 24188 27984 24326 28041
rect 24188 27965 24245 27984
rect 24188 27913 24226 27965
rect 24291 27938 24326 27984
rect 24278 27913 24326 27938
rect 24188 27880 24326 27913
rect 24188 27873 24245 27880
rect 23797 27821 23843 27829
rect 22949 27761 22995 27820
rect 22949 27656 22995 27715
rect 22725 27552 22771 27610
rect 22501 27448 22547 27506
rect 22501 27344 22547 27402
rect 22501 27265 22547 27298
rect 22725 27448 22771 27506
rect 22725 27344 22771 27402
rect 22277 27181 22323 27194
rect 22466 27240 22581 27265
rect 22466 27194 22501 27240
rect 22547 27194 22581 27240
rect 21571 26986 22134 27105
rect 21571 26888 21686 26986
rect 22018 26985 22134 26986
rect 21571 26842 21605 26888
rect 21651 26842 21686 26888
rect 21571 26841 21686 26842
rect 21829 26888 21875 26901
rect 21091 26678 21137 26737
rect 21091 26573 21137 26632
rect 21091 26468 21137 26527
rect 21091 26363 21137 26422
rect 21091 26258 21137 26317
rect 21091 26153 21137 26212
rect 21091 26048 21137 26107
rect 21091 25943 21137 26002
rect 21091 25838 21137 25897
rect 21091 25733 21137 25792
rect 21091 25628 21137 25687
rect 21091 25524 21137 25582
rect 21091 25420 21137 25478
rect 21091 25339 21137 25374
rect 21315 26783 21361 26841
rect 21315 26678 21361 26737
rect 21315 26573 21361 26632
rect 21315 26468 21361 26527
rect 21315 26363 21361 26422
rect 21315 26258 21361 26317
rect 21315 26153 21361 26212
rect 21315 26048 21361 26107
rect 21315 25943 21361 26002
rect 21315 25838 21361 25897
rect 21315 25733 21361 25792
rect 21315 25628 21361 25687
rect 21315 25524 21361 25582
rect 21315 25420 21361 25478
rect 20867 25212 20913 25270
rect 20867 25108 20913 25166
rect 20867 25004 20913 25062
rect 20867 24900 20913 24958
rect 20867 24796 20913 24854
rect 20643 24692 20689 24750
rect 20643 24633 20689 24646
rect 21050 25316 21178 25339
rect 21050 25300 21091 25316
rect 21137 25300 21178 25316
rect 21050 25248 21088 25300
rect 21140 25248 21178 25300
rect 21050 25212 21178 25248
rect 21050 25166 21091 25212
rect 21137 25166 21178 25212
rect 21050 25108 21178 25166
rect 21050 25082 21091 25108
rect 21137 25082 21178 25108
rect 21050 25030 21088 25082
rect 21140 25030 21178 25082
rect 21050 25004 21178 25030
rect 21050 24958 21091 25004
rect 21137 24958 21178 25004
rect 21050 24900 21178 24958
rect 21050 24864 21091 24900
rect 21137 24864 21178 24900
rect 21050 24812 21088 24864
rect 21140 24812 21178 24864
rect 21050 24796 21178 24812
rect 21050 24772 21091 24796
rect 20867 24692 20913 24750
rect 20867 24633 20913 24646
rect 21137 24772 21178 24796
rect 21315 25316 21361 25374
rect 21315 25212 21361 25270
rect 21315 25108 21361 25166
rect 21315 25004 21361 25062
rect 21315 24900 21361 24958
rect 21315 24796 21361 24854
rect 21091 24692 21137 24750
rect 21091 24633 21137 24646
rect 21315 24692 21361 24750
rect 21315 24633 21361 24646
rect 21605 26783 21651 26841
rect 21605 26678 21651 26737
rect 21605 26573 21651 26632
rect 21605 26468 21651 26527
rect 21605 26363 21651 26422
rect 21605 26258 21651 26317
rect 21605 26153 21651 26212
rect 21605 26048 21651 26107
rect 21605 25943 21651 26002
rect 21605 25838 21651 25897
rect 21605 25733 21651 25792
rect 21605 25628 21651 25687
rect 21605 25524 21651 25582
rect 21605 25420 21651 25478
rect 21605 25316 21651 25374
rect 21829 26783 21875 26842
rect 22019 26888 22134 26985
rect 22466 27105 22581 27194
rect 22725 27240 22771 27298
rect 22949 27552 22995 27610
rect 23560 27695 23900 27736
rect 23560 27643 23598 27695
rect 23650 27694 23810 27695
rect 23862 27694 23900 27695
rect 23650 27648 23661 27694
rect 23707 27648 23810 27694
rect 23865 27648 23900 27694
rect 23650 27643 23810 27648
rect 23862 27643 23900 27648
rect 23560 27603 23900 27643
rect 23986 27733 24102 27834
rect 24210 27834 24245 27873
rect 24291 27834 24326 27880
rect 24410 28185 24534 28225
rect 24410 28133 24446 28185
rect 24498 28133 24534 28185
rect 24410 28037 24534 28133
rect 25572 28126 25700 28292
rect 24410 27897 24423 28037
rect 24469 27967 24534 28037
rect 25392 28076 25438 28089
rect 24498 27915 24534 27967
rect 24469 27897 24534 27915
rect 24410 27875 24534 27897
rect 24210 27829 24326 27834
rect 25356 27830 25392 27999
rect 25572 28074 25610 28126
rect 25438 27830 25472 27999
rect 24245 27821 24291 27829
rect 23986 27614 24326 27733
rect 25356 27692 25472 27830
rect 25572 27908 25616 28074
rect 25572 27856 25610 27908
rect 25572 27830 25616 27856
rect 25662 27830 25700 28126
rect 25572 27816 25700 27830
rect 26606 27693 26730 27726
rect 26604 27692 26733 27693
rect 25356 27686 26733 27692
rect 22949 27448 22995 27506
rect 23762 27418 23878 27500
rect 22949 27344 22995 27402
rect 22949 27265 22995 27298
rect 23751 27382 23878 27418
rect 23751 27378 23797 27382
rect 23751 27326 23787 27378
rect 23843 27336 23878 27382
rect 23839 27326 23878 27336
rect 22725 27181 22771 27194
rect 22914 27240 23029 27265
rect 22914 27194 22949 27240
rect 22995 27194 23029 27240
rect 22914 27105 23029 27194
rect 22466 26986 23029 27105
rect 23751 27178 23878 27326
rect 23751 27160 23797 27178
rect 23751 27108 23787 27160
rect 23843 27132 23878 27178
rect 23839 27108 23878 27132
rect 23751 27095 23878 27108
rect 24210 27382 24326 27614
rect 24560 27673 24740 27685
rect 24560 27621 24572 27673
rect 24728 27666 24740 27673
rect 24560 27620 24683 27621
rect 24729 27620 24740 27666
rect 24560 27609 24740 27620
rect 25356 27634 26642 27686
rect 26694 27634 26733 27686
rect 25356 27559 26733 27634
rect 24210 27336 24245 27382
rect 24291 27336 24326 27382
rect 24210 27178 24326 27336
rect 24210 27132 24245 27178
rect 24291 27132 24326 27178
rect 23751 27068 23875 27095
rect 22466 26985 22582 26986
rect 22019 26842 22053 26888
rect 22099 26842 22134 26888
rect 22019 26841 22134 26842
rect 22277 26888 22323 26901
rect 21829 26678 21875 26737
rect 21829 26573 21875 26632
rect 21829 26468 21875 26527
rect 21829 26363 21875 26422
rect 21829 26258 21875 26317
rect 21829 26153 21875 26212
rect 21829 26048 21875 26107
rect 21829 25943 21875 26002
rect 21829 25838 21875 25897
rect 21829 25733 21875 25792
rect 21829 25628 21875 25687
rect 21829 25524 21875 25582
rect 21829 25420 21875 25478
rect 21829 25339 21875 25374
rect 22053 26783 22099 26841
rect 22053 26678 22099 26737
rect 22053 26573 22099 26632
rect 22053 26468 22099 26527
rect 22053 26363 22099 26422
rect 22053 26258 22099 26317
rect 22053 26153 22099 26212
rect 22053 26048 22099 26107
rect 22053 25943 22099 26002
rect 22053 25838 22099 25897
rect 22053 25733 22099 25792
rect 22053 25628 22099 25687
rect 22053 25524 22099 25582
rect 22053 25420 22099 25478
rect 21605 25212 21651 25270
rect 21605 25108 21651 25166
rect 21605 25004 21651 25062
rect 21605 24900 21651 24958
rect 21605 24796 21651 24854
rect 21788 25316 21916 25339
rect 21788 25300 21829 25316
rect 21875 25300 21916 25316
rect 21788 25248 21826 25300
rect 21878 25248 21916 25300
rect 21788 25212 21916 25248
rect 21788 25166 21829 25212
rect 21875 25166 21916 25212
rect 21788 25108 21916 25166
rect 21788 25082 21829 25108
rect 21875 25082 21916 25108
rect 21788 25030 21826 25082
rect 21878 25030 21916 25082
rect 21788 25004 21916 25030
rect 21788 24958 21829 25004
rect 21875 24958 21916 25004
rect 21788 24900 21916 24958
rect 21788 24864 21829 24900
rect 21875 24864 21916 24900
rect 21788 24812 21826 24864
rect 21878 24812 21916 24864
rect 21788 24796 21916 24812
rect 21788 24772 21829 24796
rect 21605 24692 21651 24750
rect 21605 24633 21651 24646
rect 21875 24772 21916 24796
rect 22053 25316 22099 25374
rect 22277 26783 22323 26842
rect 22466 26888 22581 26985
rect 22466 26842 22501 26888
rect 22547 26842 22581 26888
rect 22466 26841 22581 26842
rect 22725 26888 22771 26901
rect 22277 26678 22323 26737
rect 22277 26573 22323 26632
rect 22277 26468 22323 26527
rect 22277 26363 22323 26422
rect 22277 26258 22323 26317
rect 22277 26153 22323 26212
rect 22277 26048 22323 26107
rect 22277 25943 22323 26002
rect 22277 25838 22323 25897
rect 22277 25733 22323 25792
rect 22277 25628 22323 25687
rect 22277 25524 22323 25582
rect 22277 25420 22323 25478
rect 22277 25339 22323 25374
rect 22501 26783 22547 26841
rect 22501 26678 22547 26737
rect 22501 26573 22547 26632
rect 22501 26468 22547 26527
rect 22501 26363 22547 26422
rect 22501 26258 22547 26317
rect 22501 26153 22547 26212
rect 22501 26048 22547 26107
rect 22501 25943 22547 26002
rect 22501 25838 22547 25897
rect 22501 25733 22547 25792
rect 22501 25628 22547 25687
rect 22501 25524 22547 25582
rect 22501 25420 22547 25478
rect 22053 25212 22099 25270
rect 22053 25108 22099 25166
rect 22053 25004 22099 25062
rect 22053 24900 22099 24958
rect 22053 24796 22099 24854
rect 21829 24692 21875 24750
rect 21829 24633 21875 24646
rect 22236 25316 22364 25339
rect 22236 25300 22277 25316
rect 22323 25300 22364 25316
rect 22236 25248 22274 25300
rect 22326 25248 22364 25300
rect 22236 25212 22364 25248
rect 22236 25166 22277 25212
rect 22323 25166 22364 25212
rect 22236 25108 22364 25166
rect 22236 25082 22277 25108
rect 22323 25082 22364 25108
rect 22236 25030 22274 25082
rect 22326 25030 22364 25082
rect 22236 25004 22364 25030
rect 22236 24958 22277 25004
rect 22323 24958 22364 25004
rect 22236 24900 22364 24958
rect 22236 24864 22277 24900
rect 22323 24864 22364 24900
rect 22236 24812 22274 24864
rect 22326 24812 22364 24864
rect 22236 24796 22364 24812
rect 22236 24772 22277 24796
rect 22053 24692 22099 24750
rect 22053 24633 22099 24646
rect 22323 24772 22364 24796
rect 22501 25316 22547 25374
rect 22725 26783 22771 26842
rect 22914 26888 23029 26986
rect 24210 27015 24326 27132
rect 24658 27432 24774 27500
rect 24937 27437 25061 27477
rect 24937 27432 24973 27437
rect 24658 27385 24973 27432
rect 25025 27432 25061 27437
rect 25273 27432 25319 27442
rect 25025 27429 25354 27432
rect 25025 27385 25273 27429
rect 24658 27384 25273 27385
rect 24658 27382 24978 27384
rect 24658 27336 24693 27382
rect 24739 27336 24978 27382
rect 24658 27244 24978 27336
rect 25024 27383 25273 27384
rect 25319 27383 25354 27429
rect 25024 27294 25354 27383
rect 25024 27248 25273 27294
rect 25319 27248 25354 27294
rect 25024 27244 25354 27248
rect 24658 27219 25354 27244
rect 24658 27178 24973 27219
rect 24658 27132 24693 27178
rect 24739 27167 24973 27178
rect 25025 27167 25354 27219
rect 25462 27429 25578 27559
rect 26606 27468 26730 27559
rect 25721 27432 25767 27442
rect 25462 27383 25497 27429
rect 25543 27383 25578 27429
rect 25462 27294 25578 27383
rect 25462 27248 25497 27294
rect 25543 27248 25578 27294
rect 25462 27197 25578 27248
rect 25686 27429 26091 27432
rect 25686 27383 25721 27429
rect 25767 27392 26091 27429
rect 25767 27383 26001 27392
rect 25686 27340 26001 27383
rect 26053 27340 26091 27392
rect 26606 27416 26642 27468
rect 26694 27416 26730 27468
rect 26606 27376 26730 27416
rect 25686 27328 26091 27340
rect 25686 27294 26008 27328
rect 25686 27248 25721 27294
rect 25767 27248 26008 27294
rect 24739 27159 25354 27167
rect 24739 27132 25273 27159
rect 24658 27113 25273 27132
rect 25319 27113 25354 27159
rect 24658 27108 25354 27113
rect 25497 27159 25543 27197
rect 24658 27095 24774 27108
rect 25273 27100 25319 27108
rect 25497 27100 25543 27113
rect 25686 27188 26008 27248
rect 26054 27188 26091 27328
rect 25686 27174 26091 27188
rect 25686 27159 26001 27174
rect 25686 27113 25721 27159
rect 25767 27122 26001 27159
rect 26053 27122 26091 27174
rect 25767 27113 26091 27122
rect 25686 27108 26091 27113
rect 25721 27100 25767 27108
rect 25965 27082 26089 27108
rect 25381 27021 25637 27032
rect 25381 27015 25392 27021
rect 24210 26975 25392 27015
rect 25626 26975 25637 27021
rect 24210 26974 25637 26975
rect 24210 26922 24869 26974
rect 24921 26922 25081 26974
rect 25133 26922 25637 26974
rect 24210 26895 25637 26922
rect 22914 26842 22949 26888
rect 22995 26842 23029 26888
rect 24831 26882 25171 26895
rect 22914 26841 23029 26842
rect 22725 26678 22771 26737
rect 22725 26573 22771 26632
rect 22725 26468 22771 26527
rect 22725 26363 22771 26422
rect 22725 26258 22771 26317
rect 22725 26153 22771 26212
rect 22725 26048 22771 26107
rect 22725 25943 22771 26002
rect 22725 25838 22771 25897
rect 22725 25733 22771 25792
rect 22725 25628 22771 25687
rect 22725 25524 22771 25582
rect 22725 25420 22771 25478
rect 22725 25339 22771 25374
rect 22949 26783 22995 26841
rect 22949 26678 22995 26737
rect 23956 26733 24002 26743
rect 22949 26573 22995 26632
rect 22949 26468 22995 26527
rect 22949 26363 22995 26422
rect 22949 26258 22995 26317
rect 22949 26153 22995 26212
rect 22949 26048 22995 26107
rect 22949 25943 22995 26002
rect 22949 25838 22995 25897
rect 22949 25733 22995 25792
rect 22949 25628 22995 25687
rect 22949 25524 22995 25582
rect 22949 25420 22995 25478
rect 23605 26730 24036 26733
rect 23605 26684 23956 26730
rect 24002 26684 24036 26730
rect 23605 26636 24036 26684
rect 23605 26590 23652 26636
rect 23698 26627 24036 26636
rect 23698 26590 23956 26627
rect 23605 26581 23956 26590
rect 24002 26581 24036 26627
rect 23605 26535 24036 26581
rect 23605 26483 23739 26535
rect 23791 26483 23946 26535
rect 23998 26524 24036 26535
rect 23605 26478 23956 26483
rect 24002 26478 24036 26524
rect 23605 26473 24036 26478
rect 23605 26427 23652 26473
rect 23698 26427 24036 26473
rect 23605 26421 24036 26427
rect 23605 26375 23956 26421
rect 24002 26375 24036 26421
rect 23605 26318 24036 26375
rect 23605 26317 23956 26318
rect 23605 26309 23739 26317
rect 23605 26263 23652 26309
rect 23698 26265 23739 26309
rect 23791 26265 23946 26317
rect 24002 26272 24036 26318
rect 23998 26265 24036 26272
rect 23698 26263 24036 26265
rect 23605 26214 24036 26263
rect 23605 26168 23956 26214
rect 24002 26168 24036 26214
rect 23605 26146 24036 26168
rect 23605 26100 23652 26146
rect 23698 26110 24036 26146
rect 23698 26100 23956 26110
rect 23605 26099 23956 26100
rect 23605 26047 23739 26099
rect 23791 26047 23946 26099
rect 24002 26064 24036 26110
rect 23998 26047 24036 26064
rect 23605 26006 24036 26047
rect 23605 25983 23956 26006
rect 23605 25937 23652 25983
rect 23698 25960 23956 25983
rect 24002 25960 24036 26006
rect 23698 25937 24036 25960
rect 23605 25902 24036 25937
rect 23605 25881 23956 25902
rect 23605 25829 23739 25881
rect 23791 25829 23946 25881
rect 24002 25856 24036 25902
rect 23998 25829 24036 25856
rect 23605 25819 24036 25829
rect 23605 25773 23652 25819
rect 23698 25798 24036 25819
rect 23698 25773 23956 25798
rect 23605 25752 23956 25773
rect 24002 25752 24036 25798
rect 23605 25694 24036 25752
rect 23605 25656 23956 25694
rect 23605 25610 23652 25656
rect 23698 25648 23956 25656
rect 24002 25648 24036 25694
rect 23698 25610 24036 25648
rect 23605 25590 24036 25610
rect 23605 25544 23956 25590
rect 24002 25544 24036 25590
rect 23605 25486 24036 25544
rect 24180 26730 24226 26743
rect 24180 26627 24226 26684
rect 24180 26524 24226 26581
rect 24470 26730 24516 26743
rect 24470 26627 24516 26684
rect 24470 26575 24516 26581
rect 24694 26730 24740 26743
rect 25646 26733 25692 26743
rect 24694 26627 24740 26684
rect 24180 26421 24226 26478
rect 24180 26318 24226 26375
rect 24180 26214 24226 26272
rect 24180 26110 24226 26168
rect 24180 26006 24226 26064
rect 24180 25902 24226 25960
rect 24180 25798 24226 25856
rect 24428 26535 24556 26575
rect 24428 26483 24466 26535
rect 24518 26483 24556 26535
rect 24428 26478 24470 26483
rect 24516 26478 24556 26483
rect 24428 26421 24556 26478
rect 24428 26375 24470 26421
rect 24516 26375 24556 26421
rect 24428 26318 24556 26375
rect 24428 26317 24470 26318
rect 24516 26317 24556 26318
rect 24428 26265 24466 26317
rect 24518 26265 24556 26317
rect 24428 26214 24556 26265
rect 24428 26168 24470 26214
rect 24516 26168 24556 26214
rect 24428 26110 24556 26168
rect 24428 26099 24470 26110
rect 24516 26099 24556 26110
rect 24428 26047 24466 26099
rect 24518 26047 24556 26099
rect 24428 26006 24556 26047
rect 24428 25960 24470 26006
rect 24516 25960 24556 26006
rect 24428 25902 24556 25960
rect 24428 25881 24470 25902
rect 24516 25881 24556 25902
rect 24428 25829 24466 25881
rect 24518 25829 24556 25881
rect 24428 25798 24556 25829
rect 24428 25789 24470 25798
rect 24180 25694 24226 25752
rect 24180 25590 24226 25648
rect 24180 25496 24226 25544
rect 24516 25789 24556 25798
rect 24694 26524 24740 26581
rect 24694 26421 24740 26478
rect 24694 26318 24740 26375
rect 24694 26214 24740 26272
rect 24694 26110 24740 26168
rect 24694 26006 24740 26064
rect 24694 25902 24740 25960
rect 24694 25798 24740 25856
rect 24470 25694 24516 25752
rect 24470 25590 24516 25648
rect 23605 25440 23956 25486
rect 24002 25440 24036 25486
rect 23605 25435 24036 25440
rect 24145 25486 24260 25496
rect 24145 25440 24180 25486
rect 24226 25440 24260 25486
rect 23956 25427 24002 25435
rect 22501 25212 22547 25270
rect 22501 25108 22547 25166
rect 22501 25004 22547 25062
rect 22501 24900 22547 24958
rect 22501 24796 22547 24854
rect 22277 24692 22323 24750
rect 22277 24633 22323 24646
rect 22684 25316 22812 25339
rect 22684 25300 22725 25316
rect 22771 25300 22812 25316
rect 22684 25248 22722 25300
rect 22774 25248 22812 25300
rect 22684 25212 22812 25248
rect 22684 25166 22725 25212
rect 22771 25166 22812 25212
rect 22684 25108 22812 25166
rect 22684 25082 22725 25108
rect 22771 25082 22812 25108
rect 22684 25030 22722 25082
rect 22774 25030 22812 25082
rect 22684 25004 22812 25030
rect 22684 24958 22725 25004
rect 22771 24958 22812 25004
rect 22684 24900 22812 24958
rect 22684 24864 22725 24900
rect 22771 24864 22812 24900
rect 22684 24812 22722 24864
rect 22774 24812 22812 24864
rect 22684 24796 22812 24812
rect 22684 24772 22725 24796
rect 22501 24692 22547 24750
rect 22501 24633 22547 24646
rect 22771 24772 22812 24796
rect 22949 25316 22995 25374
rect 22949 25212 22995 25270
rect 23701 25346 24041 25353
rect 24145 25346 24260 25440
rect 24470 25486 24516 25544
rect 24694 25694 24740 25752
rect 24694 25590 24740 25648
rect 24694 25496 24740 25544
rect 25295 26730 25726 26733
rect 25295 26684 25646 26730
rect 25692 26684 25726 26730
rect 25295 26636 25726 26684
rect 25295 26590 25342 26636
rect 25388 26627 25726 26636
rect 25388 26590 25646 26627
rect 25295 26581 25646 26590
rect 25692 26581 25726 26627
rect 25295 26535 25726 26581
rect 25295 26483 25429 26535
rect 25481 26483 25636 26535
rect 25688 26524 25726 26535
rect 25295 26478 25646 26483
rect 25692 26478 25726 26524
rect 25295 26473 25726 26478
rect 25295 26427 25342 26473
rect 25388 26427 25726 26473
rect 25295 26421 25726 26427
rect 25295 26375 25646 26421
rect 25692 26375 25726 26421
rect 25295 26318 25726 26375
rect 25295 26317 25646 26318
rect 25295 26309 25429 26317
rect 25295 26263 25342 26309
rect 25388 26265 25429 26309
rect 25481 26265 25636 26317
rect 25692 26272 25726 26318
rect 25688 26265 25726 26272
rect 25388 26263 25726 26265
rect 25295 26214 25726 26263
rect 25295 26168 25646 26214
rect 25692 26168 25726 26214
rect 25295 26146 25726 26168
rect 25295 26100 25342 26146
rect 25388 26110 25726 26146
rect 25388 26100 25646 26110
rect 25295 26099 25646 26100
rect 25295 26047 25429 26099
rect 25481 26047 25636 26099
rect 25692 26064 25726 26110
rect 25688 26047 25726 26064
rect 25295 26006 25726 26047
rect 25295 25983 25646 26006
rect 25295 25937 25342 25983
rect 25388 25960 25646 25983
rect 25692 25960 25726 26006
rect 25388 25937 25726 25960
rect 25295 25902 25726 25937
rect 25295 25881 25646 25902
rect 25295 25829 25429 25881
rect 25481 25829 25636 25881
rect 25692 25856 25726 25902
rect 25688 25829 25726 25856
rect 25295 25819 25726 25829
rect 25295 25773 25342 25819
rect 25388 25798 25726 25819
rect 25388 25773 25646 25798
rect 25295 25752 25646 25773
rect 25692 25752 25726 25798
rect 25295 25694 25726 25752
rect 25295 25656 25646 25694
rect 25295 25610 25342 25656
rect 25388 25648 25646 25656
rect 25692 25648 25726 25694
rect 25388 25610 25726 25648
rect 25295 25590 25726 25610
rect 25295 25544 25646 25590
rect 25692 25544 25726 25590
rect 24470 25427 24516 25440
rect 24659 25486 24774 25496
rect 24659 25440 24694 25486
rect 24740 25440 24774 25486
rect 23701 25312 24058 25346
rect 23701 25260 23739 25312
rect 23791 25309 23951 25312
rect 24003 25309 24058 25312
rect 23791 25263 23819 25309
rect 23865 25263 23951 25309
rect 24023 25263 24058 25309
rect 23791 25260 23951 25263
rect 24003 25260 24058 25263
rect 23701 25226 24058 25260
rect 24145 25309 24568 25346
rect 24145 25263 24329 25309
rect 24375 25263 24487 25309
rect 24533 25263 24568 25309
rect 24145 25226 24568 25263
rect 23701 25220 24041 25226
rect 22949 25108 22995 25166
rect 23956 25137 24002 25147
rect 22949 25004 22995 25062
rect 22949 24900 22995 24958
rect 22949 24796 22995 24854
rect 23631 25134 24036 25137
rect 23631 25088 23956 25134
rect 24002 25088 24036 25134
rect 23631 25038 24036 25088
rect 24145 25134 24260 25226
rect 24145 25088 24180 25134
rect 24226 25088 24260 25134
rect 24145 25072 24260 25088
rect 24470 25134 24516 25147
rect 23631 25031 24049 25038
rect 23631 24985 23956 25031
rect 24002 24997 24049 25031
rect 23631 24945 23959 24985
rect 24011 24945 24049 24997
rect 23631 24928 24049 24945
rect 23631 24882 23956 24928
rect 24002 24882 24049 24928
rect 23631 24825 24049 24882
rect 23631 24802 23956 24825
rect 22725 24692 22771 24750
rect 22725 24633 22771 24646
rect 22949 24692 22995 24750
rect 22949 24633 22995 24646
rect 23556 24779 23956 24802
rect 24002 24780 24049 24825
rect 23556 24766 23959 24779
rect 23556 24720 23591 24766
rect 23637 24728 23959 24766
rect 24011 24728 24049 24780
rect 23637 24722 24049 24728
rect 23637 24720 23956 24722
rect 23556 24676 23956 24720
rect 24002 24676 24049 24722
rect 23556 24619 24049 24676
rect 23556 24602 23956 24619
rect 16670 24527 17345 24562
rect 16670 24481 16889 24527
rect 17217 24481 17345 24527
rect 16670 24443 17345 24481
rect 17453 24527 18128 24562
rect 17453 24481 17581 24527
rect 17909 24481 18128 24527
rect 17453 24443 18128 24481
rect 16670 23984 16785 24443
rect 16894 24290 17904 24326
rect 16894 24244 16981 24290
rect 17027 24244 17139 24290
rect 17185 24244 17297 24290
rect 17343 24244 17455 24290
rect 17501 24244 17613 24290
rect 17659 24244 17771 24290
rect 17817 24244 17904 24290
rect 16894 24219 17904 24244
rect 16670 23892 16704 23984
rect 15899 23370 15945 23427
rect 15899 23267 15945 23324
rect 15675 23164 15721 23195
rect 15675 23061 15721 23118
rect 15675 22958 15721 23015
rect 15675 22855 15721 22912
rect 15675 22752 15721 22809
rect 15899 23164 15945 23221
rect 15899 23061 15945 23118
rect 15899 22958 15945 23015
rect 15899 22855 15945 22912
rect 15899 22752 15945 22809
rect 15675 22649 15721 22706
rect 15675 22546 15721 22603
rect 15675 22443 15721 22500
rect 15675 22384 15721 22397
rect 15859 22706 15899 22743
rect 15945 22706 15983 22743
rect 15859 22703 15983 22706
rect 15859 22651 15895 22703
rect 15947 22651 15983 22703
rect 15859 22649 15983 22651
rect 15859 22603 15899 22649
rect 15945 22603 15983 22649
rect 15859 22546 15983 22603
rect 15859 22500 15899 22546
rect 15945 22500 15983 22546
rect 15859 22485 15983 22500
rect 15859 22433 15895 22485
rect 15947 22433 15983 22485
rect 15859 22397 15899 22433
rect 15945 22397 15983 22433
rect 15859 22393 15983 22397
rect 15899 22384 15945 22393
rect 16665 22230 16704 22270
rect 16750 23892 16785 23984
rect 16891 24207 17907 24219
rect 16891 24180 17019 24207
rect 16891 24128 16929 24180
rect 16981 24128 17019 24180
rect 16891 23984 17019 24128
rect 17335 24180 17463 24207
rect 17335 24128 17373 24180
rect 17425 24128 17463 24180
rect 16891 22781 16928 23984
rect 16974 23962 17019 23984
rect 16981 23910 17019 23962
rect 16974 23745 17019 23910
rect 16981 23693 17019 23745
rect 16974 23527 17019 23693
rect 16981 23475 17019 23527
rect 16974 23309 17019 23475
rect 16981 23257 17019 23309
rect 16974 23092 17019 23257
rect 16981 23040 17019 23092
rect 16974 22874 17019 23040
rect 16981 22822 17019 22874
rect 16750 22230 16789 22270
rect 16665 22178 16701 22230
rect 16753 22178 16789 22230
rect 16665 22012 16704 22178
rect 16750 22012 16789 22178
rect 16665 21960 16701 22012
rect 16753 21960 16789 22012
rect 16665 21924 16704 21960
rect 16750 21924 16789 21960
rect 16665 21920 16789 21924
rect 16974 22782 17019 22822
rect 17152 23984 17198 23997
rect 16974 22781 17006 22782
rect 16704 21911 16750 21920
rect 16928 21911 16974 21924
rect 17113 22230 17152 22270
rect 17335 23984 17463 24128
rect 17779 24180 17907 24207
rect 17779 24128 17817 24180
rect 17869 24128 17907 24180
rect 17335 23962 17376 23984
rect 17422 23962 17463 23984
rect 17335 23910 17373 23962
rect 17425 23910 17463 23962
rect 17335 23745 17376 23910
rect 17422 23745 17463 23910
rect 17335 23693 17373 23745
rect 17425 23693 17463 23745
rect 17335 23527 17376 23693
rect 17422 23527 17463 23693
rect 17335 23475 17373 23527
rect 17425 23475 17463 23527
rect 17335 23309 17376 23475
rect 17422 23309 17463 23475
rect 17335 23257 17373 23309
rect 17425 23257 17463 23309
rect 17335 23092 17376 23257
rect 17422 23092 17463 23257
rect 17335 23040 17373 23092
rect 17425 23040 17463 23092
rect 17335 22874 17376 23040
rect 17422 22874 17463 23040
rect 17335 22822 17373 22874
rect 17425 22822 17463 22874
rect 17335 22781 17376 22822
rect 17198 22230 17237 22270
rect 17113 22178 17149 22230
rect 17201 22178 17237 22230
rect 17113 22012 17152 22178
rect 17198 22012 17237 22178
rect 17113 21960 17149 22012
rect 17201 21960 17237 22012
rect 17113 21924 17152 21960
rect 17198 21924 17237 21960
rect 17113 21920 17237 21924
rect 17422 22781 17463 22822
rect 17600 23984 17646 23997
rect 17152 21911 17198 21920
rect 17376 21911 17422 21924
rect 17561 22230 17600 22270
rect 17779 23984 17907 24128
rect 17779 23962 17824 23984
rect 17779 23910 17817 23962
rect 17779 23745 17824 23910
rect 17779 23693 17817 23745
rect 17779 23527 17824 23693
rect 17779 23475 17817 23527
rect 17779 23309 17824 23475
rect 17779 23257 17817 23309
rect 17779 23092 17824 23257
rect 17779 23040 17817 23092
rect 17779 22874 17824 23040
rect 17779 22822 17817 22874
rect 17779 22782 17824 22822
rect 17792 22781 17824 22782
rect 17646 22230 17685 22270
rect 17561 22178 17597 22230
rect 17649 22178 17685 22230
rect 17561 22012 17600 22178
rect 17646 22012 17685 22178
rect 17561 21960 17597 22012
rect 17649 21960 17685 22012
rect 17561 21924 17600 21960
rect 17646 21924 17685 21960
rect 17561 21920 17685 21924
rect 17870 22781 17907 23984
rect 18013 23984 18128 24443
rect 18013 23892 18048 23984
rect 17600 21911 17646 21920
rect 17824 21911 17870 21924
rect 18009 22230 18048 22270
rect 18094 23892 18128 23984
rect 18304 24527 18979 24562
rect 18304 24481 18523 24527
rect 18851 24481 18979 24527
rect 18304 24443 18979 24481
rect 19087 24527 19762 24562
rect 19087 24481 19215 24527
rect 19543 24481 19762 24527
rect 19087 24443 19762 24481
rect 18304 23984 18419 24443
rect 18528 24290 19538 24326
rect 18528 24244 18615 24290
rect 18661 24244 18773 24290
rect 18819 24244 18931 24290
rect 18977 24244 19089 24290
rect 19135 24244 19247 24290
rect 19293 24244 19405 24290
rect 19451 24244 19538 24290
rect 18528 24219 19538 24244
rect 18304 23892 18338 23984
rect 18094 22230 18133 22270
rect 18009 22178 18045 22230
rect 18097 22178 18133 22230
rect 18009 22012 18048 22178
rect 18094 22012 18133 22178
rect 18009 21960 18045 22012
rect 18097 21960 18133 22012
rect 18009 21924 18048 21960
rect 18094 21924 18133 21960
rect 18009 21920 18133 21924
rect 18299 22230 18338 22270
rect 18384 23892 18419 23984
rect 18525 24207 19541 24219
rect 18525 24180 18653 24207
rect 18525 24128 18563 24180
rect 18615 24128 18653 24180
rect 18525 23984 18653 24128
rect 18969 24180 19097 24207
rect 18969 24128 19007 24180
rect 19059 24128 19097 24180
rect 18525 22781 18562 23984
rect 18608 23962 18653 23984
rect 18615 23910 18653 23962
rect 18608 23745 18653 23910
rect 18615 23693 18653 23745
rect 18608 23527 18653 23693
rect 18615 23475 18653 23527
rect 18608 23309 18653 23475
rect 18615 23257 18653 23309
rect 18608 23092 18653 23257
rect 18615 23040 18653 23092
rect 18608 22874 18653 23040
rect 18615 22822 18653 22874
rect 18384 22230 18423 22270
rect 18299 22178 18335 22230
rect 18387 22178 18423 22230
rect 18299 22012 18338 22178
rect 18384 22012 18423 22178
rect 18299 21960 18335 22012
rect 18387 21960 18423 22012
rect 18299 21924 18338 21960
rect 18384 21924 18423 21960
rect 18299 21920 18423 21924
rect 18608 22782 18653 22822
rect 18786 23984 18832 23997
rect 18608 22781 18640 22782
rect 18048 21911 18094 21920
rect 18338 21911 18384 21920
rect 18562 21911 18608 21924
rect 18747 22230 18786 22270
rect 18969 23984 19097 24128
rect 19413 24180 19541 24207
rect 19413 24128 19451 24180
rect 19503 24128 19541 24180
rect 18969 23962 19010 23984
rect 19056 23962 19097 23984
rect 18969 23910 19007 23962
rect 19059 23910 19097 23962
rect 18969 23745 19010 23910
rect 19056 23745 19097 23910
rect 18969 23693 19007 23745
rect 19059 23693 19097 23745
rect 18969 23527 19010 23693
rect 19056 23527 19097 23693
rect 18969 23475 19007 23527
rect 19059 23475 19097 23527
rect 18969 23309 19010 23475
rect 19056 23309 19097 23475
rect 18969 23257 19007 23309
rect 19059 23257 19097 23309
rect 18969 23092 19010 23257
rect 19056 23092 19097 23257
rect 18969 23040 19007 23092
rect 19059 23040 19097 23092
rect 18969 22874 19010 23040
rect 19056 22874 19097 23040
rect 18969 22822 19007 22874
rect 19059 22822 19097 22874
rect 18969 22781 19010 22822
rect 18832 22230 18871 22270
rect 18747 22178 18783 22230
rect 18835 22178 18871 22230
rect 18747 22012 18786 22178
rect 18832 22012 18871 22178
rect 18747 21960 18783 22012
rect 18835 21960 18871 22012
rect 18747 21924 18786 21960
rect 18832 21924 18871 21960
rect 18747 21920 18871 21924
rect 19056 22781 19097 22822
rect 19234 23984 19280 23997
rect 18786 21911 18832 21920
rect 19010 21911 19056 21924
rect 19195 22230 19234 22270
rect 19413 23984 19541 24128
rect 19413 23962 19458 23984
rect 19413 23910 19451 23962
rect 19413 23745 19458 23910
rect 19413 23693 19451 23745
rect 19413 23527 19458 23693
rect 19413 23475 19451 23527
rect 19413 23309 19458 23475
rect 19413 23257 19451 23309
rect 19413 23092 19458 23257
rect 19413 23040 19451 23092
rect 19413 22874 19458 23040
rect 19413 22822 19451 22874
rect 19413 22782 19458 22822
rect 19426 22781 19458 22782
rect 19280 22230 19319 22270
rect 19195 22178 19231 22230
rect 19283 22178 19319 22230
rect 19195 22012 19234 22178
rect 19280 22012 19319 22178
rect 19195 21960 19231 22012
rect 19283 21960 19319 22012
rect 19195 21924 19234 21960
rect 19280 21924 19319 21960
rect 19195 21920 19319 21924
rect 19504 22781 19541 23984
rect 19647 23984 19762 24443
rect 19647 23892 19682 23984
rect 19234 21911 19280 21920
rect 19458 21911 19504 21924
rect 19643 22230 19682 22270
rect 19728 23892 19762 23984
rect 19937 24527 20612 24562
rect 19937 24481 20156 24527
rect 20484 24481 20612 24527
rect 19937 24443 20612 24481
rect 20720 24527 21395 24562
rect 20720 24481 20848 24527
rect 21176 24481 21395 24527
rect 20720 24443 21395 24481
rect 19937 23984 20052 24443
rect 20161 24290 21171 24326
rect 20161 24244 20248 24290
rect 20294 24244 20406 24290
rect 20452 24244 20564 24290
rect 20610 24244 20722 24290
rect 20768 24244 20880 24290
rect 20926 24244 21038 24290
rect 21084 24244 21171 24290
rect 20161 24219 21171 24244
rect 19937 23892 19971 23984
rect 19728 22230 19767 22270
rect 19643 22178 19679 22230
rect 19731 22178 19767 22230
rect 19643 22012 19682 22178
rect 19728 22012 19767 22178
rect 19643 21960 19679 22012
rect 19731 21960 19767 22012
rect 19643 21924 19682 21960
rect 19728 21924 19767 21960
rect 19643 21920 19767 21924
rect 19932 22230 19971 22270
rect 20017 23892 20052 23984
rect 20158 24207 21174 24219
rect 20158 24180 20286 24207
rect 20158 24128 20196 24180
rect 20248 24128 20286 24180
rect 20158 23984 20286 24128
rect 20602 24180 20730 24207
rect 20602 24128 20640 24180
rect 20692 24128 20730 24180
rect 20158 22781 20195 23984
rect 20241 23962 20286 23984
rect 20248 23910 20286 23962
rect 20241 23745 20286 23910
rect 20248 23693 20286 23745
rect 20241 23527 20286 23693
rect 20248 23475 20286 23527
rect 20241 23309 20286 23475
rect 20248 23257 20286 23309
rect 20241 23092 20286 23257
rect 20248 23040 20286 23092
rect 20241 22874 20286 23040
rect 20248 22822 20286 22874
rect 20017 22230 20056 22270
rect 19932 22178 19968 22230
rect 20020 22178 20056 22230
rect 19932 22012 19971 22178
rect 20017 22012 20056 22178
rect 19932 21960 19968 22012
rect 20020 21960 20056 22012
rect 19932 21924 19971 21960
rect 20017 21924 20056 21960
rect 19932 21920 20056 21924
rect 20241 22782 20286 22822
rect 20419 23984 20465 23997
rect 20241 22781 20273 22782
rect 19682 21911 19728 21920
rect 19971 21911 20017 21920
rect 20195 21911 20241 21924
rect 20380 22230 20419 22270
rect 20602 23984 20730 24128
rect 21046 24180 21174 24207
rect 21046 24128 21084 24180
rect 21136 24128 21174 24180
rect 20602 23962 20643 23984
rect 20689 23962 20730 23984
rect 20602 23910 20640 23962
rect 20692 23910 20730 23962
rect 20602 23745 20643 23910
rect 20689 23745 20730 23910
rect 20602 23693 20640 23745
rect 20692 23693 20730 23745
rect 20602 23527 20643 23693
rect 20689 23527 20730 23693
rect 20602 23475 20640 23527
rect 20692 23475 20730 23527
rect 20602 23309 20643 23475
rect 20689 23309 20730 23475
rect 20602 23257 20640 23309
rect 20692 23257 20730 23309
rect 20602 23092 20643 23257
rect 20689 23092 20730 23257
rect 20602 23040 20640 23092
rect 20692 23040 20730 23092
rect 20602 22874 20643 23040
rect 20689 22874 20730 23040
rect 20602 22822 20640 22874
rect 20692 22822 20730 22874
rect 20602 22781 20643 22822
rect 20465 22230 20504 22270
rect 20380 22178 20416 22230
rect 20468 22178 20504 22230
rect 20380 22012 20419 22178
rect 20465 22012 20504 22178
rect 20380 21960 20416 22012
rect 20468 21960 20504 22012
rect 20380 21924 20419 21960
rect 20465 21924 20504 21960
rect 20380 21920 20504 21924
rect 20689 22781 20730 22822
rect 20867 23984 20913 23997
rect 20419 21911 20465 21920
rect 20643 21911 20689 21924
rect 20828 22230 20867 22270
rect 21046 23984 21174 24128
rect 21046 23962 21091 23984
rect 21046 23910 21084 23962
rect 21046 23745 21091 23910
rect 21046 23693 21084 23745
rect 21046 23527 21091 23693
rect 21046 23475 21084 23527
rect 21046 23309 21091 23475
rect 21046 23257 21084 23309
rect 21046 23092 21091 23257
rect 21046 23040 21084 23092
rect 21046 22874 21091 23040
rect 21046 22822 21084 22874
rect 21046 22782 21091 22822
rect 21059 22781 21091 22782
rect 20913 22230 20952 22270
rect 20828 22178 20864 22230
rect 20916 22178 20952 22230
rect 20828 22012 20867 22178
rect 20913 22012 20952 22178
rect 20828 21960 20864 22012
rect 20916 21960 20952 22012
rect 20828 21924 20867 21960
rect 20913 21924 20952 21960
rect 20828 21920 20952 21924
rect 21137 22781 21174 23984
rect 21280 23984 21395 24443
rect 21280 23892 21315 23984
rect 20867 21911 20913 21920
rect 21091 21911 21137 21924
rect 21276 22230 21315 22270
rect 21361 23892 21395 23984
rect 21571 24527 22246 24562
rect 21571 24481 21790 24527
rect 22118 24481 22246 24527
rect 21571 24443 22246 24481
rect 22354 24527 23029 24562
rect 22354 24481 22482 24527
rect 22810 24481 23029 24527
rect 22354 24443 23029 24481
rect 21571 23984 21686 24443
rect 21795 24290 22805 24326
rect 21795 24244 21882 24290
rect 21928 24244 22040 24290
rect 22086 24244 22198 24290
rect 22244 24244 22356 24290
rect 22402 24244 22514 24290
rect 22560 24244 22672 24290
rect 22718 24244 22805 24290
rect 21795 24219 22805 24244
rect 21571 23892 21605 23984
rect 21361 22230 21400 22270
rect 21276 22178 21312 22230
rect 21364 22178 21400 22230
rect 21276 22012 21315 22178
rect 21361 22012 21400 22178
rect 21276 21960 21312 22012
rect 21364 21960 21400 22012
rect 21276 21924 21315 21960
rect 21361 21924 21400 21960
rect 21276 21920 21400 21924
rect 21566 22230 21605 22270
rect 21651 23892 21686 23984
rect 21792 24207 22808 24219
rect 21792 24180 21920 24207
rect 21792 24128 21830 24180
rect 21882 24128 21920 24180
rect 21792 23984 21920 24128
rect 22236 24180 22364 24207
rect 22236 24128 22274 24180
rect 22326 24128 22364 24180
rect 21792 22781 21829 23984
rect 21875 23962 21920 23984
rect 21882 23910 21920 23962
rect 21875 23745 21920 23910
rect 21882 23693 21920 23745
rect 21875 23527 21920 23693
rect 21882 23475 21920 23527
rect 21875 23309 21920 23475
rect 21882 23257 21920 23309
rect 21875 23092 21920 23257
rect 21882 23040 21920 23092
rect 21875 22874 21920 23040
rect 21882 22822 21920 22874
rect 21651 22230 21690 22270
rect 21566 22178 21602 22230
rect 21654 22178 21690 22230
rect 21566 22012 21605 22178
rect 21651 22012 21690 22178
rect 21566 21960 21602 22012
rect 21654 21960 21690 22012
rect 21566 21924 21605 21960
rect 21651 21924 21690 21960
rect 21566 21920 21690 21924
rect 21875 22782 21920 22822
rect 22053 23984 22099 23997
rect 21875 22781 21907 22782
rect 21315 21911 21361 21920
rect 21605 21911 21651 21920
rect 21829 21911 21875 21924
rect 22014 22230 22053 22270
rect 22236 23984 22364 24128
rect 22680 24180 22808 24207
rect 22680 24128 22718 24180
rect 22770 24128 22808 24180
rect 22236 23962 22277 23984
rect 22323 23962 22364 23984
rect 22236 23910 22274 23962
rect 22326 23910 22364 23962
rect 22236 23745 22277 23910
rect 22323 23745 22364 23910
rect 22236 23693 22274 23745
rect 22326 23693 22364 23745
rect 22236 23527 22277 23693
rect 22323 23527 22364 23693
rect 22236 23475 22274 23527
rect 22326 23475 22364 23527
rect 22236 23309 22277 23475
rect 22323 23309 22364 23475
rect 22236 23257 22274 23309
rect 22326 23257 22364 23309
rect 22236 23092 22277 23257
rect 22323 23092 22364 23257
rect 22236 23040 22274 23092
rect 22326 23040 22364 23092
rect 22236 22874 22277 23040
rect 22323 22874 22364 23040
rect 22236 22822 22274 22874
rect 22326 22822 22364 22874
rect 22236 22781 22277 22822
rect 22099 22230 22138 22270
rect 22014 22178 22050 22230
rect 22102 22178 22138 22230
rect 22014 22012 22053 22178
rect 22099 22012 22138 22178
rect 22014 21960 22050 22012
rect 22102 21960 22138 22012
rect 22014 21924 22053 21960
rect 22099 21924 22138 21960
rect 22014 21920 22138 21924
rect 22323 22781 22364 22822
rect 22501 23984 22547 23997
rect 22053 21911 22099 21920
rect 22277 21911 22323 21924
rect 22462 22230 22501 22270
rect 22680 23984 22808 24128
rect 22680 23962 22725 23984
rect 22680 23910 22718 23962
rect 22680 23745 22725 23910
rect 22680 23693 22718 23745
rect 22680 23527 22725 23693
rect 22680 23475 22718 23527
rect 22680 23309 22725 23475
rect 22680 23257 22718 23309
rect 22680 23092 22725 23257
rect 22680 23040 22718 23092
rect 22680 22874 22725 23040
rect 22680 22822 22718 22874
rect 22680 22782 22725 22822
rect 22693 22781 22725 22782
rect 22547 22230 22586 22270
rect 22462 22178 22498 22230
rect 22550 22178 22586 22230
rect 22462 22012 22501 22178
rect 22547 22012 22586 22178
rect 22462 21960 22498 22012
rect 22550 21960 22586 22012
rect 22462 21924 22501 21960
rect 22547 21924 22586 21960
rect 22462 21920 22586 21924
rect 22771 22781 22808 23984
rect 22914 23984 23029 24443
rect 22914 23892 22949 23984
rect 22501 21911 22547 21920
rect 22725 21911 22771 21924
rect 22910 22230 22949 22270
rect 22995 23892 23029 23984
rect 23556 24556 23591 24602
rect 23637 24573 23956 24602
rect 24002 24573 24049 24619
rect 23637 24562 24049 24573
rect 23637 24556 23959 24562
rect 23556 24516 23959 24556
rect 23556 24470 23956 24516
rect 24011 24510 24049 24562
rect 24002 24470 24049 24510
rect 23556 24439 24049 24470
rect 23556 24393 23591 24439
rect 23637 24413 24049 24439
rect 23637 24393 23956 24413
rect 23556 24367 23956 24393
rect 24002 24367 24049 24413
rect 23556 24344 24049 24367
rect 23556 24310 23959 24344
rect 23556 24276 23956 24310
rect 24011 24292 24049 24344
rect 23556 24230 23591 24276
rect 23637 24264 23956 24276
rect 24002 24264 24049 24292
rect 23637 24230 24049 24264
rect 23556 24207 24049 24230
rect 23556 24161 23956 24207
rect 24002 24161 24049 24207
rect 23556 24126 24049 24161
rect 23556 24113 23959 24126
rect 23556 24067 23591 24113
rect 23637 24104 23959 24113
rect 23637 24067 23956 24104
rect 24011 24074 24049 24126
rect 23556 24058 23956 24067
rect 24002 24058 24049 24074
rect 23556 24001 24049 24058
rect 23556 23955 23956 24001
rect 24002 23955 24049 24001
rect 23556 23950 24049 23955
rect 23556 23904 23591 23950
rect 23637 23909 24049 23950
rect 23637 23904 23959 23909
rect 23556 23898 23959 23904
rect 23556 23852 23956 23898
rect 24011 23857 24049 23909
rect 24002 23852 24049 23857
rect 23556 23817 24049 23852
rect 24180 25031 24226 25072
rect 24470 25038 24516 25088
rect 24659 25134 24774 25440
rect 25295 25486 25726 25544
rect 25870 26730 25916 26743
rect 25870 26627 25916 26684
rect 25870 26524 25916 26581
rect 26160 26730 26206 26743
rect 26160 26627 26206 26684
rect 26160 26575 26206 26581
rect 26384 26730 26430 26743
rect 27337 26733 27383 26743
rect 26384 26627 26430 26684
rect 25870 26421 25916 26478
rect 25870 26318 25916 26375
rect 25870 26214 25916 26272
rect 25870 26110 25916 26168
rect 25870 26006 25916 26064
rect 25870 25902 25916 25960
rect 25870 25798 25916 25856
rect 26118 26535 26246 26575
rect 26118 26483 26156 26535
rect 26208 26483 26246 26535
rect 26118 26478 26160 26483
rect 26206 26478 26246 26483
rect 26118 26421 26246 26478
rect 26118 26375 26160 26421
rect 26206 26375 26246 26421
rect 26118 26318 26246 26375
rect 26118 26317 26160 26318
rect 26206 26317 26246 26318
rect 26118 26265 26156 26317
rect 26208 26265 26246 26317
rect 26118 26214 26246 26265
rect 26118 26168 26160 26214
rect 26206 26168 26246 26214
rect 26118 26110 26246 26168
rect 26118 26099 26160 26110
rect 26206 26099 26246 26110
rect 26118 26047 26156 26099
rect 26208 26047 26246 26099
rect 26118 26006 26246 26047
rect 26118 25960 26160 26006
rect 26206 25960 26246 26006
rect 26118 25902 26246 25960
rect 26118 25881 26160 25902
rect 26206 25881 26246 25902
rect 26118 25829 26156 25881
rect 26208 25829 26246 25881
rect 26118 25798 26246 25829
rect 26118 25789 26160 25798
rect 25870 25694 25916 25752
rect 25870 25590 25916 25648
rect 25870 25496 25916 25544
rect 26206 25789 26246 25798
rect 26384 26524 26430 26581
rect 26384 26421 26430 26478
rect 26384 26318 26430 26375
rect 26384 26214 26430 26272
rect 26384 26110 26430 26168
rect 26384 26006 26430 26064
rect 26384 25902 26430 25960
rect 26384 25798 26430 25856
rect 26160 25694 26206 25752
rect 26160 25590 26206 25648
rect 25295 25440 25646 25486
rect 25692 25440 25726 25486
rect 25295 25435 25726 25440
rect 25835 25486 25950 25496
rect 25835 25440 25870 25486
rect 25916 25440 25950 25486
rect 25646 25427 25692 25435
rect 25391 25346 25731 25353
rect 25835 25346 25950 25440
rect 26160 25486 26206 25544
rect 26384 25694 26430 25752
rect 26384 25590 26430 25648
rect 26384 25496 26430 25544
rect 26986 26730 27417 26733
rect 26986 26684 27337 26730
rect 27383 26684 27417 26730
rect 26986 26636 27417 26684
rect 26986 26590 27033 26636
rect 27079 26627 27417 26636
rect 27079 26590 27337 26627
rect 26986 26581 27337 26590
rect 27383 26581 27417 26627
rect 26986 26535 27417 26581
rect 26986 26483 27120 26535
rect 27172 26483 27327 26535
rect 27379 26524 27417 26535
rect 26986 26478 27337 26483
rect 27383 26478 27417 26524
rect 26986 26473 27417 26478
rect 26986 26427 27033 26473
rect 27079 26427 27417 26473
rect 26986 26421 27417 26427
rect 26986 26375 27337 26421
rect 27383 26375 27417 26421
rect 26986 26318 27417 26375
rect 26986 26317 27337 26318
rect 26986 26309 27120 26317
rect 26986 26263 27033 26309
rect 27079 26265 27120 26309
rect 27172 26265 27327 26317
rect 27383 26272 27417 26318
rect 27379 26265 27417 26272
rect 27079 26263 27417 26265
rect 26986 26214 27417 26263
rect 26986 26168 27337 26214
rect 27383 26168 27417 26214
rect 26986 26146 27417 26168
rect 26986 26100 27033 26146
rect 27079 26110 27417 26146
rect 27079 26100 27337 26110
rect 26986 26099 27337 26100
rect 26986 26047 27120 26099
rect 27172 26047 27327 26099
rect 27383 26064 27417 26110
rect 27379 26047 27417 26064
rect 26986 26006 27417 26047
rect 26986 25983 27337 26006
rect 26986 25937 27033 25983
rect 27079 25960 27337 25983
rect 27383 25960 27417 26006
rect 27079 25937 27417 25960
rect 26986 25902 27417 25937
rect 26986 25881 27337 25902
rect 26986 25829 27120 25881
rect 27172 25829 27327 25881
rect 27383 25856 27417 25902
rect 27379 25829 27417 25856
rect 26986 25819 27417 25829
rect 26986 25773 27033 25819
rect 27079 25798 27417 25819
rect 27079 25773 27337 25798
rect 26986 25752 27337 25773
rect 27383 25752 27417 25798
rect 26986 25694 27417 25752
rect 26986 25656 27337 25694
rect 26986 25610 27033 25656
rect 27079 25648 27337 25656
rect 27383 25648 27417 25694
rect 27079 25610 27417 25648
rect 26986 25590 27417 25610
rect 26986 25544 27337 25590
rect 27383 25544 27417 25590
rect 26160 25427 26206 25440
rect 26349 25486 26464 25496
rect 26349 25440 26384 25486
rect 26430 25440 26464 25486
rect 25391 25312 25748 25346
rect 25391 25260 25429 25312
rect 25481 25309 25641 25312
rect 25693 25309 25748 25312
rect 25481 25263 25509 25309
rect 25555 25263 25641 25309
rect 25713 25263 25748 25309
rect 25481 25260 25641 25263
rect 25693 25260 25748 25263
rect 25391 25226 25748 25260
rect 25835 25309 26258 25346
rect 25835 25263 26019 25309
rect 26065 25263 26177 25309
rect 26223 25263 26258 25309
rect 25835 25226 26258 25263
rect 25391 25220 25731 25226
rect 25646 25137 25692 25147
rect 24659 25088 24694 25134
rect 24740 25088 24774 25134
rect 24659 25072 24774 25088
rect 25321 25134 25726 25137
rect 25321 25088 25646 25134
rect 25692 25088 25726 25134
rect 24180 24928 24226 24985
rect 24180 24825 24226 24882
rect 24180 24722 24226 24779
rect 24180 24619 24226 24676
rect 24180 24516 24226 24573
rect 24180 24413 24226 24470
rect 24180 24310 24226 24367
rect 24180 24207 24226 24264
rect 24180 24104 24226 24161
rect 24180 24001 24226 24058
rect 24180 23898 24226 23955
rect 23556 23816 24043 23817
rect 23556 23795 24036 23816
rect 23556 23786 23956 23795
rect 23556 23740 23591 23786
rect 23637 23749 23956 23786
rect 24002 23749 24036 23795
rect 23637 23740 24036 23749
rect 23556 23692 24036 23740
rect 23556 23646 23956 23692
rect 24002 23646 24036 23692
rect 23556 23623 24036 23646
rect 23556 23577 23591 23623
rect 23637 23589 24036 23623
rect 23637 23577 23956 23589
rect 23556 23543 23956 23577
rect 24002 23543 24036 23589
rect 23556 23486 24036 23543
rect 23556 23460 23956 23486
rect 23556 23414 23591 23460
rect 23637 23440 23956 23460
rect 24002 23440 24036 23486
rect 23637 23414 24036 23440
rect 23556 23383 24036 23414
rect 23556 23337 23956 23383
rect 24002 23337 24036 23383
rect 23556 23296 24036 23337
rect 23556 23250 23591 23296
rect 23637 23280 24036 23296
rect 23637 23250 23956 23280
rect 23556 23234 23956 23250
rect 24002 23234 24036 23280
rect 23556 23177 24036 23234
rect 23556 23133 23956 23177
rect 23556 23087 23591 23133
rect 23637 23131 23956 23133
rect 24002 23131 24036 23177
rect 23637 23087 24036 23131
rect 23556 23074 24036 23087
rect 23556 23028 23956 23074
rect 24002 23028 24036 23074
rect 23556 22971 24036 23028
rect 23556 22970 23956 22971
rect 23556 22924 23591 22970
rect 23637 22925 23956 22970
rect 24002 22925 24036 22971
rect 23637 22924 24036 22925
rect 23556 22868 24036 22924
rect 23556 22822 23956 22868
rect 24002 22822 24036 22868
rect 23556 22806 24036 22822
rect 23556 22760 23591 22806
rect 23637 22765 24036 22806
rect 23637 22760 23956 22765
rect 23556 22719 23956 22760
rect 24002 22719 24036 22765
rect 23556 22662 24036 22719
rect 23556 22643 23956 22662
rect 23556 22597 23591 22643
rect 23637 22616 23956 22643
rect 24002 22616 24036 22662
rect 23637 22597 24036 22616
rect 23556 22559 24036 22597
rect 23556 22513 23956 22559
rect 24002 22513 24036 22559
rect 23556 22480 24036 22513
rect 23556 22434 23591 22480
rect 23637 22456 24036 22480
rect 23637 22434 23956 22456
rect 23556 22410 23956 22434
rect 24002 22410 24036 22456
rect 23556 22353 24036 22410
rect 23556 22317 23956 22353
rect 23556 22271 23591 22317
rect 23637 22307 23956 22317
rect 24002 22307 24036 22353
rect 23637 22271 24036 22307
rect 22995 22230 23034 22270
rect 22910 22178 22946 22230
rect 22998 22178 23034 22230
rect 22910 22012 22949 22178
rect 22995 22012 23034 22178
rect 22910 21960 22946 22012
rect 22998 21960 23034 22012
rect 22910 21924 22949 21960
rect 22995 21924 23034 21960
rect 22910 21920 23034 21924
rect 23556 22250 24036 22271
rect 23556 22204 23956 22250
rect 24002 22204 24036 22250
rect 24180 23795 24226 23852
rect 24435 25031 24563 25038
rect 24435 24985 24470 25031
rect 24516 24997 24563 25031
rect 24435 24945 24473 24985
rect 24525 24945 24563 24997
rect 24435 24928 24563 24945
rect 24435 24882 24470 24928
rect 24516 24882 24563 24928
rect 24435 24825 24563 24882
rect 24435 24779 24470 24825
rect 24516 24780 24563 24825
rect 24435 24728 24473 24779
rect 24525 24728 24563 24780
rect 24435 24722 24563 24728
rect 24435 24676 24470 24722
rect 24516 24676 24563 24722
rect 24435 24619 24563 24676
rect 24435 24573 24470 24619
rect 24516 24573 24563 24619
rect 24435 24562 24563 24573
rect 24435 24516 24473 24562
rect 24435 24470 24470 24516
rect 24525 24510 24563 24562
rect 24516 24470 24563 24510
rect 24435 24413 24563 24470
rect 24435 24367 24470 24413
rect 24516 24367 24563 24413
rect 24435 24344 24563 24367
rect 24435 24310 24473 24344
rect 24435 24264 24470 24310
rect 24525 24292 24563 24344
rect 24516 24264 24563 24292
rect 24435 24207 24563 24264
rect 24435 24161 24470 24207
rect 24516 24161 24563 24207
rect 24435 24126 24563 24161
rect 24435 24104 24473 24126
rect 24435 24058 24470 24104
rect 24525 24074 24563 24126
rect 24516 24058 24563 24074
rect 24435 24001 24563 24058
rect 24435 23955 24470 24001
rect 24516 23955 24563 24001
rect 24435 23909 24563 23955
rect 24435 23898 24473 23909
rect 24435 23852 24470 23898
rect 24525 23857 24563 23909
rect 24516 23852 24563 23857
rect 24435 23817 24563 23852
rect 24694 25031 24740 25072
rect 24694 24928 24740 24985
rect 24694 24825 24740 24882
rect 25321 25038 25726 25088
rect 25835 25134 25950 25226
rect 25835 25088 25870 25134
rect 25916 25088 25950 25134
rect 25835 25072 25950 25088
rect 26160 25134 26206 25147
rect 25321 25031 25739 25038
rect 25321 24985 25646 25031
rect 25692 24997 25739 25031
rect 25321 24945 25649 24985
rect 25701 24945 25739 24997
rect 25321 24928 25739 24945
rect 25321 24882 25646 24928
rect 25692 24882 25739 24928
rect 25321 24825 25739 24882
rect 25321 24802 25646 24825
rect 24694 24722 24740 24779
rect 24694 24619 24740 24676
rect 24694 24516 24740 24573
rect 24694 24413 24740 24470
rect 24694 24310 24740 24367
rect 24694 24207 24740 24264
rect 24694 24104 24740 24161
rect 24694 24001 24740 24058
rect 24694 23898 24740 23955
rect 24441 23816 24557 23817
rect 24180 23692 24226 23749
rect 24180 23589 24226 23646
rect 24180 23486 24226 23543
rect 24180 23383 24226 23440
rect 24180 23280 24226 23337
rect 24180 23177 24226 23234
rect 24180 23074 24226 23131
rect 24180 22971 24226 23028
rect 24180 22868 24226 22925
rect 24180 22765 24226 22822
rect 24180 22662 24226 22719
rect 24180 22559 24226 22616
rect 24180 22456 24226 22513
rect 24180 22353 24226 22410
rect 24180 22250 24226 22307
rect 24144 22240 24180 22241
rect 23556 22154 24036 22204
rect 23556 22108 23591 22154
rect 23637 22147 24036 22154
rect 23637 22108 23956 22147
rect 23556 22101 23956 22108
rect 24002 22101 24036 22147
rect 23556 22044 24036 22101
rect 23556 21998 23956 22044
rect 24002 21998 24036 22044
rect 23556 21990 24036 21998
rect 23556 21944 23591 21990
rect 23637 21944 24036 21990
rect 23556 21940 24036 21944
rect 22949 21911 22995 21920
rect 23556 21908 23956 21940
rect 23630 21907 23956 21908
rect 23631 21894 23956 21907
rect 24002 21894 24036 21940
rect 23631 21889 24036 21894
rect 24137 22204 24180 22240
rect 24470 23795 24516 23816
rect 24470 23692 24516 23749
rect 24470 23589 24516 23646
rect 24470 23486 24516 23543
rect 24470 23383 24516 23440
rect 24470 23280 24516 23337
rect 24470 23177 24516 23234
rect 24470 23074 24516 23131
rect 24470 22971 24516 23028
rect 24470 22868 24516 22925
rect 24470 22765 24516 22822
rect 24470 22662 24516 22719
rect 24470 22559 24516 22616
rect 24470 22456 24516 22513
rect 24470 22353 24516 22410
rect 24470 22250 24516 22307
rect 24226 22240 24260 22241
rect 24226 22204 24267 22240
rect 24137 22200 24267 22204
rect 24137 22148 24176 22200
rect 24228 22148 24267 22200
rect 24137 22147 24267 22148
rect 24137 22101 24180 22147
rect 24226 22101 24267 22147
rect 24137 22044 24267 22101
rect 24137 21998 24180 22044
rect 24226 21998 24267 22044
rect 24137 21982 24267 21998
rect 24137 21930 24176 21982
rect 24228 21930 24267 21982
rect 24137 21894 24180 21930
rect 24226 21894 24267 21930
rect 23956 21881 24002 21889
rect 15431 21796 15469 21836
rect 15345 21744 15381 21796
rect 15433 21744 15469 21796
rect 16781 21787 16896 21800
rect 17901 21787 18016 21800
rect 18414 21787 18529 21800
rect 19534 21787 19649 21800
rect 24137 21787 24267 21894
rect 24694 23795 24740 23852
rect 24694 23692 24740 23749
rect 24694 23589 24740 23646
rect 24694 23486 24740 23543
rect 24694 23383 24740 23440
rect 24694 23280 24740 23337
rect 24694 23177 24740 23234
rect 24694 23074 24740 23131
rect 24694 22971 24740 23028
rect 24694 22868 24740 22925
rect 24694 22765 24740 22822
rect 24694 22662 24740 22719
rect 24694 22559 24740 22616
rect 24694 22456 24740 22513
rect 24694 22353 24740 22410
rect 24694 22250 24740 22307
rect 24470 22147 24516 22204
rect 24470 22044 24516 22101
rect 24470 21940 24516 21998
rect 24470 21881 24516 21894
rect 24654 22204 24694 22240
rect 25246 24779 25646 24802
rect 25692 24780 25739 24825
rect 25246 24766 25649 24779
rect 25246 24720 25281 24766
rect 25327 24728 25649 24766
rect 25701 24728 25739 24780
rect 25327 24722 25739 24728
rect 25327 24720 25646 24722
rect 25246 24676 25646 24720
rect 25692 24676 25739 24722
rect 25246 24619 25739 24676
rect 25246 24602 25646 24619
rect 25246 24556 25281 24602
rect 25327 24573 25646 24602
rect 25692 24573 25739 24619
rect 25327 24562 25739 24573
rect 25327 24556 25649 24562
rect 25246 24516 25649 24556
rect 25246 24470 25646 24516
rect 25701 24510 25739 24562
rect 25692 24470 25739 24510
rect 25246 24439 25739 24470
rect 25246 24393 25281 24439
rect 25327 24413 25739 24439
rect 25327 24393 25646 24413
rect 25246 24367 25646 24393
rect 25692 24367 25739 24413
rect 25246 24344 25739 24367
rect 25246 24310 25649 24344
rect 25246 24276 25646 24310
rect 25701 24292 25739 24344
rect 25246 24230 25281 24276
rect 25327 24264 25646 24276
rect 25692 24264 25739 24292
rect 25327 24230 25739 24264
rect 25246 24207 25739 24230
rect 25246 24161 25646 24207
rect 25692 24161 25739 24207
rect 25246 24126 25739 24161
rect 25246 24113 25649 24126
rect 25246 24067 25281 24113
rect 25327 24104 25649 24113
rect 25327 24067 25646 24104
rect 25701 24074 25739 24126
rect 25246 24058 25646 24067
rect 25692 24058 25739 24074
rect 25246 24001 25739 24058
rect 25246 23955 25646 24001
rect 25692 23955 25739 24001
rect 25246 23950 25739 23955
rect 25246 23904 25281 23950
rect 25327 23909 25739 23950
rect 25327 23904 25649 23909
rect 25246 23898 25649 23904
rect 25246 23852 25646 23898
rect 25701 23857 25739 23909
rect 25692 23852 25739 23857
rect 25246 23817 25739 23852
rect 25870 25031 25916 25072
rect 26160 25038 26206 25088
rect 26349 25134 26464 25440
rect 26986 25486 27417 25544
rect 27561 26730 27607 26743
rect 27561 26627 27607 26684
rect 27561 26524 27607 26581
rect 27851 26730 27897 26743
rect 27851 26627 27897 26684
rect 27851 26575 27897 26581
rect 28075 26730 28121 26743
rect 28075 26627 28121 26684
rect 27561 26421 27607 26478
rect 27561 26318 27607 26375
rect 27561 26214 27607 26272
rect 27561 26110 27607 26168
rect 27561 26006 27607 26064
rect 27561 25902 27607 25960
rect 27561 25798 27607 25856
rect 27809 26535 27937 26575
rect 27809 26483 27847 26535
rect 27899 26483 27937 26535
rect 27809 26478 27851 26483
rect 27897 26478 27937 26483
rect 27809 26421 27937 26478
rect 27809 26375 27851 26421
rect 27897 26375 27937 26421
rect 27809 26318 27937 26375
rect 27809 26317 27851 26318
rect 27897 26317 27937 26318
rect 27809 26265 27847 26317
rect 27899 26265 27937 26317
rect 27809 26214 27937 26265
rect 27809 26168 27851 26214
rect 27897 26168 27937 26214
rect 27809 26110 27937 26168
rect 27809 26099 27851 26110
rect 27897 26099 27937 26110
rect 27809 26047 27847 26099
rect 27899 26047 27937 26099
rect 27809 26006 27937 26047
rect 27809 25960 27851 26006
rect 27897 25960 27937 26006
rect 27809 25902 27937 25960
rect 27809 25881 27851 25902
rect 27897 25881 27937 25902
rect 27809 25829 27847 25881
rect 27899 25829 27937 25881
rect 27809 25798 27937 25829
rect 27809 25789 27851 25798
rect 27561 25694 27607 25752
rect 27561 25590 27607 25648
rect 27561 25496 27607 25544
rect 27897 25789 27937 25798
rect 28075 26524 28121 26581
rect 28075 26421 28121 26478
rect 28075 26318 28121 26375
rect 28075 26214 28121 26272
rect 28075 26110 28121 26168
rect 28075 26006 28121 26064
rect 28075 25902 28121 25960
rect 28075 25798 28121 25856
rect 27851 25694 27897 25752
rect 27851 25590 27897 25648
rect 26986 25440 27337 25486
rect 27383 25440 27417 25486
rect 26986 25435 27417 25440
rect 27526 25486 27641 25496
rect 27526 25440 27561 25486
rect 27607 25440 27641 25486
rect 27337 25427 27383 25435
rect 27082 25346 27422 25353
rect 27526 25346 27641 25440
rect 27851 25486 27897 25544
rect 28075 25694 28121 25752
rect 28075 25590 28121 25648
rect 28075 25496 28121 25544
rect 27851 25427 27897 25440
rect 28040 25486 28155 25496
rect 28040 25440 28075 25486
rect 28121 25440 28155 25486
rect 27082 25312 27439 25346
rect 27082 25260 27120 25312
rect 27172 25309 27332 25312
rect 27384 25309 27439 25312
rect 27172 25263 27200 25309
rect 27246 25263 27332 25309
rect 27404 25263 27439 25309
rect 27172 25260 27332 25263
rect 27384 25260 27439 25263
rect 27082 25226 27439 25260
rect 27526 25309 27949 25346
rect 27526 25263 27710 25309
rect 27756 25263 27868 25309
rect 27914 25263 27949 25309
rect 27526 25226 27949 25263
rect 27082 25220 27422 25226
rect 27337 25137 27383 25147
rect 26349 25088 26384 25134
rect 26430 25088 26464 25134
rect 26349 25072 26464 25088
rect 27012 25134 27417 25137
rect 27012 25088 27337 25134
rect 27383 25088 27417 25134
rect 25870 24928 25916 24985
rect 25870 24825 25916 24882
rect 25870 24722 25916 24779
rect 25870 24619 25916 24676
rect 25870 24516 25916 24573
rect 25870 24413 25916 24470
rect 25870 24310 25916 24367
rect 25870 24207 25916 24264
rect 25870 24104 25916 24161
rect 25870 24001 25916 24058
rect 25870 23898 25916 23955
rect 25246 23816 25733 23817
rect 25246 23795 25726 23816
rect 25246 23786 25646 23795
rect 25246 23740 25281 23786
rect 25327 23749 25646 23786
rect 25692 23749 25726 23795
rect 25327 23740 25726 23749
rect 25246 23692 25726 23740
rect 25246 23646 25646 23692
rect 25692 23646 25726 23692
rect 25246 23623 25726 23646
rect 25246 23577 25281 23623
rect 25327 23589 25726 23623
rect 25327 23577 25646 23589
rect 25246 23543 25646 23577
rect 25692 23543 25726 23589
rect 25246 23486 25726 23543
rect 25246 23460 25646 23486
rect 25246 23414 25281 23460
rect 25327 23440 25646 23460
rect 25692 23440 25726 23486
rect 25327 23414 25726 23440
rect 25246 23383 25726 23414
rect 25246 23337 25646 23383
rect 25692 23337 25726 23383
rect 25246 23296 25726 23337
rect 25246 23250 25281 23296
rect 25327 23280 25726 23296
rect 25327 23250 25646 23280
rect 25246 23234 25646 23250
rect 25692 23234 25726 23280
rect 25246 23177 25726 23234
rect 25246 23133 25646 23177
rect 25246 23087 25281 23133
rect 25327 23131 25646 23133
rect 25692 23131 25726 23177
rect 25327 23087 25726 23131
rect 25246 23074 25726 23087
rect 25246 23028 25646 23074
rect 25692 23028 25726 23074
rect 25246 22971 25726 23028
rect 25246 22970 25646 22971
rect 25246 22924 25281 22970
rect 25327 22925 25646 22970
rect 25692 22925 25726 22971
rect 25327 22924 25726 22925
rect 25246 22868 25726 22924
rect 25246 22822 25646 22868
rect 25692 22822 25726 22868
rect 25246 22806 25726 22822
rect 25246 22760 25281 22806
rect 25327 22765 25726 22806
rect 25327 22760 25646 22765
rect 25246 22719 25646 22760
rect 25692 22719 25726 22765
rect 25246 22662 25726 22719
rect 25246 22643 25646 22662
rect 25246 22597 25281 22643
rect 25327 22616 25646 22643
rect 25692 22616 25726 22662
rect 25327 22597 25726 22616
rect 25246 22559 25726 22597
rect 25246 22513 25646 22559
rect 25692 22513 25726 22559
rect 25246 22480 25726 22513
rect 25246 22434 25281 22480
rect 25327 22456 25726 22480
rect 25327 22434 25646 22456
rect 25246 22410 25646 22434
rect 25692 22410 25726 22456
rect 25246 22353 25726 22410
rect 25246 22317 25646 22353
rect 25246 22271 25281 22317
rect 25327 22307 25646 22317
rect 25692 22307 25726 22353
rect 25327 22271 25726 22307
rect 25246 22250 25726 22271
rect 24740 22204 24778 22240
rect 24654 22200 24778 22204
rect 24654 22148 24690 22200
rect 24742 22148 24778 22200
rect 24654 22147 24778 22148
rect 24654 22101 24694 22147
rect 24740 22101 24778 22147
rect 24654 22044 24778 22101
rect 24654 21998 24694 22044
rect 24740 21998 24778 22044
rect 24654 21982 24778 21998
rect 24654 21930 24690 21982
rect 24742 21930 24778 21982
rect 24654 21894 24694 21930
rect 24740 21894 24778 21930
rect 25246 22204 25646 22250
rect 25692 22204 25726 22250
rect 25870 23795 25916 23852
rect 26125 25031 26253 25038
rect 26125 24985 26160 25031
rect 26206 24997 26253 25031
rect 26125 24945 26163 24985
rect 26215 24945 26253 24997
rect 26125 24928 26253 24945
rect 26125 24882 26160 24928
rect 26206 24882 26253 24928
rect 26125 24825 26253 24882
rect 26125 24779 26160 24825
rect 26206 24780 26253 24825
rect 26125 24728 26163 24779
rect 26215 24728 26253 24780
rect 26125 24722 26253 24728
rect 26125 24676 26160 24722
rect 26206 24676 26253 24722
rect 26125 24619 26253 24676
rect 26125 24573 26160 24619
rect 26206 24573 26253 24619
rect 26125 24562 26253 24573
rect 26125 24516 26163 24562
rect 26125 24470 26160 24516
rect 26215 24510 26253 24562
rect 26206 24470 26253 24510
rect 26125 24413 26253 24470
rect 26125 24367 26160 24413
rect 26206 24367 26253 24413
rect 26125 24344 26253 24367
rect 26125 24310 26163 24344
rect 26125 24264 26160 24310
rect 26215 24292 26253 24344
rect 26206 24264 26253 24292
rect 26125 24207 26253 24264
rect 26125 24161 26160 24207
rect 26206 24161 26253 24207
rect 26125 24126 26253 24161
rect 26125 24104 26163 24126
rect 26125 24058 26160 24104
rect 26215 24074 26253 24126
rect 26206 24058 26253 24074
rect 26125 24001 26253 24058
rect 26125 23955 26160 24001
rect 26206 23955 26253 24001
rect 26125 23909 26253 23955
rect 26125 23898 26163 23909
rect 26125 23852 26160 23898
rect 26215 23857 26253 23909
rect 26206 23852 26253 23857
rect 26125 23817 26253 23852
rect 26384 25031 26430 25072
rect 26384 24928 26430 24985
rect 26384 24825 26430 24882
rect 27012 25038 27417 25088
rect 27526 25134 27641 25226
rect 27526 25088 27561 25134
rect 27607 25088 27641 25134
rect 27526 25072 27641 25088
rect 27851 25134 27897 25147
rect 27012 25031 27430 25038
rect 27012 24985 27337 25031
rect 27383 24997 27430 25031
rect 27012 24945 27340 24985
rect 27392 24945 27430 24997
rect 27012 24928 27430 24945
rect 27012 24882 27337 24928
rect 27383 24882 27430 24928
rect 27012 24825 27430 24882
rect 27012 24802 27337 24825
rect 26384 24722 26430 24779
rect 26384 24619 26430 24676
rect 26384 24516 26430 24573
rect 26384 24413 26430 24470
rect 26384 24310 26430 24367
rect 26384 24207 26430 24264
rect 26384 24104 26430 24161
rect 26384 24001 26430 24058
rect 26384 23898 26430 23955
rect 26131 23816 26247 23817
rect 25870 23692 25916 23749
rect 25870 23589 25916 23646
rect 25870 23486 25916 23543
rect 25870 23383 25916 23440
rect 25870 23280 25916 23337
rect 25870 23177 25916 23234
rect 25870 23074 25916 23131
rect 25870 22971 25916 23028
rect 25870 22868 25916 22925
rect 25870 22765 25916 22822
rect 25870 22662 25916 22719
rect 25870 22559 25916 22616
rect 25870 22456 25916 22513
rect 25870 22353 25916 22410
rect 25870 22250 25916 22307
rect 25246 22154 25726 22204
rect 25246 22108 25281 22154
rect 25327 22147 25726 22154
rect 25327 22108 25646 22147
rect 25246 22101 25646 22108
rect 25692 22101 25726 22147
rect 25246 22044 25726 22101
rect 25246 21998 25646 22044
rect 25692 21998 25726 22044
rect 25246 21990 25726 21998
rect 25246 21944 25281 21990
rect 25327 21944 25726 21990
rect 25246 21940 25726 21944
rect 25246 21908 25646 21940
rect 25320 21907 25646 21908
rect 24654 21890 24778 21894
rect 25321 21894 25646 21907
rect 25692 21894 25726 21940
rect 24694 21881 24740 21890
rect 25321 21889 25726 21894
rect 25830 22204 25870 22240
rect 26160 23795 26206 23816
rect 26160 23692 26206 23749
rect 26160 23589 26206 23646
rect 26160 23486 26206 23543
rect 26160 23383 26206 23440
rect 26160 23280 26206 23337
rect 26160 23177 26206 23234
rect 26160 23074 26206 23131
rect 26160 22971 26206 23028
rect 26160 22868 26206 22925
rect 26160 22765 26206 22822
rect 26160 22662 26206 22719
rect 26160 22559 26206 22616
rect 26160 22456 26206 22513
rect 26160 22353 26206 22410
rect 26160 22250 26206 22307
rect 25916 22204 25954 22240
rect 25830 22200 25954 22204
rect 25830 22148 25866 22200
rect 25918 22148 25954 22200
rect 25830 22147 25954 22148
rect 25830 22101 25870 22147
rect 25916 22101 25954 22147
rect 25830 22044 25954 22101
rect 25830 21998 25870 22044
rect 25916 21998 25954 22044
rect 25830 21982 25954 21998
rect 25830 21930 25866 21982
rect 25918 21930 25954 21982
rect 25830 21894 25870 21930
rect 25916 21894 25954 21930
rect 25830 21890 25954 21894
rect 26384 23795 26430 23852
rect 26384 23692 26430 23749
rect 26384 23589 26430 23646
rect 26384 23486 26430 23543
rect 26384 23383 26430 23440
rect 26384 23280 26430 23337
rect 26384 23177 26430 23234
rect 26384 23074 26430 23131
rect 26384 22971 26430 23028
rect 26384 22868 26430 22925
rect 26384 22765 26430 22822
rect 26384 22662 26430 22719
rect 26384 22559 26430 22616
rect 26384 22456 26430 22513
rect 26384 22353 26430 22410
rect 26384 22250 26430 22307
rect 26160 22147 26206 22204
rect 26160 22044 26206 22101
rect 26160 21940 26206 21998
rect 25646 21881 25692 21889
rect 25870 21881 25916 21890
rect 26160 21881 26206 21894
rect 26344 22204 26384 22240
rect 26937 24779 27337 24802
rect 27383 24780 27430 24825
rect 26937 24766 27340 24779
rect 26937 24720 26972 24766
rect 27018 24728 27340 24766
rect 27392 24728 27430 24780
rect 27018 24722 27430 24728
rect 27018 24720 27337 24722
rect 26937 24676 27337 24720
rect 27383 24676 27430 24722
rect 26937 24619 27430 24676
rect 26937 24602 27337 24619
rect 26937 24556 26972 24602
rect 27018 24573 27337 24602
rect 27383 24573 27430 24619
rect 27018 24562 27430 24573
rect 27018 24556 27340 24562
rect 26937 24516 27340 24556
rect 26937 24470 27337 24516
rect 27392 24510 27430 24562
rect 27383 24470 27430 24510
rect 26937 24439 27430 24470
rect 26937 24393 26972 24439
rect 27018 24413 27430 24439
rect 27018 24393 27337 24413
rect 26937 24367 27337 24393
rect 27383 24367 27430 24413
rect 26937 24344 27430 24367
rect 26937 24310 27340 24344
rect 26937 24276 27337 24310
rect 27392 24292 27430 24344
rect 26937 24230 26972 24276
rect 27018 24264 27337 24276
rect 27383 24264 27430 24292
rect 27018 24230 27430 24264
rect 26937 24207 27430 24230
rect 26937 24161 27337 24207
rect 27383 24161 27430 24207
rect 26937 24126 27430 24161
rect 26937 24113 27340 24126
rect 26937 24067 26972 24113
rect 27018 24104 27340 24113
rect 27018 24067 27337 24104
rect 27392 24074 27430 24126
rect 26937 24058 27337 24067
rect 27383 24058 27430 24074
rect 26937 24001 27430 24058
rect 26937 23955 27337 24001
rect 27383 23955 27430 24001
rect 26937 23950 27430 23955
rect 26937 23904 26972 23950
rect 27018 23909 27430 23950
rect 27018 23904 27340 23909
rect 26937 23898 27340 23904
rect 26937 23852 27337 23898
rect 27392 23857 27430 23909
rect 27383 23852 27430 23857
rect 26937 23817 27430 23852
rect 27561 25031 27607 25072
rect 27851 25038 27897 25088
rect 28040 25134 28155 25440
rect 28040 25088 28075 25134
rect 28121 25088 28155 25134
rect 28040 25072 28155 25088
rect 27561 24928 27607 24985
rect 27561 24825 27607 24882
rect 27561 24722 27607 24779
rect 27561 24619 27607 24676
rect 27561 24516 27607 24573
rect 27561 24413 27607 24470
rect 27561 24310 27607 24367
rect 27561 24207 27607 24264
rect 27561 24104 27607 24161
rect 27561 24001 27607 24058
rect 27561 23898 27607 23955
rect 26937 23816 27424 23817
rect 26937 23795 27417 23816
rect 26937 23786 27337 23795
rect 26937 23740 26972 23786
rect 27018 23749 27337 23786
rect 27383 23749 27417 23795
rect 27018 23740 27417 23749
rect 26937 23692 27417 23740
rect 26937 23646 27337 23692
rect 27383 23646 27417 23692
rect 26937 23623 27417 23646
rect 26937 23577 26972 23623
rect 27018 23589 27417 23623
rect 27018 23577 27337 23589
rect 26937 23543 27337 23577
rect 27383 23543 27417 23589
rect 26937 23486 27417 23543
rect 26937 23460 27337 23486
rect 26937 23414 26972 23460
rect 27018 23440 27337 23460
rect 27383 23440 27417 23486
rect 27018 23414 27417 23440
rect 26937 23383 27417 23414
rect 26937 23337 27337 23383
rect 27383 23337 27417 23383
rect 26937 23296 27417 23337
rect 26937 23250 26972 23296
rect 27018 23280 27417 23296
rect 27018 23250 27337 23280
rect 26937 23234 27337 23250
rect 27383 23234 27417 23280
rect 26937 23177 27417 23234
rect 26937 23133 27337 23177
rect 26937 23087 26972 23133
rect 27018 23131 27337 23133
rect 27383 23131 27417 23177
rect 27018 23087 27417 23131
rect 26937 23074 27417 23087
rect 26937 23028 27337 23074
rect 27383 23028 27417 23074
rect 26937 22971 27417 23028
rect 26937 22970 27337 22971
rect 26937 22924 26972 22970
rect 27018 22925 27337 22970
rect 27383 22925 27417 22971
rect 27018 22924 27417 22925
rect 26937 22868 27417 22924
rect 26937 22822 27337 22868
rect 27383 22822 27417 22868
rect 26937 22806 27417 22822
rect 26937 22760 26972 22806
rect 27018 22765 27417 22806
rect 27018 22760 27337 22765
rect 26937 22719 27337 22760
rect 27383 22719 27417 22765
rect 26937 22662 27417 22719
rect 26937 22643 27337 22662
rect 26937 22597 26972 22643
rect 27018 22616 27337 22643
rect 27383 22616 27417 22662
rect 27018 22597 27417 22616
rect 26937 22559 27417 22597
rect 26937 22513 27337 22559
rect 27383 22513 27417 22559
rect 26937 22480 27417 22513
rect 26937 22434 26972 22480
rect 27018 22456 27417 22480
rect 27018 22434 27337 22456
rect 26937 22410 27337 22434
rect 27383 22410 27417 22456
rect 26937 22353 27417 22410
rect 26937 22317 27337 22353
rect 26937 22271 26972 22317
rect 27018 22307 27337 22317
rect 27383 22307 27417 22353
rect 27018 22271 27417 22307
rect 26937 22250 27417 22271
rect 26430 22204 26468 22240
rect 26344 22200 26468 22204
rect 26344 22148 26380 22200
rect 26432 22148 26468 22200
rect 26344 22147 26468 22148
rect 26344 22101 26384 22147
rect 26430 22101 26468 22147
rect 26344 22044 26468 22101
rect 26344 21998 26384 22044
rect 26430 21998 26468 22044
rect 26344 21982 26468 21998
rect 26344 21930 26380 21982
rect 26432 21930 26468 21982
rect 26344 21894 26384 21930
rect 26430 21894 26468 21930
rect 26937 22204 27337 22250
rect 27383 22204 27417 22250
rect 27561 23795 27607 23852
rect 27816 25031 27944 25038
rect 27816 24985 27851 25031
rect 27897 24997 27944 25031
rect 27816 24945 27854 24985
rect 27906 24945 27944 24997
rect 27816 24928 27944 24945
rect 27816 24882 27851 24928
rect 27897 24882 27944 24928
rect 27816 24825 27944 24882
rect 27816 24779 27851 24825
rect 27897 24780 27944 24825
rect 27816 24728 27854 24779
rect 27906 24728 27944 24780
rect 27816 24722 27944 24728
rect 27816 24676 27851 24722
rect 27897 24676 27944 24722
rect 27816 24619 27944 24676
rect 27816 24573 27851 24619
rect 27897 24573 27944 24619
rect 27816 24562 27944 24573
rect 27816 24516 27854 24562
rect 27816 24470 27851 24516
rect 27906 24510 27944 24562
rect 27897 24470 27944 24510
rect 27816 24413 27944 24470
rect 27816 24367 27851 24413
rect 27897 24367 27944 24413
rect 27816 24344 27944 24367
rect 27816 24310 27854 24344
rect 27816 24264 27851 24310
rect 27906 24292 27944 24344
rect 27897 24264 27944 24292
rect 27816 24207 27944 24264
rect 27816 24161 27851 24207
rect 27897 24161 27944 24207
rect 27816 24126 27944 24161
rect 27816 24104 27854 24126
rect 27816 24058 27851 24104
rect 27906 24074 27944 24126
rect 27897 24058 27944 24074
rect 27816 24001 27944 24058
rect 27816 23955 27851 24001
rect 27897 23955 27944 24001
rect 27816 23909 27944 23955
rect 27816 23898 27854 23909
rect 27816 23852 27851 23898
rect 27906 23857 27944 23909
rect 27897 23852 27944 23857
rect 27816 23817 27944 23852
rect 28075 25031 28121 25072
rect 28075 24928 28121 24985
rect 28075 24825 28121 24882
rect 28075 24722 28121 24779
rect 28075 24619 28121 24676
rect 28075 24516 28121 24573
rect 28075 24413 28121 24470
rect 28075 24310 28121 24367
rect 28075 24207 28121 24264
rect 28075 24104 28121 24161
rect 28075 24001 28121 24058
rect 28075 23898 28121 23955
rect 27822 23816 27938 23817
rect 27561 23692 27607 23749
rect 27561 23589 27607 23646
rect 27561 23486 27607 23543
rect 27561 23383 27607 23440
rect 27561 23280 27607 23337
rect 27561 23177 27607 23234
rect 27561 23074 27607 23131
rect 27561 22971 27607 23028
rect 27561 22868 27607 22925
rect 27561 22765 27607 22822
rect 27561 22662 27607 22719
rect 27561 22559 27607 22616
rect 27561 22456 27607 22513
rect 27561 22353 27607 22410
rect 27561 22250 27607 22307
rect 26937 22154 27417 22204
rect 26937 22108 26972 22154
rect 27018 22147 27417 22154
rect 27018 22108 27337 22147
rect 26937 22101 27337 22108
rect 27383 22101 27417 22147
rect 26937 22044 27417 22101
rect 26937 21998 27337 22044
rect 27383 21998 27417 22044
rect 26937 21990 27417 21998
rect 26937 21944 26972 21990
rect 27018 21944 27417 21990
rect 26937 21940 27417 21944
rect 26937 21908 27337 21940
rect 27011 21907 27337 21908
rect 26344 21890 26468 21894
rect 27012 21894 27337 21907
rect 27383 21894 27417 21940
rect 26384 21881 26430 21890
rect 27012 21889 27417 21894
rect 27521 22204 27561 22240
rect 27851 23795 27897 23816
rect 27851 23692 27897 23749
rect 27851 23589 27897 23646
rect 27851 23486 27897 23543
rect 27851 23383 27897 23440
rect 27851 23280 27897 23337
rect 27851 23177 27897 23234
rect 27851 23074 27897 23131
rect 27851 22971 27897 23028
rect 27851 22868 27897 22925
rect 27851 22765 27897 22822
rect 27851 22662 27897 22719
rect 27851 22559 27897 22616
rect 27851 22456 27897 22513
rect 27851 22353 27897 22410
rect 27851 22250 27897 22307
rect 27607 22204 27645 22240
rect 27521 22200 27645 22204
rect 27521 22148 27557 22200
rect 27609 22148 27645 22200
rect 27521 22147 27645 22148
rect 27521 22101 27561 22147
rect 27607 22101 27645 22147
rect 27521 22044 27645 22101
rect 27521 21998 27561 22044
rect 27607 21998 27645 22044
rect 27521 21982 27645 21998
rect 27521 21930 27557 21982
rect 27609 21930 27645 21982
rect 27521 21894 27561 21930
rect 27607 21894 27645 21930
rect 27521 21890 27645 21894
rect 28075 23795 28121 23852
rect 28075 23692 28121 23749
rect 28075 23589 28121 23646
rect 28075 23486 28121 23543
rect 28075 23383 28121 23440
rect 28075 23280 28121 23337
rect 28075 23177 28121 23234
rect 28075 23074 28121 23131
rect 28075 22971 28121 23028
rect 28075 22868 28121 22925
rect 28075 22765 28121 22822
rect 28075 22662 28121 22719
rect 28075 22559 28121 22616
rect 28075 22456 28121 22513
rect 28075 22353 28121 22410
rect 28075 22250 28121 22307
rect 27851 22147 27897 22204
rect 27851 22044 27897 22101
rect 27851 21940 27897 21998
rect 27337 21881 27383 21889
rect 27561 21881 27607 21890
rect 27851 21881 27897 21894
rect 28035 22204 28075 22240
rect 28121 22204 28159 22240
rect 28035 22200 28159 22204
rect 28035 22148 28071 22200
rect 28123 22148 28159 22200
rect 28035 22147 28159 22148
rect 28035 22101 28075 22147
rect 28121 22101 28159 22147
rect 28035 22044 28159 22101
rect 28035 21998 28075 22044
rect 28121 21998 28159 22044
rect 28035 21982 28159 21998
rect 28035 21930 28071 21982
rect 28123 21930 28159 21982
rect 28035 21894 28075 21930
rect 28121 21894 28159 21930
rect 28035 21890 28159 21894
rect 28075 21881 28121 21890
rect 15345 21578 15385 21744
rect 15431 21578 15469 21744
rect 16524 21764 28485 21787
rect 16524 21718 16816 21764
rect 16862 21718 17936 21764
rect 17982 21718 18449 21764
rect 18495 21718 19569 21764
rect 19615 21718 28485 21764
rect 16524 21695 28485 21718
rect 16781 21681 16896 21695
rect 17901 21681 18016 21695
rect 18414 21681 18529 21695
rect 19534 21681 19649 21695
rect 23174 21694 28485 21695
rect 17005 21585 17120 21600
rect 17677 21585 17792 21600
rect 20272 21585 20387 21600
rect 20944 21585 21059 21600
rect 25828 21585 25957 21606
rect 15345 21526 15381 21578
rect 15433 21526 15469 21578
rect 15345 21490 15385 21526
rect 15431 21490 15469 21526
rect 16524 21565 28485 21585
rect 16524 21564 25867 21565
rect 16524 21518 17040 21564
rect 17086 21518 17712 21564
rect 17758 21518 20307 21564
rect 20353 21518 20979 21564
rect 21025 21518 25867 21564
rect 16524 21513 25867 21518
rect 25919 21513 28485 21565
rect 16524 21493 28485 21513
rect 15345 21486 15469 21490
rect 15161 21477 15207 21486
rect 15385 21477 15431 21486
rect 17005 21481 17120 21493
rect 17677 21481 17792 21493
rect 20272 21481 20387 21493
rect 20944 21481 21059 21493
rect 23174 21492 28485 21493
rect 25828 21472 25957 21492
rect 17229 21383 17344 21396
rect 18862 21383 18977 21396
rect 20496 21383 20611 21396
rect 22130 21383 22245 21396
rect 27519 21383 27648 21404
rect 1583 21363 8866 21383
rect 1583 21317 1929 21363
rect 1975 21317 3181 21363
rect 3227 21317 8866 21363
rect 1583 21291 8866 21317
rect 8962 21363 16245 21383
rect 8962 21317 9308 21363
rect 9354 21317 10560 21363
rect 10606 21317 16245 21363
rect 8962 21291 16245 21317
rect 16524 21363 28485 21383
rect 16524 21360 27558 21363
rect 16524 21314 17264 21360
rect 17310 21314 18897 21360
rect 18943 21314 20531 21360
rect 20577 21314 22165 21360
rect 22211 21314 27558 21360
rect 16524 21311 27558 21314
rect 27610 21311 28485 21363
rect 16524 21292 28485 21311
rect 1894 21280 2009 21291
rect 3146 21280 3261 21291
rect 9273 21280 9388 21291
rect 10525 21280 10640 21291
rect 17229 21277 17344 21292
rect 18862 21277 18977 21292
rect 20496 21277 20611 21292
rect 22130 21277 22245 21292
rect 23174 21291 28485 21292
rect 27519 21270 27648 21291
rect 3686 21182 3801 21195
rect 4938 21182 5053 21195
rect 6787 21182 6916 21203
rect 11065 21182 11180 21195
rect 12317 21182 12432 21195
rect 14166 21182 14295 21203
rect 20048 21182 20163 21195
rect 21168 21182 21283 21195
rect 21682 21182 21797 21195
rect 22802 21182 22917 21195
rect 24651 21182 24780 21203
rect 1583 21162 8866 21182
rect 1583 21159 6825 21162
rect 1583 21113 3721 21159
rect 3767 21113 4973 21159
rect 5019 21113 6825 21159
rect 1583 21110 6825 21113
rect 6877 21110 8866 21162
rect 1583 21089 8866 21110
rect 8962 21162 16245 21182
rect 8962 21159 14204 21162
rect 8962 21113 11100 21159
rect 11146 21113 12352 21159
rect 12398 21113 14204 21159
rect 8962 21110 14204 21113
rect 14256 21110 16245 21162
rect 8962 21089 16245 21110
rect 16524 21162 28485 21182
rect 16524 21159 24690 21162
rect 16524 21113 20083 21159
rect 20129 21113 21203 21159
rect 21249 21113 21717 21159
rect 21763 21113 22837 21159
rect 22883 21113 24690 21159
rect 16524 21110 24690 21113
rect 24742 21110 28485 21162
rect 16524 21090 28485 21110
rect 3686 21076 3801 21089
rect 4938 21076 5053 21089
rect 6787 21069 6916 21089
rect 11065 21076 11180 21089
rect 12317 21076 12432 21089
rect 14166 21069 14295 21089
rect 20048 21076 20163 21090
rect 21168 21076 21283 21090
rect 21682 21076 21797 21090
rect 22802 21076 22917 21090
rect 23174 21089 28485 21090
rect 24651 21069 24780 21089
rect 2118 20980 2233 20991
rect 3910 20980 4025 20991
rect 7964 20980 8093 21001
rect 9497 20980 9612 20991
rect 11289 20980 11404 20991
rect 15343 20980 15472 21001
rect 18638 20980 18753 20993
rect 19310 20980 19425 20993
rect 21906 20980 22021 20993
rect 22578 20980 22693 20993
rect 26342 20980 26471 21001
rect 1583 20960 8866 20980
rect 1583 20955 8002 20960
rect 1583 20909 2153 20955
rect 2199 20909 3945 20955
rect 3991 20909 8002 20955
rect 1583 20908 8002 20909
rect 8054 20908 8866 20960
rect 1583 20888 8866 20908
rect 8962 20960 16245 20980
rect 8962 20955 15381 20960
rect 8962 20909 9532 20955
rect 9578 20909 11324 20955
rect 11370 20909 15381 20955
rect 8962 20908 15381 20909
rect 15433 20908 16245 20960
rect 8962 20888 16245 20908
rect 16524 20960 28485 20980
rect 16524 20957 26381 20960
rect 16524 20911 18673 20957
rect 18719 20911 19345 20957
rect 19391 20911 21941 20957
rect 21987 20911 22613 20957
rect 22659 20911 26381 20957
rect 16524 20908 26381 20911
rect 26433 20908 28485 20960
rect 16524 20888 28485 20908
rect 2118 20872 2233 20888
rect 3910 20872 4025 20888
rect 5309 20887 8866 20888
rect 7964 20867 8093 20887
rect 9497 20872 9612 20888
rect 11289 20872 11404 20888
rect 12688 20887 16245 20888
rect 15343 20867 15472 20887
rect 18638 20874 18753 20888
rect 19310 20874 19425 20888
rect 21906 20874 22021 20888
rect 22578 20874 22693 20888
rect 23174 20887 28485 20888
rect 26342 20867 26471 20887
rect 2922 20778 3037 20791
rect 4714 20778 4829 20791
rect 8478 20778 8607 20799
rect 10301 20778 10416 20791
rect 12093 20778 12208 20791
rect 15857 20778 15986 20799
rect 17453 20778 17568 20791
rect 19086 20778 19201 20791
rect 20720 20778 20835 20791
rect 22354 20778 22469 20791
rect 28033 20778 28162 20799
rect 1583 20758 8866 20778
rect 1583 20755 8516 20758
rect 1583 20709 2957 20755
rect 3003 20709 4749 20755
rect 4795 20709 8516 20755
rect 1583 20706 8516 20709
rect 8568 20706 8866 20758
rect 1583 20686 8866 20706
rect 8962 20758 16245 20778
rect 8962 20755 15895 20758
rect 8962 20709 10336 20755
rect 10382 20709 12128 20755
rect 12174 20709 15895 20755
rect 8962 20706 15895 20709
rect 15947 20706 16245 20758
rect 8962 20686 16245 20706
rect 16524 20758 28485 20778
rect 16524 20755 28072 20758
rect 16524 20709 17488 20755
rect 17534 20709 19121 20755
rect 19167 20709 20755 20755
rect 20801 20709 22389 20755
rect 22435 20709 28072 20755
rect 16524 20706 28072 20709
rect 28124 20706 28485 20758
rect 16524 20686 28485 20706
rect 2922 20672 3037 20686
rect 4714 20672 4829 20686
rect 5309 20685 8866 20686
rect 8478 20665 8607 20685
rect 10301 20672 10416 20686
rect 12093 20672 12208 20686
rect 12688 20685 16245 20686
rect 15857 20665 15986 20685
rect 17453 20672 17568 20686
rect 19086 20672 19201 20686
rect 20720 20672 20835 20686
rect 22354 20672 22469 20686
rect 23174 20685 28485 20686
rect 28033 20665 28162 20685
rect 1776 20506 1903 20542
rect 1776 20502 1817 20506
rect 1863 20502 1903 20506
rect 1776 20450 1814 20502
rect 1866 20450 1903 20502
rect 1776 20338 1903 20450
rect 1776 20292 1817 20338
rect 1863 20292 1903 20338
rect 1776 20284 1903 20292
rect 1776 20232 1814 20284
rect 1866 20232 1903 20284
rect 1776 20171 1903 20232
rect 1776 20125 1817 20171
rect 1863 20125 1903 20171
rect 1776 20067 1903 20125
rect 1776 20015 1814 20067
rect 1866 20015 1903 20067
rect 1776 20003 1903 20015
rect 1776 19957 1817 20003
rect 1863 19957 1903 20003
rect 1776 19849 1903 19957
rect 1776 19797 1814 19849
rect 1866 19797 1903 19849
rect 1776 19789 1817 19797
rect 1863 19789 1903 19797
rect 1776 19667 1903 19789
rect 1776 19631 1817 19667
rect 1863 19631 1903 19667
rect 1776 19579 1814 19631
rect 1866 19579 1903 19631
rect 1776 19499 1903 19579
rect 1776 19453 1817 19499
rect 1863 19453 1903 19499
rect 1776 19413 1903 19453
rect 1776 19361 1814 19413
rect 1866 19361 1903 19413
rect 1776 19332 1903 19361
rect 1776 19286 1817 19332
rect 1863 19286 1903 19332
rect 1776 19196 1903 19286
rect 1776 19144 1814 19196
rect 1866 19144 1903 19196
rect 1776 19118 1817 19144
rect 1863 19118 1903 19144
rect 1776 18996 1903 19118
rect 1776 18978 1817 18996
rect 1863 18978 1903 18996
rect 1776 18926 1814 18978
rect 1866 18926 1903 18978
rect 1776 18886 1903 18926
rect 2230 20506 2926 20542
rect 2230 20460 2266 20506
rect 2312 20492 2844 20506
rect 2312 20460 2555 20492
rect 2230 20446 2555 20460
rect 2601 20460 2844 20492
rect 2890 20460 2926 20506
rect 2601 20446 2926 20460
rect 2230 20364 2926 20446
rect 2230 20338 2269 20364
rect 2230 20292 2266 20338
rect 2321 20312 2552 20364
rect 2604 20312 2835 20364
rect 2887 20338 2926 20364
rect 2312 20292 2555 20312
rect 2230 20283 2555 20292
rect 2601 20292 2844 20312
rect 2890 20292 2926 20338
rect 2601 20283 2926 20292
rect 2230 20171 2926 20283
rect 2230 20125 2266 20171
rect 2312 20166 2844 20171
rect 2312 20146 2555 20166
rect 2601 20146 2844 20166
rect 2230 20094 2269 20125
rect 2321 20094 2552 20146
rect 2604 20094 2835 20146
rect 2890 20125 2926 20171
rect 2887 20094 2926 20125
rect 2230 20003 2926 20094
rect 2230 19957 2266 20003
rect 2312 19957 2555 20003
rect 2601 19957 2844 20003
rect 2890 19957 2926 20003
rect 2230 19929 2926 19957
rect 2230 19877 2269 19929
rect 2321 19877 2552 19929
rect 2604 19877 2835 19929
rect 2887 19877 2926 19929
rect 2230 19840 2926 19877
rect 2230 19835 2555 19840
rect 2230 19789 2266 19835
rect 2312 19794 2555 19835
rect 2601 19835 2926 19840
rect 2601 19794 2844 19835
rect 2312 19789 2844 19794
rect 2890 19789 2926 19835
rect 2230 19711 2926 19789
rect 2230 19667 2269 19711
rect 2230 19621 2266 19667
rect 2321 19659 2552 19711
rect 2604 19659 2835 19711
rect 2887 19667 2926 19711
rect 2312 19630 2555 19659
rect 2601 19630 2844 19659
rect 2312 19621 2844 19630
rect 2890 19621 2926 19667
rect 2230 19513 2926 19621
rect 2230 19499 2555 19513
rect 2230 19453 2266 19499
rect 2312 19494 2555 19499
rect 2601 19499 2926 19513
rect 2601 19494 2844 19499
rect 2230 19442 2269 19453
rect 2321 19442 2552 19494
rect 2604 19442 2835 19494
rect 2890 19453 2926 19499
rect 2887 19442 2926 19453
rect 2230 19350 2926 19442
rect 2230 19332 2555 19350
rect 2230 19286 2266 19332
rect 2312 19304 2555 19332
rect 2601 19332 2926 19350
rect 2601 19304 2844 19332
rect 2312 19286 2844 19304
rect 2890 19286 2926 19332
rect 2230 19276 2926 19286
rect 2230 19224 2269 19276
rect 2321 19224 2552 19276
rect 2604 19224 2835 19276
rect 2887 19224 2926 19276
rect 2230 19187 2926 19224
rect 2230 19164 2555 19187
rect 2230 19118 2266 19164
rect 2312 19141 2555 19164
rect 2601 19164 2926 19187
rect 2601 19141 2844 19164
rect 2312 19118 2844 19141
rect 2890 19118 2926 19164
rect 2230 19058 2926 19118
rect 2230 19006 2269 19058
rect 2321 19006 2552 19058
rect 2604 19006 2835 19058
rect 2887 19006 2926 19058
rect 2230 18996 2555 19006
rect 2230 18950 2266 18996
rect 2312 18977 2555 18996
rect 2601 18996 2926 19006
rect 2601 18977 2844 18996
rect 2312 18950 2844 18977
rect 2890 18950 2926 18996
rect 1781 18885 1898 18886
rect 1781 18828 1897 18885
rect 1781 18782 1817 18828
rect 1863 18782 1897 18828
rect 1781 18658 1897 18782
rect 1781 18612 1817 18658
rect 1863 18612 1897 18658
rect 1781 18488 1897 18612
rect 1781 18442 1817 18488
rect 1863 18442 1897 18488
rect 1781 18318 1897 18442
rect 1781 18272 1817 18318
rect 1863 18272 1897 18318
rect 1781 18110 1897 18272
rect 2230 18860 2926 18950
rect 3253 20506 3380 20542
rect 3253 20502 3293 20506
rect 3339 20502 3380 20506
rect 3253 20450 3290 20502
rect 3342 20450 3380 20502
rect 3253 20338 3380 20450
rect 3253 20292 3293 20338
rect 3339 20292 3380 20338
rect 3253 20284 3380 20292
rect 3253 20232 3290 20284
rect 3342 20232 3380 20284
rect 3253 20171 3380 20232
rect 3253 20125 3293 20171
rect 3339 20125 3380 20171
rect 3253 20067 3380 20125
rect 3253 20015 3290 20067
rect 3342 20015 3380 20067
rect 3253 20003 3380 20015
rect 3253 19957 3293 20003
rect 3339 19957 3380 20003
rect 3253 19849 3380 19957
rect 3253 19797 3290 19849
rect 3342 19797 3380 19849
rect 3253 19789 3293 19797
rect 3339 19789 3380 19797
rect 3253 19667 3380 19789
rect 3253 19631 3293 19667
rect 3339 19631 3380 19667
rect 3253 19579 3290 19631
rect 3342 19579 3380 19631
rect 3253 19499 3380 19579
rect 3253 19453 3293 19499
rect 3339 19453 3380 19499
rect 3253 19413 3380 19453
rect 3253 19361 3290 19413
rect 3342 19361 3380 19413
rect 3253 19332 3380 19361
rect 3253 19286 3293 19332
rect 3339 19286 3380 19332
rect 3253 19196 3380 19286
rect 3253 19144 3290 19196
rect 3342 19144 3380 19196
rect 3253 19118 3293 19144
rect 3339 19118 3380 19144
rect 3253 18996 3380 19118
rect 3253 18978 3293 18996
rect 3339 18978 3380 18996
rect 3253 18926 3290 18978
rect 3342 18926 3380 18978
rect 3253 18886 3380 18926
rect 3568 20506 3695 20542
rect 3568 20502 3609 20506
rect 3655 20502 3695 20506
rect 3568 20450 3606 20502
rect 3658 20450 3695 20502
rect 3568 20338 3695 20450
rect 3568 20292 3609 20338
rect 3655 20292 3695 20338
rect 3568 20284 3695 20292
rect 3568 20232 3606 20284
rect 3658 20232 3695 20284
rect 3568 20171 3695 20232
rect 3568 20125 3609 20171
rect 3655 20125 3695 20171
rect 3568 20067 3695 20125
rect 3568 20015 3606 20067
rect 3658 20015 3695 20067
rect 3568 20003 3695 20015
rect 3568 19957 3609 20003
rect 3655 19957 3695 20003
rect 3568 19849 3695 19957
rect 3568 19797 3606 19849
rect 3658 19797 3695 19849
rect 3568 19789 3609 19797
rect 3655 19789 3695 19797
rect 3568 19667 3695 19789
rect 3568 19631 3609 19667
rect 3655 19631 3695 19667
rect 3568 19579 3606 19631
rect 3658 19579 3695 19631
rect 3568 19499 3695 19579
rect 3568 19453 3609 19499
rect 3655 19453 3695 19499
rect 3568 19413 3695 19453
rect 3568 19361 3606 19413
rect 3658 19361 3695 19413
rect 3568 19332 3695 19361
rect 3568 19286 3609 19332
rect 3655 19286 3695 19332
rect 3568 19196 3695 19286
rect 3568 19144 3606 19196
rect 3658 19144 3695 19196
rect 3568 19118 3609 19144
rect 3655 19118 3695 19144
rect 3568 18996 3695 19118
rect 3568 18978 3609 18996
rect 3655 18978 3695 18996
rect 3568 18926 3606 18978
rect 3658 18926 3695 18978
rect 3568 18886 3695 18926
rect 4022 20506 4718 20542
rect 4022 20460 4058 20506
rect 4104 20492 4636 20506
rect 4104 20460 4347 20492
rect 4022 20446 4347 20460
rect 4393 20460 4636 20492
rect 4682 20460 4718 20506
rect 4393 20446 4718 20460
rect 4022 20364 4718 20446
rect 4022 20338 4061 20364
rect 4022 20292 4058 20338
rect 4113 20312 4344 20364
rect 4396 20312 4627 20364
rect 4679 20338 4718 20364
rect 4104 20292 4347 20312
rect 4022 20283 4347 20292
rect 4393 20292 4636 20312
rect 4682 20292 4718 20338
rect 4393 20283 4718 20292
rect 4022 20171 4718 20283
rect 4022 20125 4058 20171
rect 4104 20166 4636 20171
rect 4104 20146 4347 20166
rect 4393 20146 4636 20166
rect 4022 20094 4061 20125
rect 4113 20094 4344 20146
rect 4396 20094 4627 20146
rect 4682 20125 4718 20171
rect 4679 20094 4718 20125
rect 4022 20003 4718 20094
rect 4022 19957 4058 20003
rect 4104 19957 4347 20003
rect 4393 19957 4636 20003
rect 4682 19957 4718 20003
rect 4022 19929 4718 19957
rect 4022 19877 4061 19929
rect 4113 19877 4344 19929
rect 4396 19877 4627 19929
rect 4679 19877 4718 19929
rect 4022 19840 4718 19877
rect 4022 19835 4347 19840
rect 4022 19789 4058 19835
rect 4104 19794 4347 19835
rect 4393 19835 4718 19840
rect 4393 19794 4636 19835
rect 4104 19789 4636 19794
rect 4682 19789 4718 19835
rect 4022 19711 4718 19789
rect 4022 19667 4061 19711
rect 4022 19621 4058 19667
rect 4113 19659 4344 19711
rect 4396 19659 4627 19711
rect 4679 19667 4718 19711
rect 4104 19630 4347 19659
rect 4393 19630 4636 19659
rect 4104 19621 4636 19630
rect 4682 19621 4718 19667
rect 4022 19513 4718 19621
rect 4022 19499 4347 19513
rect 4022 19453 4058 19499
rect 4104 19494 4347 19499
rect 4393 19499 4718 19513
rect 4393 19494 4636 19499
rect 4022 19442 4061 19453
rect 4113 19442 4344 19494
rect 4396 19442 4627 19494
rect 4682 19453 4718 19499
rect 4679 19442 4718 19453
rect 4022 19350 4718 19442
rect 4022 19332 4347 19350
rect 4022 19286 4058 19332
rect 4104 19304 4347 19332
rect 4393 19332 4718 19350
rect 4393 19304 4636 19332
rect 4104 19286 4636 19304
rect 4682 19286 4718 19332
rect 4022 19276 4718 19286
rect 4022 19224 4061 19276
rect 4113 19224 4344 19276
rect 4396 19224 4627 19276
rect 4679 19224 4718 19276
rect 4022 19187 4718 19224
rect 4022 19164 4347 19187
rect 4022 19118 4058 19164
rect 4104 19141 4347 19164
rect 4393 19164 4718 19187
rect 4393 19141 4636 19164
rect 4104 19118 4636 19141
rect 4682 19118 4718 19164
rect 4022 19058 4718 19118
rect 4022 19006 4061 19058
rect 4113 19006 4344 19058
rect 4396 19006 4627 19058
rect 4679 19006 4718 19058
rect 4022 18996 4347 19006
rect 4022 18950 4058 18996
rect 4104 18977 4347 18996
rect 4393 18996 4718 19006
rect 4393 18977 4636 18996
rect 4104 18950 4636 18977
rect 4682 18950 4718 18996
rect 3258 18885 3375 18886
rect 2230 18840 2555 18860
rect 2601 18840 2926 18860
rect 2230 18828 2269 18840
rect 2230 18782 2266 18828
rect 2321 18788 2552 18840
rect 2604 18788 2835 18840
rect 2887 18828 2926 18840
rect 2312 18782 2844 18788
rect 2890 18782 2926 18828
rect 2230 18697 2926 18782
rect 2230 18658 2555 18697
rect 2230 18612 2266 18658
rect 2312 18651 2555 18658
rect 2601 18658 2926 18697
rect 2601 18651 2844 18658
rect 2312 18623 2844 18651
rect 2230 18571 2269 18612
rect 2321 18571 2552 18623
rect 2604 18571 2835 18623
rect 2890 18612 2926 18658
rect 2887 18571 2926 18612
rect 2230 18534 2926 18571
rect 2230 18488 2555 18534
rect 2601 18488 2926 18534
rect 2230 18442 2266 18488
rect 2312 18442 2844 18488
rect 2890 18442 2926 18488
rect 2230 18405 2926 18442
rect 2230 18353 2269 18405
rect 2321 18353 2552 18405
rect 2604 18353 2835 18405
rect 2887 18353 2926 18405
rect 2230 18325 2555 18353
rect 2601 18325 2926 18353
rect 2230 18318 2926 18325
rect 2230 18272 2266 18318
rect 2312 18272 2844 18318
rect 2890 18272 2926 18318
rect 2230 18207 2926 18272
rect 2230 18188 2555 18207
rect 2601 18188 2926 18207
rect 2230 18136 2269 18188
rect 2321 18136 2552 18188
rect 2604 18136 2835 18188
rect 2887 18136 2926 18188
rect 2230 17970 2926 18136
rect 3259 18828 3375 18885
rect 3259 18782 3293 18828
rect 3339 18782 3375 18828
rect 3259 18658 3375 18782
rect 3259 18612 3293 18658
rect 3339 18612 3375 18658
rect 3259 18488 3375 18612
rect 3259 18442 3293 18488
rect 3339 18442 3375 18488
rect 3259 18318 3375 18442
rect 3259 18272 3293 18318
rect 3339 18272 3375 18318
rect 3259 18110 3375 18272
rect 3573 18885 3690 18886
rect 3573 18828 3689 18885
rect 3573 18782 3609 18828
rect 3655 18782 3689 18828
rect 3573 18658 3689 18782
rect 3573 18612 3609 18658
rect 3655 18612 3689 18658
rect 3573 18488 3689 18612
rect 3573 18442 3609 18488
rect 3655 18442 3689 18488
rect 3573 18318 3689 18442
rect 3573 18272 3609 18318
rect 3655 18272 3689 18318
rect 3573 18110 3689 18272
rect 4022 18860 4718 18950
rect 5045 20506 5172 20542
rect 5045 20502 5085 20506
rect 5131 20502 5172 20506
rect 5045 20450 5082 20502
rect 5134 20450 5172 20502
rect 5045 20338 5172 20450
rect 5045 20292 5085 20338
rect 5131 20292 5172 20338
rect 5045 20284 5172 20292
rect 5045 20232 5082 20284
rect 5134 20232 5172 20284
rect 5045 20171 5172 20232
rect 5045 20125 5085 20171
rect 5131 20125 5172 20171
rect 5045 20067 5172 20125
rect 5045 20015 5082 20067
rect 5134 20015 5172 20067
rect 5045 20003 5172 20015
rect 5045 19957 5085 20003
rect 5131 19957 5172 20003
rect 5045 19849 5172 19957
rect 9155 20506 9282 20542
rect 9155 20502 9196 20506
rect 9242 20502 9282 20506
rect 9155 20450 9193 20502
rect 9245 20450 9282 20502
rect 9155 20338 9282 20450
rect 9155 20292 9196 20338
rect 9242 20292 9282 20338
rect 9155 20284 9282 20292
rect 9155 20232 9193 20284
rect 9245 20232 9282 20284
rect 9155 20171 9282 20232
rect 9155 20125 9196 20171
rect 9242 20125 9282 20171
rect 9155 20067 9282 20125
rect 9155 20015 9193 20067
rect 9245 20015 9282 20067
rect 9155 20003 9282 20015
rect 9155 19957 9196 20003
rect 9242 19957 9282 20003
rect 5045 19797 5082 19849
rect 5134 19797 5172 19849
rect 5045 19789 5085 19797
rect 5131 19789 5172 19797
rect 5045 19667 5172 19789
rect 5045 19631 5085 19667
rect 5131 19631 5172 19667
rect 5045 19579 5082 19631
rect 5134 19579 5172 19631
rect 5045 19499 5172 19579
rect 5838 19837 5962 19877
rect 5838 19785 5874 19837
rect 5926 19785 5962 19837
rect 5838 19619 5962 19785
rect 5838 19567 5874 19619
rect 5926 19567 5962 19619
rect 5838 19527 5962 19567
rect 7529 19837 7653 19877
rect 7529 19785 7565 19837
rect 7617 19785 7653 19837
rect 7529 19619 7653 19785
rect 7529 19567 7565 19619
rect 7617 19567 7653 19619
rect 7529 19527 7653 19567
rect 9155 19849 9282 19957
rect 9155 19797 9193 19849
rect 9245 19797 9282 19849
rect 9155 19789 9196 19797
rect 9242 19789 9282 19797
rect 9155 19667 9282 19789
rect 9155 19631 9196 19667
rect 9242 19631 9282 19667
rect 9155 19579 9193 19631
rect 9245 19579 9282 19631
rect 5045 19453 5085 19499
rect 5131 19453 5172 19499
rect 5045 19413 5172 19453
rect 5045 19361 5082 19413
rect 5134 19361 5172 19413
rect 5045 19332 5172 19361
rect 5045 19286 5085 19332
rect 5131 19286 5172 19332
rect 5045 19196 5172 19286
rect 5045 19144 5082 19196
rect 5134 19144 5172 19196
rect 5045 19118 5085 19144
rect 5131 19118 5172 19144
rect 5045 18996 5172 19118
rect 5045 18978 5085 18996
rect 5131 18978 5172 18996
rect 5045 18926 5082 18978
rect 5134 18926 5172 18978
rect 5045 18886 5172 18926
rect 9155 19499 9282 19579
rect 9155 19453 9196 19499
rect 9242 19453 9282 19499
rect 9155 19413 9282 19453
rect 9155 19361 9193 19413
rect 9245 19361 9282 19413
rect 9155 19332 9282 19361
rect 9155 19286 9196 19332
rect 9242 19286 9282 19332
rect 9155 19196 9282 19286
rect 9155 19144 9193 19196
rect 9245 19144 9282 19196
rect 9155 19118 9196 19144
rect 9242 19118 9282 19144
rect 9155 18996 9282 19118
rect 9155 18978 9196 18996
rect 9242 18978 9282 18996
rect 9155 18926 9193 18978
rect 9245 18926 9282 18978
rect 9155 18886 9282 18926
rect 9609 20506 10305 20542
rect 9609 20460 9645 20506
rect 9691 20492 10223 20506
rect 9691 20460 9934 20492
rect 9609 20446 9934 20460
rect 9980 20460 10223 20492
rect 10269 20460 10305 20506
rect 9980 20446 10305 20460
rect 9609 20364 10305 20446
rect 9609 20338 9648 20364
rect 9609 20292 9645 20338
rect 9700 20312 9931 20364
rect 9983 20312 10214 20364
rect 10266 20338 10305 20364
rect 9691 20292 9934 20312
rect 9609 20283 9934 20292
rect 9980 20292 10223 20312
rect 10269 20292 10305 20338
rect 9980 20283 10305 20292
rect 9609 20171 10305 20283
rect 9609 20125 9645 20171
rect 9691 20166 10223 20171
rect 9691 20146 9934 20166
rect 9980 20146 10223 20166
rect 9609 20094 9648 20125
rect 9700 20094 9931 20146
rect 9983 20094 10214 20146
rect 10269 20125 10305 20171
rect 10266 20094 10305 20125
rect 9609 20003 10305 20094
rect 9609 19957 9645 20003
rect 9691 19957 9934 20003
rect 9980 19957 10223 20003
rect 10269 19957 10305 20003
rect 9609 19929 10305 19957
rect 9609 19877 9648 19929
rect 9700 19877 9931 19929
rect 9983 19877 10214 19929
rect 10266 19877 10305 19929
rect 9609 19840 10305 19877
rect 9609 19835 9934 19840
rect 9609 19789 9645 19835
rect 9691 19794 9934 19835
rect 9980 19835 10305 19840
rect 9980 19794 10223 19835
rect 9691 19789 10223 19794
rect 10269 19789 10305 19835
rect 9609 19711 10305 19789
rect 9609 19667 9648 19711
rect 9609 19621 9645 19667
rect 9700 19659 9931 19711
rect 9983 19659 10214 19711
rect 10266 19667 10305 19711
rect 9691 19630 9934 19659
rect 9980 19630 10223 19659
rect 9691 19621 10223 19630
rect 10269 19621 10305 19667
rect 9609 19513 10305 19621
rect 9609 19499 9934 19513
rect 9609 19453 9645 19499
rect 9691 19494 9934 19499
rect 9980 19499 10305 19513
rect 9980 19494 10223 19499
rect 9609 19442 9648 19453
rect 9700 19442 9931 19494
rect 9983 19442 10214 19494
rect 10269 19453 10305 19499
rect 10266 19442 10305 19453
rect 9609 19350 10305 19442
rect 9609 19332 9934 19350
rect 9609 19286 9645 19332
rect 9691 19304 9934 19332
rect 9980 19332 10305 19350
rect 9980 19304 10223 19332
rect 9691 19286 10223 19304
rect 10269 19286 10305 19332
rect 9609 19276 10305 19286
rect 9609 19224 9648 19276
rect 9700 19224 9931 19276
rect 9983 19224 10214 19276
rect 10266 19224 10305 19276
rect 9609 19187 10305 19224
rect 9609 19164 9934 19187
rect 9609 19118 9645 19164
rect 9691 19141 9934 19164
rect 9980 19164 10305 19187
rect 9980 19141 10223 19164
rect 9691 19118 10223 19141
rect 10269 19118 10305 19164
rect 9609 19058 10305 19118
rect 9609 19006 9648 19058
rect 9700 19006 9931 19058
rect 9983 19006 10214 19058
rect 10266 19006 10305 19058
rect 9609 18996 9934 19006
rect 9609 18950 9645 18996
rect 9691 18977 9934 18996
rect 9980 18996 10305 19006
rect 9980 18977 10223 18996
rect 9691 18950 10223 18977
rect 10269 18950 10305 18996
rect 5050 18885 5167 18886
rect 4022 18840 4347 18860
rect 4393 18840 4718 18860
rect 4022 18828 4061 18840
rect 4022 18782 4058 18828
rect 4113 18788 4344 18840
rect 4396 18788 4627 18840
rect 4679 18828 4718 18840
rect 4104 18782 4636 18788
rect 4682 18782 4718 18828
rect 4022 18697 4718 18782
rect 4022 18658 4347 18697
rect 4022 18612 4058 18658
rect 4104 18651 4347 18658
rect 4393 18658 4718 18697
rect 4393 18651 4636 18658
rect 4104 18623 4636 18651
rect 4022 18571 4061 18612
rect 4113 18571 4344 18623
rect 4396 18571 4627 18623
rect 4682 18612 4718 18658
rect 4679 18571 4718 18612
rect 4022 18534 4718 18571
rect 4022 18488 4347 18534
rect 4393 18488 4718 18534
rect 4022 18442 4058 18488
rect 4104 18442 4636 18488
rect 4682 18442 4718 18488
rect 4022 18405 4718 18442
rect 4022 18353 4061 18405
rect 4113 18353 4344 18405
rect 4396 18353 4627 18405
rect 4679 18353 4718 18405
rect 4022 18325 4347 18353
rect 4393 18325 4718 18353
rect 4022 18318 4718 18325
rect 4022 18272 4058 18318
rect 4104 18272 4636 18318
rect 4682 18272 4718 18318
rect 4022 18207 4718 18272
rect 4022 18188 4347 18207
rect 4393 18188 4718 18207
rect 4022 18136 4061 18188
rect 4113 18136 4344 18188
rect 4396 18136 4627 18188
rect 4679 18136 4718 18188
rect 2230 17918 2269 17970
rect 2321 17918 2552 17970
rect 2604 17918 2835 17970
rect 2887 17918 2926 17970
rect 2230 17874 2926 17918
rect 4022 17970 4718 18136
rect 5051 18828 5167 18885
rect 5051 18782 5085 18828
rect 5131 18782 5167 18828
rect 5051 18658 5167 18782
rect 5051 18612 5085 18658
rect 5131 18612 5167 18658
rect 5051 18488 5167 18612
rect 5051 18442 5085 18488
rect 5131 18442 5167 18488
rect 5051 18318 5167 18442
rect 5051 18272 5085 18318
rect 5131 18272 5167 18318
rect 5051 18110 5167 18272
rect 9160 18885 9277 18886
rect 9160 18828 9276 18885
rect 9160 18782 9196 18828
rect 9242 18782 9276 18828
rect 9160 18658 9276 18782
rect 9160 18612 9196 18658
rect 9242 18612 9276 18658
rect 9160 18488 9276 18612
rect 9160 18442 9196 18488
rect 9242 18442 9276 18488
rect 9160 18318 9276 18442
rect 9160 18272 9196 18318
rect 9242 18272 9276 18318
rect 9160 18110 9276 18272
rect 9609 18860 10305 18950
rect 10632 20506 10759 20542
rect 10632 20502 10672 20506
rect 10718 20502 10759 20506
rect 10632 20450 10669 20502
rect 10721 20450 10759 20502
rect 10632 20338 10759 20450
rect 10632 20292 10672 20338
rect 10718 20292 10759 20338
rect 10632 20284 10759 20292
rect 10632 20232 10669 20284
rect 10721 20232 10759 20284
rect 10632 20171 10759 20232
rect 10632 20125 10672 20171
rect 10718 20125 10759 20171
rect 10632 20067 10759 20125
rect 10632 20015 10669 20067
rect 10721 20015 10759 20067
rect 10632 20003 10759 20015
rect 10632 19957 10672 20003
rect 10718 19957 10759 20003
rect 10632 19849 10759 19957
rect 10632 19797 10669 19849
rect 10721 19797 10759 19849
rect 10632 19789 10672 19797
rect 10718 19789 10759 19797
rect 10632 19667 10759 19789
rect 10632 19631 10672 19667
rect 10718 19631 10759 19667
rect 10632 19579 10669 19631
rect 10721 19579 10759 19631
rect 10632 19499 10759 19579
rect 10632 19453 10672 19499
rect 10718 19453 10759 19499
rect 10632 19413 10759 19453
rect 10632 19361 10669 19413
rect 10721 19361 10759 19413
rect 10632 19332 10759 19361
rect 10632 19286 10672 19332
rect 10718 19286 10759 19332
rect 10632 19196 10759 19286
rect 10632 19144 10669 19196
rect 10721 19144 10759 19196
rect 10632 19118 10672 19144
rect 10718 19118 10759 19144
rect 10632 18996 10759 19118
rect 10632 18978 10672 18996
rect 10718 18978 10759 18996
rect 10632 18926 10669 18978
rect 10721 18926 10759 18978
rect 10632 18886 10759 18926
rect 10947 20506 11074 20542
rect 10947 20502 10988 20506
rect 11034 20502 11074 20506
rect 10947 20450 10985 20502
rect 11037 20450 11074 20502
rect 10947 20338 11074 20450
rect 10947 20292 10988 20338
rect 11034 20292 11074 20338
rect 10947 20284 11074 20292
rect 10947 20232 10985 20284
rect 11037 20232 11074 20284
rect 10947 20171 11074 20232
rect 10947 20125 10988 20171
rect 11034 20125 11074 20171
rect 10947 20067 11074 20125
rect 10947 20015 10985 20067
rect 11037 20015 11074 20067
rect 10947 20003 11074 20015
rect 10947 19957 10988 20003
rect 11034 19957 11074 20003
rect 10947 19849 11074 19957
rect 10947 19797 10985 19849
rect 11037 19797 11074 19849
rect 10947 19789 10988 19797
rect 11034 19789 11074 19797
rect 10947 19667 11074 19789
rect 10947 19631 10988 19667
rect 11034 19631 11074 19667
rect 10947 19579 10985 19631
rect 11037 19579 11074 19631
rect 10947 19499 11074 19579
rect 10947 19453 10988 19499
rect 11034 19453 11074 19499
rect 10947 19413 11074 19453
rect 10947 19361 10985 19413
rect 11037 19361 11074 19413
rect 10947 19332 11074 19361
rect 10947 19286 10988 19332
rect 11034 19286 11074 19332
rect 10947 19196 11074 19286
rect 10947 19144 10985 19196
rect 11037 19144 11074 19196
rect 10947 19118 10988 19144
rect 11034 19118 11074 19144
rect 10947 18996 11074 19118
rect 10947 18978 10988 18996
rect 11034 18978 11074 18996
rect 10947 18926 10985 18978
rect 11037 18926 11074 18978
rect 10947 18886 11074 18926
rect 11401 20506 12097 20542
rect 11401 20460 11437 20506
rect 11483 20492 12015 20506
rect 11483 20460 11726 20492
rect 11401 20446 11726 20460
rect 11772 20460 12015 20492
rect 12061 20460 12097 20506
rect 11772 20446 12097 20460
rect 11401 20364 12097 20446
rect 11401 20338 11440 20364
rect 11401 20292 11437 20338
rect 11492 20312 11723 20364
rect 11775 20312 12006 20364
rect 12058 20338 12097 20364
rect 11483 20292 11726 20312
rect 11401 20283 11726 20292
rect 11772 20292 12015 20312
rect 12061 20292 12097 20338
rect 11772 20283 12097 20292
rect 11401 20171 12097 20283
rect 11401 20125 11437 20171
rect 11483 20166 12015 20171
rect 11483 20146 11726 20166
rect 11772 20146 12015 20166
rect 11401 20094 11440 20125
rect 11492 20094 11723 20146
rect 11775 20094 12006 20146
rect 12061 20125 12097 20171
rect 12058 20094 12097 20125
rect 11401 20003 12097 20094
rect 11401 19957 11437 20003
rect 11483 19957 11726 20003
rect 11772 19957 12015 20003
rect 12061 19957 12097 20003
rect 11401 19929 12097 19957
rect 11401 19877 11440 19929
rect 11492 19877 11723 19929
rect 11775 19877 12006 19929
rect 12058 19877 12097 19929
rect 11401 19840 12097 19877
rect 11401 19835 11726 19840
rect 11401 19789 11437 19835
rect 11483 19794 11726 19835
rect 11772 19835 12097 19840
rect 11772 19794 12015 19835
rect 11483 19789 12015 19794
rect 12061 19789 12097 19835
rect 11401 19711 12097 19789
rect 11401 19667 11440 19711
rect 11401 19621 11437 19667
rect 11492 19659 11723 19711
rect 11775 19659 12006 19711
rect 12058 19667 12097 19711
rect 11483 19630 11726 19659
rect 11772 19630 12015 19659
rect 11483 19621 12015 19630
rect 12061 19621 12097 19667
rect 11401 19513 12097 19621
rect 11401 19499 11726 19513
rect 11401 19453 11437 19499
rect 11483 19494 11726 19499
rect 11772 19499 12097 19513
rect 11772 19494 12015 19499
rect 11401 19442 11440 19453
rect 11492 19442 11723 19494
rect 11775 19442 12006 19494
rect 12061 19453 12097 19499
rect 12058 19442 12097 19453
rect 11401 19350 12097 19442
rect 11401 19332 11726 19350
rect 11401 19286 11437 19332
rect 11483 19304 11726 19332
rect 11772 19332 12097 19350
rect 11772 19304 12015 19332
rect 11483 19286 12015 19304
rect 12061 19286 12097 19332
rect 11401 19276 12097 19286
rect 11401 19224 11440 19276
rect 11492 19224 11723 19276
rect 11775 19224 12006 19276
rect 12058 19224 12097 19276
rect 11401 19187 12097 19224
rect 11401 19164 11726 19187
rect 11401 19118 11437 19164
rect 11483 19141 11726 19164
rect 11772 19164 12097 19187
rect 11772 19141 12015 19164
rect 11483 19118 12015 19141
rect 12061 19118 12097 19164
rect 11401 19058 12097 19118
rect 11401 19006 11440 19058
rect 11492 19006 11723 19058
rect 11775 19006 12006 19058
rect 12058 19006 12097 19058
rect 11401 18996 11726 19006
rect 11401 18950 11437 18996
rect 11483 18977 11726 18996
rect 11772 18996 12097 19006
rect 11772 18977 12015 18996
rect 11483 18950 12015 18977
rect 12061 18950 12097 18996
rect 10637 18885 10754 18886
rect 9609 18840 9934 18860
rect 9980 18840 10305 18860
rect 9609 18828 9648 18840
rect 9609 18782 9645 18828
rect 9700 18788 9931 18840
rect 9983 18788 10214 18840
rect 10266 18828 10305 18840
rect 9691 18782 10223 18788
rect 10269 18782 10305 18828
rect 9609 18697 10305 18782
rect 9609 18658 9934 18697
rect 9609 18612 9645 18658
rect 9691 18651 9934 18658
rect 9980 18658 10305 18697
rect 9980 18651 10223 18658
rect 9691 18623 10223 18651
rect 9609 18571 9648 18612
rect 9700 18571 9931 18623
rect 9983 18571 10214 18623
rect 10269 18612 10305 18658
rect 10266 18571 10305 18612
rect 9609 18534 10305 18571
rect 9609 18488 9934 18534
rect 9980 18488 10305 18534
rect 9609 18442 9645 18488
rect 9691 18442 10223 18488
rect 10269 18442 10305 18488
rect 9609 18405 10305 18442
rect 9609 18353 9648 18405
rect 9700 18353 9931 18405
rect 9983 18353 10214 18405
rect 10266 18353 10305 18405
rect 9609 18325 9934 18353
rect 9980 18325 10305 18353
rect 9609 18318 10305 18325
rect 9609 18272 9645 18318
rect 9691 18272 10223 18318
rect 10269 18272 10305 18318
rect 9609 18207 10305 18272
rect 9609 18188 9934 18207
rect 9980 18188 10305 18207
rect 9609 18136 9648 18188
rect 9700 18136 9931 18188
rect 9983 18136 10214 18188
rect 10266 18136 10305 18188
rect 4022 17918 4061 17970
rect 4113 17918 4344 17970
rect 4396 17918 4627 17970
rect 4679 17918 4718 17970
rect 4022 17874 4718 17918
rect 9609 17970 10305 18136
rect 10638 18828 10754 18885
rect 10638 18782 10672 18828
rect 10718 18782 10754 18828
rect 10638 18658 10754 18782
rect 10638 18612 10672 18658
rect 10718 18612 10754 18658
rect 10638 18488 10754 18612
rect 10638 18442 10672 18488
rect 10718 18442 10754 18488
rect 10638 18318 10754 18442
rect 10638 18272 10672 18318
rect 10718 18272 10754 18318
rect 10638 18110 10754 18272
rect 10952 18885 11069 18886
rect 10952 18828 11068 18885
rect 10952 18782 10988 18828
rect 11034 18782 11068 18828
rect 10952 18658 11068 18782
rect 10952 18612 10988 18658
rect 11034 18612 11068 18658
rect 10952 18488 11068 18612
rect 10952 18442 10988 18488
rect 11034 18442 11068 18488
rect 10952 18318 11068 18442
rect 10952 18272 10988 18318
rect 11034 18272 11068 18318
rect 10952 18110 11068 18272
rect 11401 18860 12097 18950
rect 12424 20506 12551 20542
rect 12424 20502 12464 20506
rect 12510 20502 12551 20506
rect 12424 20450 12461 20502
rect 12513 20450 12551 20502
rect 12424 20338 12551 20450
rect 12424 20292 12464 20338
rect 12510 20292 12551 20338
rect 12424 20284 12551 20292
rect 12424 20232 12461 20284
rect 12513 20232 12551 20284
rect 12424 20171 12551 20232
rect 12424 20125 12464 20171
rect 12510 20125 12551 20171
rect 12424 20067 12551 20125
rect 12424 20015 12461 20067
rect 12513 20015 12551 20067
rect 12424 20003 12551 20015
rect 12424 19957 12464 20003
rect 12510 19957 12551 20003
rect 12424 19849 12551 19957
rect 16663 20492 16790 20529
rect 16663 20489 16704 20492
rect 16750 20489 16790 20492
rect 16663 20437 16701 20489
rect 16753 20437 16790 20489
rect 16663 20325 16790 20437
rect 17341 20492 17457 20529
rect 17341 20446 17376 20492
rect 17422 20446 17457 20492
rect 17341 20424 17457 20446
rect 18008 20492 18135 20529
rect 18008 20489 18048 20492
rect 18094 20489 18135 20492
rect 18008 20437 18045 20489
rect 18097 20437 18135 20489
rect 16663 20279 16704 20325
rect 16750 20279 16790 20325
rect 16663 20271 16790 20279
rect 16663 20219 16701 20271
rect 16753 20219 16790 20271
rect 16663 20157 16790 20219
rect 16663 20111 16704 20157
rect 16750 20111 16790 20157
rect 16663 20054 16790 20111
rect 16663 20002 16701 20054
rect 16753 20002 16790 20054
rect 16663 19989 16790 20002
rect 16663 19943 16704 19989
rect 16750 19943 16790 19989
rect 12424 19797 12461 19849
rect 12513 19797 12551 19849
rect 12424 19789 12464 19797
rect 12510 19789 12551 19797
rect 12424 19667 12551 19789
rect 12424 19631 12464 19667
rect 12510 19631 12551 19667
rect 12424 19579 12461 19631
rect 12513 19579 12551 19631
rect 12424 19499 12551 19579
rect 13217 19837 13341 19877
rect 13217 19785 13253 19837
rect 13305 19785 13341 19837
rect 13217 19619 13341 19785
rect 13217 19567 13253 19619
rect 13305 19567 13341 19619
rect 13217 19527 13341 19567
rect 14908 19837 15032 19877
rect 14908 19785 14944 19837
rect 14996 19785 15032 19837
rect 14908 19619 15032 19785
rect 14908 19567 14944 19619
rect 14996 19567 15032 19619
rect 14908 19527 15032 19567
rect 16663 19836 16790 19943
rect 16663 19784 16701 19836
rect 16753 19784 16790 19836
rect 16663 19775 16704 19784
rect 16750 19775 16790 19784
rect 16663 19654 16790 19775
rect 16663 19618 16704 19654
rect 16750 19618 16790 19654
rect 16663 19566 16701 19618
rect 16753 19566 16790 19618
rect 12424 19453 12464 19499
rect 12510 19453 12551 19499
rect 12424 19413 12551 19453
rect 12424 19361 12461 19413
rect 12513 19361 12551 19413
rect 12424 19332 12551 19361
rect 12424 19286 12464 19332
rect 12510 19286 12551 19332
rect 12424 19196 12551 19286
rect 12424 19144 12461 19196
rect 12513 19144 12551 19196
rect 12424 19118 12464 19144
rect 12510 19118 12551 19144
rect 12424 18996 12551 19118
rect 12424 18978 12464 18996
rect 12510 18978 12551 18996
rect 12424 18926 12461 18978
rect 12513 18926 12551 18978
rect 12424 18886 12551 18926
rect 16663 19486 16790 19566
rect 16663 19440 16704 19486
rect 16750 19440 16790 19486
rect 16663 19400 16790 19440
rect 16663 19348 16701 19400
rect 16753 19348 16790 19400
rect 16663 19318 16790 19348
rect 16663 19272 16704 19318
rect 16750 19272 16790 19318
rect 16663 19183 16790 19272
rect 16663 19131 16701 19183
rect 16753 19131 16790 19183
rect 16663 19104 16704 19131
rect 16750 19104 16790 19131
rect 16663 18982 16790 19104
rect 16663 18965 16704 18982
rect 16750 18965 16790 18982
rect 16663 18913 16701 18965
rect 16753 18913 16790 18965
rect 12429 18885 12546 18886
rect 11401 18840 11726 18860
rect 11772 18840 12097 18860
rect 11401 18828 11440 18840
rect 11401 18782 11437 18828
rect 11492 18788 11723 18840
rect 11775 18788 12006 18840
rect 12058 18828 12097 18840
rect 11483 18782 12015 18788
rect 12061 18782 12097 18828
rect 11401 18697 12097 18782
rect 11401 18658 11726 18697
rect 11401 18612 11437 18658
rect 11483 18651 11726 18658
rect 11772 18658 12097 18697
rect 11772 18651 12015 18658
rect 11483 18623 12015 18651
rect 11401 18571 11440 18612
rect 11492 18571 11723 18623
rect 11775 18571 12006 18623
rect 12061 18612 12097 18658
rect 12058 18571 12097 18612
rect 11401 18534 12097 18571
rect 11401 18488 11726 18534
rect 11772 18488 12097 18534
rect 11401 18442 11437 18488
rect 11483 18442 12015 18488
rect 12061 18442 12097 18488
rect 11401 18405 12097 18442
rect 11401 18353 11440 18405
rect 11492 18353 11723 18405
rect 11775 18353 12006 18405
rect 12058 18353 12097 18405
rect 11401 18325 11726 18353
rect 11772 18325 12097 18353
rect 11401 18318 12097 18325
rect 11401 18272 11437 18318
rect 11483 18272 12015 18318
rect 12061 18272 12097 18318
rect 11401 18207 12097 18272
rect 11401 18188 11726 18207
rect 11772 18188 12097 18207
rect 11401 18136 11440 18188
rect 11492 18136 11723 18188
rect 11775 18136 12006 18188
rect 12058 18136 12097 18188
rect 9609 17918 9648 17970
rect 9700 17918 9931 17970
rect 9983 17918 10214 17970
rect 10266 17918 10305 17970
rect 9609 17874 10305 17918
rect 11401 17970 12097 18136
rect 12430 18828 12546 18885
rect 16663 18873 16790 18913
rect 17335 20385 17463 20424
rect 17335 20333 17373 20385
rect 17425 20333 17463 20385
rect 17335 20325 17463 20333
rect 17335 20279 17376 20325
rect 17422 20279 17463 20325
rect 17335 20167 17463 20279
rect 17335 20115 17373 20167
rect 17425 20115 17463 20167
rect 17335 20111 17376 20115
rect 17422 20111 17463 20115
rect 17335 19989 17463 20111
rect 17335 19950 17376 19989
rect 17422 19950 17463 19989
rect 17335 19898 17373 19950
rect 17425 19898 17463 19950
rect 17335 19821 17463 19898
rect 17335 19775 17376 19821
rect 17422 19775 17463 19821
rect 17335 19732 17463 19775
rect 17335 19680 17373 19732
rect 17425 19680 17463 19732
rect 17335 19654 17463 19680
rect 17335 19608 17376 19654
rect 17422 19608 17463 19654
rect 17335 19514 17463 19608
rect 17335 19462 17373 19514
rect 17425 19462 17463 19514
rect 17335 19440 17376 19462
rect 17422 19440 17463 19462
rect 17335 19318 17463 19440
rect 17335 19297 17376 19318
rect 17422 19297 17463 19318
rect 17335 19245 17373 19297
rect 17425 19245 17463 19297
rect 17335 19150 17463 19245
rect 17335 19104 17376 19150
rect 17422 19104 17463 19150
rect 17335 19079 17463 19104
rect 17335 19027 17373 19079
rect 17425 19027 17463 19079
rect 17335 18982 17463 19027
rect 17335 18936 17376 18982
rect 17422 18936 17463 18982
rect 16669 18872 16785 18873
rect 12430 18782 12464 18828
rect 12510 18782 12546 18828
rect 12430 18658 12546 18782
rect 12430 18612 12464 18658
rect 12510 18612 12546 18658
rect 12430 18488 12546 18612
rect 12430 18442 12464 18488
rect 12510 18442 12546 18488
rect 12430 18318 12546 18442
rect 12430 18272 12464 18318
rect 12510 18272 12546 18318
rect 12430 18110 12546 18272
rect 16670 18815 16785 18872
rect 16670 18769 16704 18815
rect 16750 18769 16785 18815
rect 16670 18645 16785 18769
rect 16670 18599 16704 18645
rect 16750 18599 16785 18645
rect 16670 18475 16785 18599
rect 16670 18429 16704 18475
rect 16750 18429 16785 18475
rect 16670 18305 16785 18429
rect 16670 18259 16704 18305
rect 16750 18259 16785 18305
rect 16670 18135 16785 18259
rect 16670 18089 16704 18135
rect 16750 18089 16785 18135
rect 16670 18052 16785 18089
rect 17335 18861 17463 18936
rect 18008 20325 18135 20437
rect 18008 20279 18048 20325
rect 18094 20279 18135 20325
rect 18008 20271 18135 20279
rect 18008 20219 18045 20271
rect 18097 20219 18135 20271
rect 18008 20157 18135 20219
rect 18008 20111 18048 20157
rect 18094 20111 18135 20157
rect 18008 20054 18135 20111
rect 18008 20002 18045 20054
rect 18097 20002 18135 20054
rect 18008 19989 18135 20002
rect 18008 19943 18048 19989
rect 18094 19943 18135 19989
rect 18008 19836 18135 19943
rect 18008 19784 18045 19836
rect 18097 19784 18135 19836
rect 18008 19775 18048 19784
rect 18094 19775 18135 19784
rect 18008 19654 18135 19775
rect 18008 19618 18048 19654
rect 18094 19618 18135 19654
rect 18008 19566 18045 19618
rect 18097 19566 18135 19618
rect 18008 19486 18135 19566
rect 18008 19440 18048 19486
rect 18094 19440 18135 19486
rect 18008 19400 18135 19440
rect 18008 19348 18045 19400
rect 18097 19348 18135 19400
rect 18008 19318 18135 19348
rect 18008 19272 18048 19318
rect 18094 19272 18135 19318
rect 18008 19183 18135 19272
rect 18008 19131 18045 19183
rect 18097 19131 18135 19183
rect 18008 19104 18048 19131
rect 18094 19104 18135 19131
rect 18008 18982 18135 19104
rect 18008 18965 18048 18982
rect 18094 18965 18135 18982
rect 18008 18913 18045 18965
rect 18097 18913 18135 18965
rect 18008 18873 18135 18913
rect 18297 20492 18424 20529
rect 18297 20489 18338 20492
rect 18384 20489 18424 20492
rect 18297 20437 18335 20489
rect 18387 20437 18424 20489
rect 18297 20325 18424 20437
rect 18975 20492 19091 20529
rect 18975 20446 19010 20492
rect 19056 20446 19091 20492
rect 18975 20424 19091 20446
rect 19642 20492 19769 20529
rect 19642 20489 19682 20492
rect 19728 20489 19769 20492
rect 19642 20437 19679 20489
rect 19731 20437 19769 20489
rect 18297 20279 18338 20325
rect 18384 20279 18424 20325
rect 18297 20271 18424 20279
rect 18297 20219 18335 20271
rect 18387 20219 18424 20271
rect 18297 20157 18424 20219
rect 18297 20111 18338 20157
rect 18384 20111 18424 20157
rect 18297 20054 18424 20111
rect 18297 20002 18335 20054
rect 18387 20002 18424 20054
rect 18297 19989 18424 20002
rect 18297 19943 18338 19989
rect 18384 19943 18424 19989
rect 18297 19836 18424 19943
rect 18297 19784 18335 19836
rect 18387 19784 18424 19836
rect 18297 19775 18338 19784
rect 18384 19775 18424 19784
rect 18297 19654 18424 19775
rect 18297 19618 18338 19654
rect 18384 19618 18424 19654
rect 18297 19566 18335 19618
rect 18387 19566 18424 19618
rect 18297 19486 18424 19566
rect 18297 19440 18338 19486
rect 18384 19440 18424 19486
rect 18297 19400 18424 19440
rect 18297 19348 18335 19400
rect 18387 19348 18424 19400
rect 18297 19318 18424 19348
rect 18297 19272 18338 19318
rect 18384 19272 18424 19318
rect 18297 19183 18424 19272
rect 18297 19131 18335 19183
rect 18387 19131 18424 19183
rect 18297 19104 18338 19131
rect 18384 19104 18424 19131
rect 18297 18982 18424 19104
rect 18297 18965 18338 18982
rect 18384 18965 18424 18982
rect 18297 18913 18335 18965
rect 18387 18913 18424 18965
rect 18297 18873 18424 18913
rect 18969 20385 19097 20424
rect 18969 20333 19007 20385
rect 19059 20333 19097 20385
rect 18969 20325 19097 20333
rect 18969 20279 19010 20325
rect 19056 20279 19097 20325
rect 18969 20167 19097 20279
rect 18969 20115 19007 20167
rect 19059 20115 19097 20167
rect 18969 20111 19010 20115
rect 19056 20111 19097 20115
rect 18969 19989 19097 20111
rect 18969 19950 19010 19989
rect 19056 19950 19097 19989
rect 18969 19898 19007 19950
rect 19059 19898 19097 19950
rect 18969 19821 19097 19898
rect 18969 19775 19010 19821
rect 19056 19775 19097 19821
rect 18969 19732 19097 19775
rect 18969 19680 19007 19732
rect 19059 19680 19097 19732
rect 18969 19654 19097 19680
rect 18969 19608 19010 19654
rect 19056 19608 19097 19654
rect 18969 19514 19097 19608
rect 18969 19462 19007 19514
rect 19059 19462 19097 19514
rect 18969 19440 19010 19462
rect 19056 19440 19097 19462
rect 18969 19318 19097 19440
rect 18969 19297 19010 19318
rect 19056 19297 19097 19318
rect 18969 19245 19007 19297
rect 19059 19245 19097 19297
rect 18969 19150 19097 19245
rect 18969 19104 19010 19150
rect 19056 19104 19097 19150
rect 18969 19079 19097 19104
rect 18969 19027 19007 19079
rect 19059 19027 19097 19079
rect 18969 18982 19097 19027
rect 18969 18936 19010 18982
rect 19056 18936 19097 18982
rect 17335 18809 17373 18861
rect 17425 18809 17463 18861
rect 17335 18769 17376 18809
rect 17422 18769 17463 18809
rect 17335 18645 17463 18769
rect 17335 18644 17376 18645
rect 17422 18644 17463 18645
rect 17335 18592 17373 18644
rect 17425 18592 17463 18644
rect 17335 18475 17463 18592
rect 17335 18429 17376 18475
rect 17422 18429 17463 18475
rect 17335 18426 17463 18429
rect 17335 18374 17373 18426
rect 17425 18374 17463 18426
rect 17335 18305 17463 18374
rect 17335 18259 17376 18305
rect 17422 18259 17463 18305
rect 17335 18208 17463 18259
rect 17335 18156 17373 18208
rect 17425 18156 17463 18208
rect 17335 18135 17463 18156
rect 17335 18089 17376 18135
rect 17422 18089 17463 18135
rect 11401 17918 11440 17970
rect 11492 17918 11723 17970
rect 11775 17918 12006 17970
rect 12058 17918 12097 17970
rect 17335 17991 17463 18089
rect 18013 18872 18129 18873
rect 18303 18872 18419 18873
rect 18013 18815 18128 18872
rect 18013 18769 18048 18815
rect 18094 18769 18128 18815
rect 18013 18645 18128 18769
rect 18013 18599 18048 18645
rect 18094 18599 18128 18645
rect 18013 18475 18128 18599
rect 18013 18429 18048 18475
rect 18094 18429 18128 18475
rect 18013 18305 18128 18429
rect 18013 18259 18048 18305
rect 18094 18259 18128 18305
rect 18013 18135 18128 18259
rect 18013 18089 18048 18135
rect 18094 18089 18128 18135
rect 18013 18052 18128 18089
rect 18304 18815 18419 18872
rect 18304 18769 18338 18815
rect 18384 18769 18419 18815
rect 18304 18645 18419 18769
rect 18304 18599 18338 18645
rect 18384 18599 18419 18645
rect 18304 18475 18419 18599
rect 18304 18429 18338 18475
rect 18384 18429 18419 18475
rect 18304 18305 18419 18429
rect 18304 18259 18338 18305
rect 18384 18259 18419 18305
rect 18304 18135 18419 18259
rect 18304 18089 18338 18135
rect 18384 18089 18419 18135
rect 18304 18052 18419 18089
rect 18969 18861 19097 18936
rect 19642 20325 19769 20437
rect 19642 20279 19682 20325
rect 19728 20279 19769 20325
rect 19642 20271 19769 20279
rect 19642 20219 19679 20271
rect 19731 20219 19769 20271
rect 19642 20157 19769 20219
rect 19642 20111 19682 20157
rect 19728 20111 19769 20157
rect 19642 20054 19769 20111
rect 19642 20002 19679 20054
rect 19731 20002 19769 20054
rect 19642 19989 19769 20002
rect 19642 19943 19682 19989
rect 19728 19943 19769 19989
rect 19642 19836 19769 19943
rect 19642 19784 19679 19836
rect 19731 19784 19769 19836
rect 19642 19775 19682 19784
rect 19728 19775 19769 19784
rect 19642 19654 19769 19775
rect 19642 19618 19682 19654
rect 19728 19618 19769 19654
rect 19642 19566 19679 19618
rect 19731 19566 19769 19618
rect 19642 19486 19769 19566
rect 19642 19440 19682 19486
rect 19728 19440 19769 19486
rect 19642 19400 19769 19440
rect 19642 19348 19679 19400
rect 19731 19348 19769 19400
rect 19642 19318 19769 19348
rect 19642 19272 19682 19318
rect 19728 19272 19769 19318
rect 19642 19183 19769 19272
rect 19642 19131 19679 19183
rect 19731 19131 19769 19183
rect 19642 19104 19682 19131
rect 19728 19104 19769 19131
rect 19642 18982 19769 19104
rect 19642 18965 19682 18982
rect 19728 18965 19769 18982
rect 19642 18913 19679 18965
rect 19731 18913 19769 18965
rect 19642 18873 19769 18913
rect 19930 20492 20057 20529
rect 19930 20489 19971 20492
rect 20017 20489 20057 20492
rect 19930 20437 19968 20489
rect 20020 20437 20057 20489
rect 19930 20325 20057 20437
rect 20608 20492 20724 20529
rect 20608 20446 20643 20492
rect 20689 20446 20724 20492
rect 20608 20424 20724 20446
rect 21275 20492 21402 20529
rect 21275 20489 21315 20492
rect 21361 20489 21402 20492
rect 21275 20437 21312 20489
rect 21364 20437 21402 20489
rect 19930 20279 19971 20325
rect 20017 20279 20057 20325
rect 19930 20271 20057 20279
rect 19930 20219 19968 20271
rect 20020 20219 20057 20271
rect 19930 20157 20057 20219
rect 19930 20111 19971 20157
rect 20017 20111 20057 20157
rect 19930 20054 20057 20111
rect 19930 20002 19968 20054
rect 20020 20002 20057 20054
rect 19930 19989 20057 20002
rect 19930 19943 19971 19989
rect 20017 19943 20057 19989
rect 19930 19836 20057 19943
rect 19930 19784 19968 19836
rect 20020 19784 20057 19836
rect 19930 19775 19971 19784
rect 20017 19775 20057 19784
rect 19930 19654 20057 19775
rect 19930 19618 19971 19654
rect 20017 19618 20057 19654
rect 19930 19566 19968 19618
rect 20020 19566 20057 19618
rect 19930 19486 20057 19566
rect 19930 19440 19971 19486
rect 20017 19440 20057 19486
rect 19930 19400 20057 19440
rect 19930 19348 19968 19400
rect 20020 19348 20057 19400
rect 19930 19318 20057 19348
rect 19930 19272 19971 19318
rect 20017 19272 20057 19318
rect 19930 19183 20057 19272
rect 19930 19131 19968 19183
rect 20020 19131 20057 19183
rect 19930 19104 19971 19131
rect 20017 19104 20057 19131
rect 19930 18982 20057 19104
rect 19930 18965 19971 18982
rect 20017 18965 20057 18982
rect 19930 18913 19968 18965
rect 20020 18913 20057 18965
rect 19930 18873 20057 18913
rect 20602 20385 20730 20424
rect 20602 20333 20640 20385
rect 20692 20333 20730 20385
rect 20602 20325 20730 20333
rect 20602 20279 20643 20325
rect 20689 20279 20730 20325
rect 20602 20167 20730 20279
rect 20602 20115 20640 20167
rect 20692 20115 20730 20167
rect 20602 20111 20643 20115
rect 20689 20111 20730 20115
rect 20602 19989 20730 20111
rect 20602 19950 20643 19989
rect 20689 19950 20730 19989
rect 20602 19898 20640 19950
rect 20692 19898 20730 19950
rect 20602 19821 20730 19898
rect 20602 19775 20643 19821
rect 20689 19775 20730 19821
rect 20602 19732 20730 19775
rect 20602 19680 20640 19732
rect 20692 19680 20730 19732
rect 20602 19654 20730 19680
rect 20602 19608 20643 19654
rect 20689 19608 20730 19654
rect 20602 19514 20730 19608
rect 20602 19462 20640 19514
rect 20692 19462 20730 19514
rect 20602 19440 20643 19462
rect 20689 19440 20730 19462
rect 20602 19318 20730 19440
rect 20602 19297 20643 19318
rect 20689 19297 20730 19318
rect 20602 19245 20640 19297
rect 20692 19245 20730 19297
rect 20602 19150 20730 19245
rect 20602 19104 20643 19150
rect 20689 19104 20730 19150
rect 20602 19079 20730 19104
rect 20602 19027 20640 19079
rect 20692 19027 20730 19079
rect 20602 18982 20730 19027
rect 20602 18936 20643 18982
rect 20689 18936 20730 18982
rect 18969 18809 19007 18861
rect 19059 18809 19097 18861
rect 18969 18769 19010 18809
rect 19056 18769 19097 18809
rect 18969 18645 19097 18769
rect 18969 18644 19010 18645
rect 19056 18644 19097 18645
rect 18969 18592 19007 18644
rect 19059 18592 19097 18644
rect 18969 18475 19097 18592
rect 18969 18429 19010 18475
rect 19056 18429 19097 18475
rect 18969 18426 19097 18429
rect 18969 18374 19007 18426
rect 19059 18374 19097 18426
rect 18969 18305 19097 18374
rect 18969 18259 19010 18305
rect 19056 18259 19097 18305
rect 18969 18208 19097 18259
rect 18969 18156 19007 18208
rect 19059 18156 19097 18208
rect 18969 18135 19097 18156
rect 18969 18089 19010 18135
rect 19056 18089 19097 18135
rect 17335 17962 17373 17991
rect 11401 17874 12097 17918
rect 16581 17939 17373 17962
rect 17425 17962 17463 17991
rect 18969 17991 19097 18089
rect 19647 18872 19763 18873
rect 19936 18872 20052 18873
rect 19647 18815 19762 18872
rect 19647 18769 19682 18815
rect 19728 18769 19762 18815
rect 19647 18645 19762 18769
rect 19647 18599 19682 18645
rect 19728 18599 19762 18645
rect 19647 18475 19762 18599
rect 19647 18429 19682 18475
rect 19728 18429 19762 18475
rect 19647 18305 19762 18429
rect 19647 18259 19682 18305
rect 19728 18259 19762 18305
rect 19647 18135 19762 18259
rect 19647 18089 19682 18135
rect 19728 18089 19762 18135
rect 19647 18052 19762 18089
rect 19937 18815 20052 18872
rect 19937 18769 19971 18815
rect 20017 18769 20052 18815
rect 19937 18645 20052 18769
rect 19937 18599 19971 18645
rect 20017 18599 20052 18645
rect 19937 18475 20052 18599
rect 19937 18429 19971 18475
rect 20017 18429 20052 18475
rect 19937 18305 20052 18429
rect 19937 18259 19971 18305
rect 20017 18259 20052 18305
rect 19937 18135 20052 18259
rect 19937 18089 19971 18135
rect 20017 18089 20052 18135
rect 19937 18052 20052 18089
rect 20602 18861 20730 18936
rect 21275 20325 21402 20437
rect 21275 20279 21315 20325
rect 21361 20279 21402 20325
rect 21275 20271 21402 20279
rect 21275 20219 21312 20271
rect 21364 20219 21402 20271
rect 21275 20157 21402 20219
rect 21275 20111 21315 20157
rect 21361 20111 21402 20157
rect 21275 20054 21402 20111
rect 21275 20002 21312 20054
rect 21364 20002 21402 20054
rect 21275 19989 21402 20002
rect 21275 19943 21315 19989
rect 21361 19943 21402 19989
rect 21275 19836 21402 19943
rect 21275 19784 21312 19836
rect 21364 19784 21402 19836
rect 21275 19775 21315 19784
rect 21361 19775 21402 19784
rect 21275 19654 21402 19775
rect 21275 19618 21315 19654
rect 21361 19618 21402 19654
rect 21275 19566 21312 19618
rect 21364 19566 21402 19618
rect 21275 19486 21402 19566
rect 21275 19440 21315 19486
rect 21361 19440 21402 19486
rect 21275 19400 21402 19440
rect 21275 19348 21312 19400
rect 21364 19348 21402 19400
rect 21275 19318 21402 19348
rect 21275 19272 21315 19318
rect 21361 19272 21402 19318
rect 21275 19183 21402 19272
rect 21275 19131 21312 19183
rect 21364 19131 21402 19183
rect 21275 19104 21315 19131
rect 21361 19104 21402 19131
rect 21275 18982 21402 19104
rect 21275 18965 21315 18982
rect 21361 18965 21402 18982
rect 21275 18913 21312 18965
rect 21364 18913 21402 18965
rect 21275 18873 21402 18913
rect 21564 20492 21691 20529
rect 21564 20489 21605 20492
rect 21651 20489 21691 20492
rect 21564 20437 21602 20489
rect 21654 20437 21691 20489
rect 21564 20325 21691 20437
rect 22242 20492 22358 20529
rect 22242 20446 22277 20492
rect 22323 20446 22358 20492
rect 22242 20424 22358 20446
rect 22909 20492 23036 20529
rect 22909 20489 22949 20492
rect 22995 20489 23036 20492
rect 22909 20437 22946 20489
rect 22998 20437 23036 20489
rect 21564 20279 21605 20325
rect 21651 20279 21691 20325
rect 21564 20271 21691 20279
rect 21564 20219 21602 20271
rect 21654 20219 21691 20271
rect 21564 20157 21691 20219
rect 21564 20111 21605 20157
rect 21651 20111 21691 20157
rect 21564 20054 21691 20111
rect 21564 20002 21602 20054
rect 21654 20002 21691 20054
rect 21564 19989 21691 20002
rect 21564 19943 21605 19989
rect 21651 19943 21691 19989
rect 21564 19836 21691 19943
rect 21564 19784 21602 19836
rect 21654 19784 21691 19836
rect 21564 19775 21605 19784
rect 21651 19775 21691 19784
rect 21564 19654 21691 19775
rect 21564 19618 21605 19654
rect 21651 19618 21691 19654
rect 21564 19566 21602 19618
rect 21654 19566 21691 19618
rect 21564 19486 21691 19566
rect 21564 19440 21605 19486
rect 21651 19440 21691 19486
rect 21564 19400 21691 19440
rect 21564 19348 21602 19400
rect 21654 19348 21691 19400
rect 21564 19318 21691 19348
rect 21564 19272 21605 19318
rect 21651 19272 21691 19318
rect 21564 19183 21691 19272
rect 21564 19131 21602 19183
rect 21654 19131 21691 19183
rect 21564 19104 21605 19131
rect 21651 19104 21691 19131
rect 21564 18982 21691 19104
rect 21564 18965 21605 18982
rect 21651 18965 21691 18982
rect 21564 18913 21602 18965
rect 21654 18913 21691 18965
rect 21564 18873 21691 18913
rect 22236 20385 22364 20424
rect 22236 20333 22274 20385
rect 22326 20333 22364 20385
rect 22236 20325 22364 20333
rect 22236 20279 22277 20325
rect 22323 20279 22364 20325
rect 22236 20167 22364 20279
rect 22236 20115 22274 20167
rect 22326 20115 22364 20167
rect 22236 20111 22277 20115
rect 22323 20111 22364 20115
rect 22236 19989 22364 20111
rect 22236 19950 22277 19989
rect 22323 19950 22364 19989
rect 22236 19898 22274 19950
rect 22326 19898 22364 19950
rect 22236 19821 22364 19898
rect 22236 19775 22277 19821
rect 22323 19775 22364 19821
rect 22236 19732 22364 19775
rect 22236 19680 22274 19732
rect 22326 19680 22364 19732
rect 22236 19654 22364 19680
rect 22236 19608 22277 19654
rect 22323 19608 22364 19654
rect 22236 19514 22364 19608
rect 22236 19462 22274 19514
rect 22326 19462 22364 19514
rect 22236 19440 22277 19462
rect 22323 19440 22364 19462
rect 22236 19318 22364 19440
rect 22236 19297 22277 19318
rect 22323 19297 22364 19318
rect 22236 19245 22274 19297
rect 22326 19245 22364 19297
rect 22236 19150 22364 19245
rect 22236 19104 22277 19150
rect 22323 19104 22364 19150
rect 22236 19079 22364 19104
rect 22236 19027 22274 19079
rect 22326 19027 22364 19079
rect 22236 18982 22364 19027
rect 22236 18936 22277 18982
rect 22323 18936 22364 18982
rect 20602 18809 20640 18861
rect 20692 18809 20730 18861
rect 20602 18769 20643 18809
rect 20689 18769 20730 18809
rect 20602 18645 20730 18769
rect 20602 18644 20643 18645
rect 20689 18644 20730 18645
rect 20602 18592 20640 18644
rect 20692 18592 20730 18644
rect 20602 18475 20730 18592
rect 20602 18429 20643 18475
rect 20689 18429 20730 18475
rect 20602 18426 20730 18429
rect 20602 18374 20640 18426
rect 20692 18374 20730 18426
rect 20602 18305 20730 18374
rect 20602 18259 20643 18305
rect 20689 18259 20730 18305
rect 20602 18208 20730 18259
rect 20602 18156 20640 18208
rect 20692 18156 20730 18208
rect 20602 18135 20730 18156
rect 20602 18089 20643 18135
rect 20689 18089 20730 18135
rect 18969 17962 19007 17991
rect 17425 17939 19007 17962
rect 19059 17962 19097 17991
rect 20602 17991 20730 18089
rect 21280 18872 21396 18873
rect 21570 18872 21686 18873
rect 21280 18815 21395 18872
rect 21280 18769 21315 18815
rect 21361 18769 21395 18815
rect 21280 18645 21395 18769
rect 21280 18599 21315 18645
rect 21361 18599 21395 18645
rect 21280 18475 21395 18599
rect 21280 18429 21315 18475
rect 21361 18429 21395 18475
rect 21280 18305 21395 18429
rect 21280 18259 21315 18305
rect 21361 18259 21395 18305
rect 21280 18135 21395 18259
rect 21280 18089 21315 18135
rect 21361 18089 21395 18135
rect 21280 18052 21395 18089
rect 21571 18815 21686 18872
rect 21571 18769 21605 18815
rect 21651 18769 21686 18815
rect 21571 18645 21686 18769
rect 21571 18599 21605 18645
rect 21651 18599 21686 18645
rect 21571 18475 21686 18599
rect 21571 18429 21605 18475
rect 21651 18429 21686 18475
rect 21571 18305 21686 18429
rect 21571 18259 21605 18305
rect 21651 18259 21686 18305
rect 21571 18135 21686 18259
rect 21571 18089 21605 18135
rect 21651 18089 21686 18135
rect 21571 18052 21686 18089
rect 22236 18861 22364 18936
rect 22909 20325 23036 20437
rect 22909 20279 22949 20325
rect 22995 20279 23036 20325
rect 22909 20271 23036 20279
rect 22909 20219 22946 20271
rect 22998 20219 23036 20271
rect 22909 20157 23036 20219
rect 22909 20111 22949 20157
rect 22995 20111 23036 20157
rect 22909 20054 23036 20111
rect 22909 20002 22946 20054
rect 22998 20002 23036 20054
rect 22909 19989 23036 20002
rect 22909 19943 22949 19989
rect 22995 19943 23036 19989
rect 22909 19836 23036 19943
rect 22909 19784 22946 19836
rect 22998 19784 23036 19836
rect 22909 19775 22949 19784
rect 22995 19775 23036 19784
rect 22909 19654 23036 19775
rect 22909 19618 22949 19654
rect 22995 19618 23036 19654
rect 22909 19566 22946 19618
rect 22998 19566 23036 19618
rect 22909 19486 23036 19566
rect 23703 19837 23827 19877
rect 23703 19785 23739 19837
rect 23791 19785 23827 19837
rect 23703 19619 23827 19785
rect 23703 19567 23739 19619
rect 23791 19567 23827 19619
rect 23703 19527 23827 19567
rect 25393 19837 25517 19877
rect 25393 19785 25429 19837
rect 25481 19785 25517 19837
rect 25393 19619 25517 19785
rect 25393 19567 25429 19619
rect 25481 19567 25517 19619
rect 25393 19527 25517 19567
rect 27084 19837 27208 19877
rect 27084 19785 27120 19837
rect 27172 19785 27208 19837
rect 27084 19619 27208 19785
rect 27084 19567 27120 19619
rect 27172 19567 27208 19619
rect 27084 19527 27208 19567
rect 22909 19440 22949 19486
rect 22995 19440 23036 19486
rect 22909 19400 23036 19440
rect 22909 19348 22946 19400
rect 22998 19348 23036 19400
rect 22909 19318 23036 19348
rect 22909 19272 22949 19318
rect 22995 19272 23036 19318
rect 22909 19183 23036 19272
rect 22909 19131 22946 19183
rect 22998 19131 23036 19183
rect 22909 19104 22949 19131
rect 22995 19104 23036 19131
rect 22909 18982 23036 19104
rect 22909 18965 22949 18982
rect 22995 18965 23036 18982
rect 22909 18913 22946 18965
rect 22998 18913 23036 18965
rect 22909 18873 23036 18913
rect 22236 18809 22274 18861
rect 22326 18809 22364 18861
rect 22236 18769 22277 18809
rect 22323 18769 22364 18809
rect 22236 18645 22364 18769
rect 22236 18644 22277 18645
rect 22323 18644 22364 18645
rect 22236 18592 22274 18644
rect 22326 18592 22364 18644
rect 22236 18475 22364 18592
rect 22236 18429 22277 18475
rect 22323 18429 22364 18475
rect 22236 18426 22364 18429
rect 22236 18374 22274 18426
rect 22326 18374 22364 18426
rect 22236 18305 22364 18374
rect 22236 18259 22277 18305
rect 22323 18259 22364 18305
rect 22236 18208 22364 18259
rect 22236 18156 22274 18208
rect 22326 18156 22364 18208
rect 22236 18135 22364 18156
rect 22236 18089 22277 18135
rect 22323 18089 22364 18135
rect 20602 17962 20640 17991
rect 19059 17939 20640 17962
rect 20692 17962 20730 17991
rect 22236 17991 22364 18089
rect 22914 18872 23030 18873
rect 22914 18815 23029 18872
rect 22914 18769 22949 18815
rect 22995 18769 23029 18815
rect 22914 18645 23029 18769
rect 22914 18599 22949 18645
rect 22995 18599 23029 18645
rect 22914 18475 23029 18599
rect 22914 18429 22949 18475
rect 22995 18429 23029 18475
rect 22914 18305 23029 18429
rect 22914 18259 22949 18305
rect 22995 18259 23029 18305
rect 22914 18135 23029 18259
rect 22914 18089 22949 18135
rect 22995 18089 23029 18135
rect 22914 18052 23029 18089
rect 22236 17962 22274 17991
rect 20692 17939 22274 17962
rect 22326 17962 22364 17991
rect 22326 17939 23118 17962
rect 1681 17833 5267 17874
rect 1681 17787 1763 17833
rect 1809 17787 1921 17833
rect 1967 17787 2079 17833
rect 2125 17787 2237 17833
rect 2283 17787 2395 17833
rect 2441 17787 2715 17833
rect 2761 17787 2873 17833
rect 2919 17787 3031 17833
rect 3077 17787 3189 17833
rect 3235 17787 3347 17833
rect 3393 17787 3555 17833
rect 3601 17787 3713 17833
rect 3759 17787 3871 17833
rect 3917 17787 4029 17833
rect 4075 17787 4187 17833
rect 4233 17787 4507 17833
rect 4553 17787 4665 17833
rect 4711 17787 4823 17833
rect 4869 17787 4981 17833
rect 5027 17787 5139 17833
rect 5185 17787 5267 17833
rect 9060 17833 12646 17874
rect 1681 17745 5267 17787
rect 6826 17625 6956 17826
rect 765 17491 6956 17625
rect 765 10724 894 17491
rect 8530 17398 8660 17813
rect 9060 17787 9142 17833
rect 9188 17787 9300 17833
rect 9346 17787 9458 17833
rect 9504 17787 9616 17833
rect 9662 17787 9774 17833
rect 9820 17787 10094 17833
rect 10140 17787 10252 17833
rect 10298 17787 10410 17833
rect 10456 17787 10568 17833
rect 10614 17787 10726 17833
rect 10772 17787 10934 17833
rect 10980 17787 11092 17833
rect 11138 17787 11250 17833
rect 11296 17787 11408 17833
rect 11454 17787 11566 17833
rect 11612 17787 11886 17833
rect 11932 17787 12044 17833
rect 12090 17787 12202 17833
rect 12248 17787 12360 17833
rect 12406 17787 12518 17833
rect 12564 17787 12646 17833
rect 9060 17745 12646 17787
rect 1007 17264 8660 17398
rect 1007 11101 1136 17264
rect 14218 17171 14347 17797
rect 1248 17038 14347 17171
rect 15909 17248 16038 17874
rect 16581 17773 23118 17939
rect 16581 17767 17373 17773
rect 16581 17721 16812 17767
rect 16858 17721 16970 17767
rect 17016 17721 17128 17767
rect 17174 17721 17286 17767
rect 17332 17721 17373 17767
rect 17425 17767 19007 17773
rect 17425 17721 17466 17767
rect 17512 17721 17624 17767
rect 17670 17721 17782 17767
rect 17828 17721 17940 17767
rect 17986 17721 18446 17767
rect 18492 17721 18604 17767
rect 18650 17721 18762 17767
rect 18808 17721 18920 17767
rect 18966 17721 19007 17767
rect 19059 17767 20640 17773
rect 19059 17721 19100 17767
rect 19146 17721 19258 17767
rect 19304 17721 19416 17767
rect 19462 17721 19574 17767
rect 19620 17721 20079 17767
rect 20125 17721 20237 17767
rect 20283 17721 20395 17767
rect 20441 17721 20553 17767
rect 20599 17721 20640 17767
rect 20692 17767 22274 17773
rect 20692 17721 20733 17767
rect 20779 17721 20891 17767
rect 20937 17721 21049 17767
rect 21095 17721 21207 17767
rect 21253 17721 21713 17767
rect 21759 17721 21871 17767
rect 21917 17721 22029 17767
rect 22075 17721 22187 17767
rect 22233 17721 22274 17767
rect 22326 17767 23118 17773
rect 22326 17721 22367 17767
rect 22413 17721 22525 17767
rect 22571 17721 22683 17767
rect 22729 17721 22841 17767
rect 22887 17721 23118 17767
rect 16581 17671 23118 17721
rect 24704 17475 24833 17890
rect 26395 17702 26524 17904
rect 28070 17795 28861 17928
rect 26395 17568 28619 17702
rect 24704 17342 28378 17475
rect 15909 17115 28136 17248
rect 1248 11393 1377 17038
rect 1953 16902 20175 16924
rect 1953 16850 1992 16902
rect 2044 16887 2664 16902
rect 2716 16887 3112 16902
rect 3164 16887 3784 16902
rect 3836 16887 4232 16902
rect 4284 16887 4904 16902
rect 1953 16841 2012 16850
rect 2058 16841 2171 16887
rect 2217 16841 2329 16887
rect 2375 16841 2487 16887
rect 2533 16841 2645 16887
rect 2716 16850 2803 16887
rect 2691 16841 2803 16850
rect 2849 16841 2961 16887
rect 3007 16850 3112 16887
rect 3007 16841 3119 16850
rect 3165 16841 3277 16887
rect 3323 16841 3435 16887
rect 3481 16841 3594 16887
rect 3640 16841 3752 16887
rect 3836 16850 3910 16887
rect 3798 16841 3910 16850
rect 3956 16841 4068 16887
rect 4114 16841 4226 16887
rect 4284 16850 4384 16887
rect 4272 16841 4384 16850
rect 4430 16841 4542 16887
rect 4588 16841 4700 16887
rect 4746 16841 4858 16887
rect 4956 16887 5352 16902
rect 5404 16887 6024 16902
rect 4956 16850 5017 16887
rect 4904 16841 5017 16850
rect 5063 16841 5175 16887
rect 5221 16841 5333 16887
rect 5404 16850 5491 16887
rect 5379 16841 5491 16850
rect 5537 16841 5649 16887
rect 5695 16841 5807 16887
rect 5853 16841 5965 16887
rect 6011 16850 6024 16887
rect 6076 16887 6472 16902
rect 6524 16887 7144 16902
rect 6076 16850 6123 16887
rect 6011 16841 6123 16850
rect 6169 16841 6282 16887
rect 6328 16841 6440 16887
rect 6524 16850 6598 16887
rect 6486 16841 6598 16850
rect 6644 16841 6756 16887
rect 6802 16841 6914 16887
rect 6960 16841 7072 16887
rect 7118 16850 7144 16887
rect 7196 16887 7592 16902
rect 7196 16850 7230 16887
rect 7118 16841 7230 16850
rect 7276 16841 7388 16887
rect 7434 16841 7546 16887
rect 7644 16887 8264 16902
rect 7644 16850 7705 16887
rect 7592 16841 7705 16850
rect 7751 16841 7863 16887
rect 7909 16841 8021 16887
rect 8067 16841 8179 16887
rect 8225 16850 8264 16887
rect 8316 16887 8712 16902
rect 8316 16850 8337 16887
rect 8225 16841 8337 16850
rect 8383 16841 8495 16887
rect 8541 16841 8653 16887
rect 8699 16850 8712 16887
rect 8764 16887 9384 16902
rect 8764 16850 8811 16887
rect 8699 16841 8811 16850
rect 8857 16841 8969 16887
rect 9015 16841 9128 16887
rect 9174 16841 9286 16887
rect 9332 16850 9384 16887
rect 9436 16887 9832 16902
rect 9436 16850 9444 16887
rect 9332 16841 9444 16850
rect 9490 16841 9602 16887
rect 9648 16841 9760 16887
rect 9806 16850 9832 16887
rect 9884 16887 10504 16902
rect 10556 16887 10952 16902
rect 9884 16850 9918 16887
rect 9806 16841 9918 16850
rect 9964 16841 10076 16887
rect 10122 16841 10234 16887
rect 10280 16841 10392 16887
rect 10438 16850 10504 16887
rect 10438 16841 10551 16850
rect 10597 16841 10709 16887
rect 10755 16841 10867 16887
rect 10913 16850 10952 16887
rect 11004 16887 11624 16902
rect 11676 16887 12072 16902
rect 11004 16850 11025 16887
rect 10913 16841 11025 16850
rect 11071 16841 11183 16887
rect 11229 16841 11341 16887
rect 11387 16841 11499 16887
rect 11545 16850 11624 16887
rect 11545 16841 11658 16850
rect 11704 16841 11816 16887
rect 11862 16841 11974 16887
rect 12020 16850 12072 16887
rect 12124 16887 12744 16902
rect 12796 16887 13192 16902
rect 13244 16887 13864 16902
rect 13916 16887 14312 16902
rect 14364 16887 14984 16902
rect 15036 16887 15432 16902
rect 15484 16887 16104 16902
rect 16156 16887 16552 16902
rect 16604 16887 17224 16902
rect 17276 16887 17672 16902
rect 17724 16887 18344 16902
rect 12124 16850 12132 16887
rect 12020 16841 12132 16850
rect 12178 16841 12290 16887
rect 12336 16841 12448 16887
rect 12494 16841 12606 16887
rect 12652 16850 12744 16887
rect 12652 16841 12764 16850
rect 12810 16841 12922 16887
rect 12968 16841 13081 16887
rect 13127 16850 13192 16887
rect 13127 16841 13239 16850
rect 13285 16841 13397 16887
rect 13443 16841 13555 16887
rect 13601 16841 13713 16887
rect 13759 16850 13864 16887
rect 13759 16841 13871 16850
rect 13917 16841 14029 16887
rect 14075 16841 14187 16887
rect 14233 16850 14312 16887
rect 14233 16841 14345 16850
rect 14391 16841 14504 16887
rect 14550 16841 14662 16887
rect 14708 16841 14820 16887
rect 14866 16841 14978 16887
rect 15036 16850 15136 16887
rect 15024 16841 15136 16850
rect 15182 16841 15294 16887
rect 15340 16850 15432 16887
rect 15340 16841 15452 16850
rect 15498 16841 15610 16887
rect 15656 16841 15768 16887
rect 15814 16841 15927 16887
rect 15973 16841 16085 16887
rect 16156 16850 16243 16887
rect 16131 16841 16243 16850
rect 16289 16841 16401 16887
rect 16447 16850 16552 16887
rect 16447 16841 16559 16850
rect 16605 16841 16717 16887
rect 16763 16841 16875 16887
rect 16921 16841 17033 16887
rect 17079 16841 17192 16887
rect 17276 16850 17350 16887
rect 17238 16841 17350 16850
rect 17396 16841 17508 16887
rect 17554 16841 17666 16887
rect 17724 16850 17824 16887
rect 17712 16841 17824 16850
rect 17870 16841 17982 16887
rect 18028 16841 18140 16887
rect 18186 16841 18298 16887
rect 18396 16887 18792 16902
rect 18844 16887 19464 16902
rect 18396 16850 18456 16887
rect 18344 16841 18456 16850
rect 18502 16841 18615 16887
rect 18661 16841 18773 16887
rect 18844 16850 18931 16887
rect 18819 16841 18931 16850
rect 18977 16841 19089 16887
rect 19135 16841 19247 16887
rect 19293 16841 19405 16887
rect 19451 16850 19464 16887
rect 19516 16887 19912 16902
rect 19964 16887 20175 16902
rect 19516 16850 19563 16887
rect 19451 16841 19563 16850
rect 19609 16841 19721 16887
rect 19767 16841 19879 16887
rect 19964 16850 20038 16887
rect 19925 16841 20038 16850
rect 20084 16841 20175 16887
rect 1953 16778 20175 16841
rect 1953 16726 1992 16778
rect 2044 16726 2664 16778
rect 2716 16726 3112 16778
rect 3164 16726 3784 16778
rect 3836 16726 4232 16778
rect 4284 16726 4904 16778
rect 4956 16726 5352 16778
rect 5404 16726 6024 16778
rect 6076 16726 6472 16778
rect 6524 16726 7144 16778
rect 7196 16726 7592 16778
rect 7644 16726 8264 16778
rect 8316 16726 8712 16778
rect 8764 16726 9384 16778
rect 9436 16726 9832 16778
rect 9884 16726 10504 16778
rect 10556 16726 10952 16778
rect 11004 16726 11624 16778
rect 11676 16726 12072 16778
rect 12124 16726 12744 16778
rect 12796 16726 13192 16778
rect 13244 16726 13864 16778
rect 13916 16726 14312 16778
rect 14364 16726 14984 16778
rect 15036 16726 15432 16778
rect 15484 16726 16104 16778
rect 16156 16726 16552 16778
rect 16604 16726 17224 16778
rect 17276 16726 17672 16778
rect 17724 16726 18344 16778
rect 18396 16726 18792 16778
rect 18844 16726 19464 16778
rect 19516 16726 19912 16778
rect 19964 16726 20175 16778
rect 1953 16682 20175 16726
rect 1980 16654 2056 16682
rect 1980 16602 1992 16654
rect 2044 16602 2056 16654
rect 1980 16572 2056 16602
rect 2652 16654 2728 16682
rect 2652 16602 2664 16654
rect 2716 16602 2728 16654
rect 1980 16530 1995 16572
rect 2041 16530 2056 16572
rect 1980 16478 1992 16530
rect 2044 16478 2056 16530
rect 1980 16406 1995 16478
rect 2041 16406 2056 16478
rect 1980 16354 1992 16406
rect 2044 16354 2056 16406
rect 1980 16282 1995 16354
rect 2041 16282 2056 16354
rect 1980 16230 1992 16282
rect 2044 16230 2056 16282
rect 1980 16158 1995 16230
rect 2041 16158 2056 16230
rect 1980 16106 1992 16158
rect 2044 16106 2056 16158
rect 1980 16034 1995 16106
rect 2041 16034 2056 16106
rect 1980 15982 1992 16034
rect 2044 15982 2056 16034
rect 1980 15910 1995 15982
rect 2041 15910 2056 15982
rect 1980 15858 1992 15910
rect 2044 15858 2056 15910
rect 1980 15786 1995 15858
rect 2041 15786 2056 15858
rect 1980 15734 1992 15786
rect 2044 15734 2056 15786
rect 1980 15662 1995 15734
rect 2041 15662 2056 15734
rect 1980 15610 1992 15662
rect 2044 15610 2056 15662
rect 1980 15538 1995 15610
rect 2041 15538 2056 15610
rect 1980 15486 1992 15538
rect 2044 15486 2056 15538
rect 1980 15474 1995 15486
rect 2041 15474 2056 15486
rect 2219 16572 2265 16585
rect 1995 12585 2041 12598
rect 2443 16572 2489 16585
rect 2428 14996 2443 15008
rect 2652 16572 2728 16602
rect 3100 16654 3176 16682
rect 3100 16602 3112 16654
rect 3164 16602 3176 16654
rect 2652 16530 2667 16572
rect 2713 16530 2728 16572
rect 2652 16478 2664 16530
rect 2716 16478 2728 16530
rect 2652 16406 2667 16478
rect 2713 16406 2728 16478
rect 2652 16354 2664 16406
rect 2716 16354 2728 16406
rect 2652 16282 2667 16354
rect 2713 16282 2728 16354
rect 2652 16230 2664 16282
rect 2716 16230 2728 16282
rect 2652 16158 2667 16230
rect 2713 16158 2728 16230
rect 2652 16106 2664 16158
rect 2716 16106 2728 16158
rect 2652 16034 2667 16106
rect 2713 16034 2728 16106
rect 2652 15982 2664 16034
rect 2716 15982 2728 16034
rect 2652 15910 2667 15982
rect 2713 15910 2728 15982
rect 2652 15858 2664 15910
rect 2716 15858 2728 15910
rect 2652 15786 2667 15858
rect 2713 15786 2728 15858
rect 2652 15734 2664 15786
rect 2716 15734 2728 15786
rect 2652 15662 2667 15734
rect 2713 15662 2728 15734
rect 2652 15610 2664 15662
rect 2716 15610 2728 15662
rect 2652 15538 2667 15610
rect 2713 15538 2728 15610
rect 2652 15486 2664 15538
rect 2716 15486 2728 15538
rect 2652 15474 2667 15486
rect 2489 14996 2504 15008
rect 2428 14944 2440 14996
rect 2492 14944 2504 14996
rect 2428 14872 2443 14944
rect 2489 14872 2504 14944
rect 2428 14820 2440 14872
rect 2492 14820 2504 14872
rect 2428 14748 2443 14820
rect 2489 14748 2504 14820
rect 2428 14696 2440 14748
rect 2492 14696 2504 14748
rect 2428 14624 2443 14696
rect 2489 14624 2504 14696
rect 2428 14572 2440 14624
rect 2492 14572 2504 14624
rect 2428 14500 2443 14572
rect 2489 14500 2504 14572
rect 2428 14448 2440 14500
rect 2492 14448 2504 14500
rect 2428 14376 2443 14448
rect 2489 14376 2504 14448
rect 2428 14324 2440 14376
rect 2492 14324 2504 14376
rect 2428 14252 2443 14324
rect 2489 14252 2504 14324
rect 2428 14200 2440 14252
rect 2492 14200 2504 14252
rect 2428 14128 2443 14200
rect 2489 14128 2504 14200
rect 2428 14076 2440 14128
rect 2492 14076 2504 14128
rect 2428 14004 2443 14076
rect 2489 14004 2504 14076
rect 2428 13952 2440 14004
rect 2492 13952 2504 14004
rect 2428 13880 2443 13952
rect 2489 13880 2504 13952
rect 2428 13828 2440 13880
rect 2492 13828 2504 13880
rect 2428 13756 2443 13828
rect 2489 13756 2504 13828
rect 2428 13704 2440 13756
rect 2492 13704 2504 13756
rect 2428 13632 2443 13704
rect 2489 13632 2504 13704
rect 2428 13580 2440 13632
rect 2492 13580 2504 13632
rect 2428 13508 2443 13580
rect 2489 13508 2504 13580
rect 2428 13456 2440 13508
rect 2492 13456 2504 13508
rect 2428 13384 2443 13456
rect 2489 13384 2504 13456
rect 2428 13332 2440 13384
rect 2492 13332 2504 13384
rect 2428 13260 2443 13332
rect 2489 13260 2504 13332
rect 2428 13208 2440 13260
rect 2492 13208 2504 13260
rect 2428 13136 2443 13208
rect 2489 13136 2504 13208
rect 2428 13084 2440 13136
rect 2492 13084 2504 13136
rect 2428 13012 2443 13084
rect 2489 13012 2504 13084
rect 2428 12960 2440 13012
rect 2492 12960 2504 13012
rect 2428 12888 2443 12960
rect 2489 12888 2504 12960
rect 2428 12836 2440 12888
rect 2492 12836 2504 12888
rect 2428 12824 2443 12836
rect 2078 12427 2146 12438
rect 2078 12381 2089 12427
rect 2135 12381 2146 12427
rect 2078 11923 2146 12381
rect 1996 11911 2146 11923
rect 1996 11859 2008 11911
rect 2060 11905 2146 11911
rect 2060 11859 2089 11905
rect 2135 11859 2146 11905
rect 1996 11840 2146 11859
rect 2219 11958 2265 12598
rect 2489 12824 2504 12836
rect 2443 12585 2489 12598
rect 2713 15474 2728 15486
rect 2891 16572 2937 16585
rect 2876 14996 2891 15008
rect 3100 16572 3176 16602
rect 3772 16654 3848 16682
rect 3772 16602 3784 16654
rect 3836 16602 3848 16654
rect 3100 16530 3115 16572
rect 3161 16530 3176 16572
rect 3100 16478 3112 16530
rect 3164 16478 3176 16530
rect 3100 16406 3115 16478
rect 3161 16406 3176 16478
rect 3100 16354 3112 16406
rect 3164 16354 3176 16406
rect 3100 16282 3115 16354
rect 3161 16282 3176 16354
rect 3100 16230 3112 16282
rect 3164 16230 3176 16282
rect 3100 16158 3115 16230
rect 3161 16158 3176 16230
rect 3100 16106 3112 16158
rect 3164 16106 3176 16158
rect 3100 16034 3115 16106
rect 3161 16034 3176 16106
rect 3100 15982 3112 16034
rect 3164 15982 3176 16034
rect 3100 15910 3115 15982
rect 3161 15910 3176 15982
rect 3100 15858 3112 15910
rect 3164 15858 3176 15910
rect 3100 15786 3115 15858
rect 3161 15786 3176 15858
rect 3100 15734 3112 15786
rect 3164 15734 3176 15786
rect 3100 15662 3115 15734
rect 3161 15662 3176 15734
rect 3100 15610 3112 15662
rect 3164 15610 3176 15662
rect 3100 15538 3115 15610
rect 3161 15538 3176 15610
rect 3100 15486 3112 15538
rect 3164 15486 3176 15538
rect 3100 15474 3115 15486
rect 2937 14996 2952 15008
rect 2876 14944 2888 14996
rect 2940 14944 2952 14996
rect 2876 14872 2891 14944
rect 2937 14872 2952 14944
rect 2876 14820 2888 14872
rect 2940 14820 2952 14872
rect 2876 14748 2891 14820
rect 2937 14748 2952 14820
rect 2876 14696 2888 14748
rect 2940 14696 2952 14748
rect 2876 14624 2891 14696
rect 2937 14624 2952 14696
rect 2876 14572 2888 14624
rect 2940 14572 2952 14624
rect 2876 14500 2891 14572
rect 2937 14500 2952 14572
rect 2876 14448 2888 14500
rect 2940 14448 2952 14500
rect 2876 14376 2891 14448
rect 2937 14376 2952 14448
rect 2876 14324 2888 14376
rect 2940 14324 2952 14376
rect 2876 14252 2891 14324
rect 2937 14252 2952 14324
rect 2876 14200 2888 14252
rect 2940 14200 2952 14252
rect 2876 14128 2891 14200
rect 2937 14128 2952 14200
rect 2876 14076 2888 14128
rect 2940 14076 2952 14128
rect 2876 14004 2891 14076
rect 2937 14004 2952 14076
rect 2876 13952 2888 14004
rect 2940 13952 2952 14004
rect 2876 13880 2891 13952
rect 2937 13880 2952 13952
rect 2876 13828 2888 13880
rect 2940 13828 2952 13880
rect 2876 13756 2891 13828
rect 2937 13756 2952 13828
rect 2876 13704 2888 13756
rect 2940 13704 2952 13756
rect 2876 13632 2891 13704
rect 2937 13632 2952 13704
rect 2876 13580 2888 13632
rect 2940 13580 2952 13632
rect 2876 13508 2891 13580
rect 2937 13508 2952 13580
rect 2876 13456 2888 13508
rect 2940 13456 2952 13508
rect 2876 13384 2891 13456
rect 2937 13384 2952 13456
rect 2876 13332 2888 13384
rect 2940 13332 2952 13384
rect 2876 13260 2891 13332
rect 2937 13260 2952 13332
rect 2876 13208 2888 13260
rect 2940 13208 2952 13260
rect 2876 13136 2891 13208
rect 2937 13136 2952 13208
rect 2876 13084 2888 13136
rect 2940 13084 2952 13136
rect 2876 13012 2891 13084
rect 2937 13012 2952 13084
rect 2876 12960 2888 13012
rect 2940 12960 2952 13012
rect 2876 12888 2891 12960
rect 2937 12888 2952 12960
rect 2876 12836 2888 12888
rect 2940 12836 2952 12888
rect 2876 12824 2891 12836
rect 2667 12274 2713 12598
rect 2937 12824 2952 12836
rect 2891 12585 2937 12598
rect 3161 15474 3176 15486
rect 3339 16572 3385 16585
rect 3115 12585 3161 12598
rect 3563 16572 3609 16585
rect 3548 14996 3563 15008
rect 3772 16572 3848 16602
rect 4220 16654 4296 16682
rect 4220 16602 4232 16654
rect 4284 16602 4296 16654
rect 3772 16530 3787 16572
rect 3833 16530 3848 16572
rect 3772 16478 3784 16530
rect 3836 16478 3848 16530
rect 3772 16406 3787 16478
rect 3833 16406 3848 16478
rect 3772 16354 3784 16406
rect 3836 16354 3848 16406
rect 3772 16282 3787 16354
rect 3833 16282 3848 16354
rect 3772 16230 3784 16282
rect 3836 16230 3848 16282
rect 3772 16158 3787 16230
rect 3833 16158 3848 16230
rect 3772 16106 3784 16158
rect 3836 16106 3848 16158
rect 3772 16034 3787 16106
rect 3833 16034 3848 16106
rect 3772 15982 3784 16034
rect 3836 15982 3848 16034
rect 3772 15910 3787 15982
rect 3833 15910 3848 15982
rect 3772 15858 3784 15910
rect 3836 15858 3848 15910
rect 3772 15786 3787 15858
rect 3833 15786 3848 15858
rect 3772 15734 3784 15786
rect 3836 15734 3848 15786
rect 3772 15662 3787 15734
rect 3833 15662 3848 15734
rect 3772 15610 3784 15662
rect 3836 15610 3848 15662
rect 3772 15538 3787 15610
rect 3833 15538 3848 15610
rect 3772 15486 3784 15538
rect 3836 15486 3848 15538
rect 3772 15474 3787 15486
rect 3609 14996 3624 15008
rect 3548 14944 3560 14996
rect 3612 14944 3624 14996
rect 3548 14872 3563 14944
rect 3609 14872 3624 14944
rect 3548 14820 3560 14872
rect 3612 14820 3624 14872
rect 3548 14748 3563 14820
rect 3609 14748 3624 14820
rect 3548 14696 3560 14748
rect 3612 14696 3624 14748
rect 3548 14624 3563 14696
rect 3609 14624 3624 14696
rect 3548 14572 3560 14624
rect 3612 14572 3624 14624
rect 3548 14500 3563 14572
rect 3609 14500 3624 14572
rect 3548 14448 3560 14500
rect 3612 14448 3624 14500
rect 3548 14376 3563 14448
rect 3609 14376 3624 14448
rect 3548 14324 3560 14376
rect 3612 14324 3624 14376
rect 3548 14252 3563 14324
rect 3609 14252 3624 14324
rect 3548 14200 3560 14252
rect 3612 14200 3624 14252
rect 3548 14128 3563 14200
rect 3609 14128 3624 14200
rect 3548 14076 3560 14128
rect 3612 14076 3624 14128
rect 3548 14004 3563 14076
rect 3609 14004 3624 14076
rect 3548 13952 3560 14004
rect 3612 13952 3624 14004
rect 3548 13880 3563 13952
rect 3609 13880 3624 13952
rect 3548 13828 3560 13880
rect 3612 13828 3624 13880
rect 3548 13756 3563 13828
rect 3609 13756 3624 13828
rect 3548 13704 3560 13756
rect 3612 13704 3624 13756
rect 3548 13632 3563 13704
rect 3609 13632 3624 13704
rect 3548 13580 3560 13632
rect 3612 13580 3624 13632
rect 3548 13508 3563 13580
rect 3609 13508 3624 13580
rect 3548 13456 3560 13508
rect 3612 13456 3624 13508
rect 3548 13384 3563 13456
rect 3609 13384 3624 13456
rect 3548 13332 3560 13384
rect 3612 13332 3624 13384
rect 3548 13260 3563 13332
rect 3609 13260 3624 13332
rect 3548 13208 3560 13260
rect 3612 13208 3624 13260
rect 3548 13136 3563 13208
rect 3609 13136 3624 13208
rect 3548 13084 3560 13136
rect 3612 13084 3624 13136
rect 3548 13012 3563 13084
rect 3609 13012 3624 13084
rect 3548 12960 3560 13012
rect 3612 12960 3624 13012
rect 3548 12888 3563 12960
rect 3609 12888 3624 12960
rect 3548 12836 3560 12888
rect 3612 12836 3624 12888
rect 3548 12824 3563 12836
rect 2905 12458 3067 12469
rect 2905 12412 2916 12458
rect 3056 12412 3067 12458
rect 2905 12401 3067 12412
rect 3198 12427 3266 12438
rect 2575 12263 2831 12274
rect 2575 12217 2586 12263
rect 2820 12217 2831 12263
rect 2575 12206 2831 12217
rect 3002 11958 3048 12401
rect 3198 12381 3209 12427
rect 3255 12381 3266 12427
rect 2219 11947 3067 11958
rect 2219 11901 2916 11947
rect 3056 11901 3067 11947
rect 3198 11923 3266 12381
rect 2219 11890 3067 11901
rect 3116 11911 3266 11923
rect 1995 11757 2041 11770
rect 1248 11266 1843 11393
rect 1007 10945 1602 11101
rect 765 10571 1360 10724
rect 1231 1158 1360 10571
rect 1473 1158 1602 10945
rect 408 1117 532 1155
rect 408 1065 444 1117
rect 496 1065 532 1117
rect 408 899 532 1065
rect 408 847 444 899
rect 496 847 532 899
rect 408 807 532 847
rect 1231 1117 1361 1158
rect 1231 1065 1270 1117
rect 1322 1065 1361 1117
rect 1231 899 1361 1065
rect 1231 847 1270 899
rect 1322 847 1361 899
rect 1231 807 1361 847
rect 1472 1117 1602 1158
rect 1472 1065 1511 1117
rect 1563 1065 1602 1117
rect 1472 899 1602 1065
rect 1472 847 1511 899
rect 1563 847 1602 899
rect 1472 807 1602 847
rect 1231 806 1360 807
rect 1473 806 1602 807
rect 1714 1158 1843 11266
rect 1995 10940 2041 10997
rect 1995 10837 2041 10894
rect 1995 10734 2041 10791
rect 1995 10631 2041 10688
rect 1995 10528 2041 10585
rect 1995 10425 2041 10482
rect 1995 10322 2041 10379
rect 1995 10219 2041 10276
rect 1995 10116 2041 10173
rect 1961 10070 1995 10109
rect 2219 11757 2265 11890
rect 3116 11859 3128 11911
rect 3180 11905 3266 11911
rect 3180 11859 3209 11905
rect 3255 11859 3266 11905
rect 3116 11840 3266 11859
rect 3339 11958 3385 12598
rect 3609 12824 3624 12836
rect 3563 12585 3609 12598
rect 3833 15474 3848 15486
rect 4011 16572 4057 16585
rect 3996 14996 4011 15008
rect 4220 16572 4296 16602
rect 4892 16654 4968 16682
rect 4892 16602 4904 16654
rect 4956 16602 4968 16654
rect 4220 16530 4235 16572
rect 4281 16530 4296 16572
rect 4220 16478 4232 16530
rect 4284 16478 4296 16530
rect 4220 16406 4235 16478
rect 4281 16406 4296 16478
rect 4220 16354 4232 16406
rect 4284 16354 4296 16406
rect 4220 16282 4235 16354
rect 4281 16282 4296 16354
rect 4220 16230 4232 16282
rect 4284 16230 4296 16282
rect 4220 16158 4235 16230
rect 4281 16158 4296 16230
rect 4220 16106 4232 16158
rect 4284 16106 4296 16158
rect 4220 16034 4235 16106
rect 4281 16034 4296 16106
rect 4220 15982 4232 16034
rect 4284 15982 4296 16034
rect 4220 15910 4235 15982
rect 4281 15910 4296 15982
rect 4220 15858 4232 15910
rect 4284 15858 4296 15910
rect 4220 15786 4235 15858
rect 4281 15786 4296 15858
rect 4220 15734 4232 15786
rect 4284 15734 4296 15786
rect 4220 15662 4235 15734
rect 4281 15662 4296 15734
rect 4220 15610 4232 15662
rect 4284 15610 4296 15662
rect 4220 15538 4235 15610
rect 4281 15538 4296 15610
rect 4220 15486 4232 15538
rect 4284 15486 4296 15538
rect 4220 15474 4235 15486
rect 4057 14996 4072 15008
rect 3996 14944 4008 14996
rect 4060 14944 4072 14996
rect 3996 14872 4011 14944
rect 4057 14872 4072 14944
rect 3996 14820 4008 14872
rect 4060 14820 4072 14872
rect 3996 14748 4011 14820
rect 4057 14748 4072 14820
rect 3996 14696 4008 14748
rect 4060 14696 4072 14748
rect 3996 14624 4011 14696
rect 4057 14624 4072 14696
rect 3996 14572 4008 14624
rect 4060 14572 4072 14624
rect 3996 14500 4011 14572
rect 4057 14500 4072 14572
rect 3996 14448 4008 14500
rect 4060 14448 4072 14500
rect 3996 14376 4011 14448
rect 4057 14376 4072 14448
rect 3996 14324 4008 14376
rect 4060 14324 4072 14376
rect 3996 14252 4011 14324
rect 4057 14252 4072 14324
rect 3996 14200 4008 14252
rect 4060 14200 4072 14252
rect 3996 14128 4011 14200
rect 4057 14128 4072 14200
rect 3996 14076 4008 14128
rect 4060 14076 4072 14128
rect 3996 14004 4011 14076
rect 4057 14004 4072 14076
rect 3996 13952 4008 14004
rect 4060 13952 4072 14004
rect 3996 13880 4011 13952
rect 4057 13880 4072 13952
rect 3996 13828 4008 13880
rect 4060 13828 4072 13880
rect 3996 13756 4011 13828
rect 4057 13756 4072 13828
rect 3996 13704 4008 13756
rect 4060 13704 4072 13756
rect 3996 13632 4011 13704
rect 4057 13632 4072 13704
rect 3996 13580 4008 13632
rect 4060 13580 4072 13632
rect 3996 13508 4011 13580
rect 4057 13508 4072 13580
rect 3996 13456 4008 13508
rect 4060 13456 4072 13508
rect 3996 13384 4011 13456
rect 4057 13384 4072 13456
rect 3996 13332 4008 13384
rect 4060 13332 4072 13384
rect 3996 13260 4011 13332
rect 4057 13260 4072 13332
rect 3996 13208 4008 13260
rect 4060 13208 4072 13260
rect 3996 13136 4011 13208
rect 4057 13136 4072 13208
rect 3996 13084 4008 13136
rect 4060 13084 4072 13136
rect 3996 13012 4011 13084
rect 4057 13012 4072 13084
rect 3996 12960 4008 13012
rect 4060 12960 4072 13012
rect 3996 12888 4011 12960
rect 4057 12888 4072 12960
rect 3996 12836 4008 12888
rect 4060 12836 4072 12888
rect 3996 12824 4011 12836
rect 3787 12274 3833 12598
rect 4057 12824 4072 12836
rect 4011 12585 4057 12598
rect 4281 15474 4296 15486
rect 4459 16572 4505 16585
rect 4235 12585 4281 12598
rect 4683 16572 4729 16585
rect 4668 14996 4683 15008
rect 4892 16572 4968 16602
rect 5340 16654 5416 16682
rect 5340 16602 5352 16654
rect 5404 16602 5416 16654
rect 4892 16530 4907 16572
rect 4953 16530 4968 16572
rect 4892 16478 4904 16530
rect 4956 16478 4968 16530
rect 4892 16406 4907 16478
rect 4953 16406 4968 16478
rect 4892 16354 4904 16406
rect 4956 16354 4968 16406
rect 4892 16282 4907 16354
rect 4953 16282 4968 16354
rect 4892 16230 4904 16282
rect 4956 16230 4968 16282
rect 4892 16158 4907 16230
rect 4953 16158 4968 16230
rect 4892 16106 4904 16158
rect 4956 16106 4968 16158
rect 4892 16034 4907 16106
rect 4953 16034 4968 16106
rect 4892 15982 4904 16034
rect 4956 15982 4968 16034
rect 4892 15910 4907 15982
rect 4953 15910 4968 15982
rect 4892 15858 4904 15910
rect 4956 15858 4968 15910
rect 4892 15786 4907 15858
rect 4953 15786 4968 15858
rect 4892 15734 4904 15786
rect 4956 15734 4968 15786
rect 4892 15662 4907 15734
rect 4953 15662 4968 15734
rect 4892 15610 4904 15662
rect 4956 15610 4968 15662
rect 4892 15538 4907 15610
rect 4953 15538 4968 15610
rect 4892 15486 4904 15538
rect 4956 15486 4968 15538
rect 4892 15474 4907 15486
rect 4729 14996 4744 15008
rect 4668 14944 4680 14996
rect 4732 14944 4744 14996
rect 4668 14872 4683 14944
rect 4729 14872 4744 14944
rect 4668 14820 4680 14872
rect 4732 14820 4744 14872
rect 4668 14748 4683 14820
rect 4729 14748 4744 14820
rect 4668 14696 4680 14748
rect 4732 14696 4744 14748
rect 4668 14624 4683 14696
rect 4729 14624 4744 14696
rect 4668 14572 4680 14624
rect 4732 14572 4744 14624
rect 4668 14500 4683 14572
rect 4729 14500 4744 14572
rect 4668 14448 4680 14500
rect 4732 14448 4744 14500
rect 4668 14376 4683 14448
rect 4729 14376 4744 14448
rect 4668 14324 4680 14376
rect 4732 14324 4744 14376
rect 4668 14252 4683 14324
rect 4729 14252 4744 14324
rect 4668 14200 4680 14252
rect 4732 14200 4744 14252
rect 4668 14128 4683 14200
rect 4729 14128 4744 14200
rect 4668 14076 4680 14128
rect 4732 14076 4744 14128
rect 4668 14004 4683 14076
rect 4729 14004 4744 14076
rect 4668 13952 4680 14004
rect 4732 13952 4744 14004
rect 4668 13880 4683 13952
rect 4729 13880 4744 13952
rect 4668 13828 4680 13880
rect 4732 13828 4744 13880
rect 4668 13756 4683 13828
rect 4729 13756 4744 13828
rect 4668 13704 4680 13756
rect 4732 13704 4744 13756
rect 4668 13632 4683 13704
rect 4729 13632 4744 13704
rect 4668 13580 4680 13632
rect 4732 13580 4744 13632
rect 4668 13508 4683 13580
rect 4729 13508 4744 13580
rect 4668 13456 4680 13508
rect 4732 13456 4744 13508
rect 4668 13384 4683 13456
rect 4729 13384 4744 13456
rect 4668 13332 4680 13384
rect 4732 13332 4744 13384
rect 4668 13260 4683 13332
rect 4729 13260 4744 13332
rect 4668 13208 4680 13260
rect 4732 13208 4744 13260
rect 4668 13136 4683 13208
rect 4729 13136 4744 13208
rect 4668 13084 4680 13136
rect 4732 13084 4744 13136
rect 4668 13012 4683 13084
rect 4729 13012 4744 13084
rect 4668 12960 4680 13012
rect 4732 12960 4744 13012
rect 4668 12888 4683 12960
rect 4729 12888 4744 12960
rect 4668 12836 4680 12888
rect 4732 12836 4744 12888
rect 4668 12824 4683 12836
rect 4025 12458 4187 12469
rect 4025 12412 4036 12458
rect 4176 12412 4187 12458
rect 4025 12401 4187 12412
rect 4318 12427 4386 12438
rect 3695 12263 3951 12274
rect 3695 12217 3706 12263
rect 3940 12217 3951 12263
rect 3695 12206 3951 12217
rect 4122 11958 4168 12401
rect 4318 12381 4329 12427
rect 4375 12381 4386 12427
rect 3339 11947 4187 11958
rect 3339 11901 4036 11947
rect 4176 11901 4187 11947
rect 4318 11923 4386 12381
rect 3339 11890 4187 11901
rect 4236 11911 4386 11923
rect 2428 11758 2504 11770
rect 2428 11706 2440 11758
rect 2492 11706 2504 11758
rect 2428 11634 2443 11706
rect 2489 11634 2504 11706
rect 2428 11582 2440 11634
rect 2492 11582 2504 11634
rect 2428 11510 2443 11582
rect 2489 11510 2504 11582
rect 2428 11458 2440 11510
rect 2492 11458 2504 11510
rect 2428 11446 2443 11458
rect 2219 10940 2265 10997
rect 2219 10837 2265 10894
rect 2219 10734 2265 10791
rect 2219 10631 2265 10688
rect 2219 10528 2265 10585
rect 2219 10425 2265 10482
rect 2219 10322 2265 10379
rect 2219 10219 2265 10276
rect 2219 10116 2265 10173
rect 2041 10070 2076 10109
rect 1961 10013 2076 10070
rect 1961 9967 1995 10013
rect 2041 9967 2076 10013
rect 1961 9863 2076 9967
rect 2219 10013 2265 10070
rect 2219 9954 2265 9967
rect 2489 11446 2504 11458
rect 2667 11757 2713 11770
rect 2443 10940 2489 10997
rect 2443 10837 2489 10894
rect 2443 10734 2489 10791
rect 2443 10631 2489 10688
rect 2443 10528 2489 10585
rect 2443 10425 2489 10482
rect 2443 10322 2489 10379
rect 2443 10219 2489 10276
rect 2443 10116 2489 10173
rect 2876 11758 2952 11770
rect 2876 11706 2888 11758
rect 2940 11706 2952 11758
rect 2876 11634 2891 11706
rect 2937 11634 2952 11706
rect 2876 11582 2888 11634
rect 2940 11582 2952 11634
rect 2876 11510 2891 11582
rect 2937 11510 2952 11582
rect 2876 11458 2888 11510
rect 2940 11458 2952 11510
rect 2876 11446 2891 11458
rect 2667 10940 2713 10997
rect 2667 10837 2713 10894
rect 2667 10734 2713 10791
rect 2667 10631 2713 10688
rect 2667 10528 2713 10585
rect 2667 10425 2713 10482
rect 2667 10322 2713 10379
rect 2667 10219 2713 10276
rect 2667 10116 2713 10173
rect 2443 10013 2489 10070
rect 2443 9954 2489 9967
rect 2633 10070 2667 10109
rect 2937 11446 2952 11458
rect 3115 11757 3161 11770
rect 2891 10940 2937 10997
rect 2891 10837 2937 10894
rect 2891 10734 2937 10791
rect 2891 10631 2937 10688
rect 2891 10528 2937 10585
rect 2891 10425 2937 10482
rect 2891 10322 2937 10379
rect 2891 10219 2937 10276
rect 2891 10116 2937 10173
rect 2713 10070 2748 10109
rect 2633 10013 2748 10070
rect 2633 9967 2667 10013
rect 2713 9967 2748 10013
rect 2633 9863 2748 9967
rect 3115 10940 3161 10997
rect 3115 10837 3161 10894
rect 3115 10734 3161 10791
rect 3115 10631 3161 10688
rect 3115 10528 3161 10585
rect 3115 10425 3161 10482
rect 3115 10322 3161 10379
rect 3115 10219 3161 10276
rect 3115 10116 3161 10173
rect 2891 10013 2937 10070
rect 2891 9954 2937 9967
rect 3081 10070 3115 10109
rect 3339 11757 3385 11890
rect 4236 11859 4248 11911
rect 4300 11905 4386 11911
rect 4300 11859 4329 11905
rect 4375 11859 4386 11905
rect 4236 11840 4386 11859
rect 4459 11958 4505 12598
rect 4729 12824 4744 12836
rect 4683 12585 4729 12598
rect 4953 15474 4968 15486
rect 5131 16572 5177 16585
rect 5116 14996 5131 15008
rect 5340 16572 5416 16602
rect 6012 16654 6088 16682
rect 6012 16602 6024 16654
rect 6076 16602 6088 16654
rect 5340 16530 5355 16572
rect 5401 16530 5416 16572
rect 5340 16478 5352 16530
rect 5404 16478 5416 16530
rect 5340 16406 5355 16478
rect 5401 16406 5416 16478
rect 5340 16354 5352 16406
rect 5404 16354 5416 16406
rect 5340 16282 5355 16354
rect 5401 16282 5416 16354
rect 5340 16230 5352 16282
rect 5404 16230 5416 16282
rect 5340 16158 5355 16230
rect 5401 16158 5416 16230
rect 5340 16106 5352 16158
rect 5404 16106 5416 16158
rect 5340 16034 5355 16106
rect 5401 16034 5416 16106
rect 5340 15982 5352 16034
rect 5404 15982 5416 16034
rect 5340 15910 5355 15982
rect 5401 15910 5416 15982
rect 5340 15858 5352 15910
rect 5404 15858 5416 15910
rect 5340 15786 5355 15858
rect 5401 15786 5416 15858
rect 5340 15734 5352 15786
rect 5404 15734 5416 15786
rect 5340 15662 5355 15734
rect 5401 15662 5416 15734
rect 5340 15610 5352 15662
rect 5404 15610 5416 15662
rect 5340 15538 5355 15610
rect 5401 15538 5416 15610
rect 5340 15486 5352 15538
rect 5404 15486 5416 15538
rect 5340 15474 5355 15486
rect 5177 14996 5192 15008
rect 5116 14944 5128 14996
rect 5180 14944 5192 14996
rect 5116 14872 5131 14944
rect 5177 14872 5192 14944
rect 5116 14820 5128 14872
rect 5180 14820 5192 14872
rect 5116 14748 5131 14820
rect 5177 14748 5192 14820
rect 5116 14696 5128 14748
rect 5180 14696 5192 14748
rect 5116 14624 5131 14696
rect 5177 14624 5192 14696
rect 5116 14572 5128 14624
rect 5180 14572 5192 14624
rect 5116 14500 5131 14572
rect 5177 14500 5192 14572
rect 5116 14448 5128 14500
rect 5180 14448 5192 14500
rect 5116 14376 5131 14448
rect 5177 14376 5192 14448
rect 5116 14324 5128 14376
rect 5180 14324 5192 14376
rect 5116 14252 5131 14324
rect 5177 14252 5192 14324
rect 5116 14200 5128 14252
rect 5180 14200 5192 14252
rect 5116 14128 5131 14200
rect 5177 14128 5192 14200
rect 5116 14076 5128 14128
rect 5180 14076 5192 14128
rect 5116 14004 5131 14076
rect 5177 14004 5192 14076
rect 5116 13952 5128 14004
rect 5180 13952 5192 14004
rect 5116 13880 5131 13952
rect 5177 13880 5192 13952
rect 5116 13828 5128 13880
rect 5180 13828 5192 13880
rect 5116 13756 5131 13828
rect 5177 13756 5192 13828
rect 5116 13704 5128 13756
rect 5180 13704 5192 13756
rect 5116 13632 5131 13704
rect 5177 13632 5192 13704
rect 5116 13580 5128 13632
rect 5180 13580 5192 13632
rect 5116 13508 5131 13580
rect 5177 13508 5192 13580
rect 5116 13456 5128 13508
rect 5180 13456 5192 13508
rect 5116 13384 5131 13456
rect 5177 13384 5192 13456
rect 5116 13332 5128 13384
rect 5180 13332 5192 13384
rect 5116 13260 5131 13332
rect 5177 13260 5192 13332
rect 5116 13208 5128 13260
rect 5180 13208 5192 13260
rect 5116 13136 5131 13208
rect 5177 13136 5192 13208
rect 5116 13084 5128 13136
rect 5180 13084 5192 13136
rect 5116 13012 5131 13084
rect 5177 13012 5192 13084
rect 5116 12960 5128 13012
rect 5180 12960 5192 13012
rect 5116 12888 5131 12960
rect 5177 12888 5192 12960
rect 5116 12836 5128 12888
rect 5180 12836 5192 12888
rect 5116 12824 5131 12836
rect 4907 12274 4953 12598
rect 5177 12824 5192 12836
rect 5131 12585 5177 12598
rect 5401 15474 5416 15486
rect 5579 16572 5625 16585
rect 5355 12585 5401 12598
rect 5803 16572 5849 16585
rect 5788 14996 5803 15008
rect 6012 16572 6088 16602
rect 6460 16654 6536 16682
rect 6460 16602 6472 16654
rect 6524 16602 6536 16654
rect 6012 16530 6027 16572
rect 6073 16530 6088 16572
rect 6012 16478 6024 16530
rect 6076 16478 6088 16530
rect 6012 16406 6027 16478
rect 6073 16406 6088 16478
rect 6012 16354 6024 16406
rect 6076 16354 6088 16406
rect 6012 16282 6027 16354
rect 6073 16282 6088 16354
rect 6012 16230 6024 16282
rect 6076 16230 6088 16282
rect 6012 16158 6027 16230
rect 6073 16158 6088 16230
rect 6012 16106 6024 16158
rect 6076 16106 6088 16158
rect 6012 16034 6027 16106
rect 6073 16034 6088 16106
rect 6012 15982 6024 16034
rect 6076 15982 6088 16034
rect 6012 15910 6027 15982
rect 6073 15910 6088 15982
rect 6012 15858 6024 15910
rect 6076 15858 6088 15910
rect 6012 15786 6027 15858
rect 6073 15786 6088 15858
rect 6012 15734 6024 15786
rect 6076 15734 6088 15786
rect 6012 15662 6027 15734
rect 6073 15662 6088 15734
rect 6012 15610 6024 15662
rect 6076 15610 6088 15662
rect 6012 15538 6027 15610
rect 6073 15538 6088 15610
rect 6012 15486 6024 15538
rect 6076 15486 6088 15538
rect 6012 15474 6027 15486
rect 5849 14996 5864 15008
rect 5788 14944 5800 14996
rect 5852 14944 5864 14996
rect 5788 14872 5803 14944
rect 5849 14872 5864 14944
rect 5788 14820 5800 14872
rect 5852 14820 5864 14872
rect 5788 14748 5803 14820
rect 5849 14748 5864 14820
rect 5788 14696 5800 14748
rect 5852 14696 5864 14748
rect 5788 14624 5803 14696
rect 5849 14624 5864 14696
rect 5788 14572 5800 14624
rect 5852 14572 5864 14624
rect 5788 14500 5803 14572
rect 5849 14500 5864 14572
rect 5788 14448 5800 14500
rect 5852 14448 5864 14500
rect 5788 14376 5803 14448
rect 5849 14376 5864 14448
rect 5788 14324 5800 14376
rect 5852 14324 5864 14376
rect 5788 14252 5803 14324
rect 5849 14252 5864 14324
rect 5788 14200 5800 14252
rect 5852 14200 5864 14252
rect 5788 14128 5803 14200
rect 5849 14128 5864 14200
rect 5788 14076 5800 14128
rect 5852 14076 5864 14128
rect 5788 14004 5803 14076
rect 5849 14004 5864 14076
rect 5788 13952 5800 14004
rect 5852 13952 5864 14004
rect 5788 13880 5803 13952
rect 5849 13880 5864 13952
rect 5788 13828 5800 13880
rect 5852 13828 5864 13880
rect 5788 13756 5803 13828
rect 5849 13756 5864 13828
rect 5788 13704 5800 13756
rect 5852 13704 5864 13756
rect 5788 13632 5803 13704
rect 5849 13632 5864 13704
rect 5788 13580 5800 13632
rect 5852 13580 5864 13632
rect 5788 13508 5803 13580
rect 5849 13508 5864 13580
rect 5788 13456 5800 13508
rect 5852 13456 5864 13508
rect 5788 13384 5803 13456
rect 5849 13384 5864 13456
rect 5788 13332 5800 13384
rect 5852 13332 5864 13384
rect 5788 13260 5803 13332
rect 5849 13260 5864 13332
rect 5788 13208 5800 13260
rect 5852 13208 5864 13260
rect 5788 13136 5803 13208
rect 5849 13136 5864 13208
rect 5788 13084 5800 13136
rect 5852 13084 5864 13136
rect 5788 13012 5803 13084
rect 5849 13012 5864 13084
rect 5788 12960 5800 13012
rect 5852 12960 5864 13012
rect 5788 12888 5803 12960
rect 5849 12888 5864 12960
rect 5788 12836 5800 12888
rect 5852 12836 5864 12888
rect 5788 12824 5803 12836
rect 5145 12458 5307 12469
rect 5145 12412 5156 12458
rect 5296 12412 5307 12458
rect 5145 12401 5307 12412
rect 5438 12427 5506 12438
rect 4815 12263 5071 12274
rect 4815 12217 4826 12263
rect 5060 12217 5071 12263
rect 4815 12206 5071 12217
rect 5242 11958 5288 12401
rect 5438 12381 5449 12427
rect 5495 12381 5506 12427
rect 4459 11947 5307 11958
rect 4459 11901 5156 11947
rect 5296 11901 5307 11947
rect 5438 11923 5506 12381
rect 4459 11890 5307 11901
rect 5356 11911 5506 11923
rect 3548 11758 3624 11770
rect 3548 11706 3560 11758
rect 3612 11706 3624 11758
rect 3548 11634 3563 11706
rect 3609 11634 3624 11706
rect 3548 11582 3560 11634
rect 3612 11582 3624 11634
rect 3548 11510 3563 11582
rect 3609 11510 3624 11582
rect 3548 11458 3560 11510
rect 3612 11458 3624 11510
rect 3548 11446 3563 11458
rect 3339 10940 3385 10997
rect 3339 10837 3385 10894
rect 3339 10734 3385 10791
rect 3339 10631 3385 10688
rect 3339 10528 3385 10585
rect 3339 10425 3385 10482
rect 3339 10322 3385 10379
rect 3339 10219 3385 10276
rect 3339 10116 3385 10173
rect 3161 10070 3196 10109
rect 3081 10013 3196 10070
rect 3081 9967 3115 10013
rect 3161 9967 3196 10013
rect 3081 9863 3196 9967
rect 3339 10013 3385 10070
rect 3339 9954 3385 9967
rect 3609 11446 3624 11458
rect 3787 11757 3833 11770
rect 3563 10940 3609 10997
rect 3563 10837 3609 10894
rect 3563 10734 3609 10791
rect 3563 10631 3609 10688
rect 3563 10528 3609 10585
rect 3563 10425 3609 10482
rect 3563 10322 3609 10379
rect 3563 10219 3609 10276
rect 3563 10116 3609 10173
rect 3996 11758 4072 11770
rect 3996 11706 4008 11758
rect 4060 11706 4072 11758
rect 3996 11634 4011 11706
rect 4057 11634 4072 11706
rect 3996 11582 4008 11634
rect 4060 11582 4072 11634
rect 3996 11510 4011 11582
rect 4057 11510 4072 11582
rect 3996 11458 4008 11510
rect 4060 11458 4072 11510
rect 3996 11446 4011 11458
rect 3787 10940 3833 10997
rect 3787 10837 3833 10894
rect 3787 10734 3833 10791
rect 3787 10631 3833 10688
rect 3787 10528 3833 10585
rect 3787 10425 3833 10482
rect 3787 10322 3833 10379
rect 3787 10219 3833 10276
rect 3787 10116 3833 10173
rect 3563 10013 3609 10070
rect 3563 9954 3609 9967
rect 3753 10070 3787 10109
rect 4057 11446 4072 11458
rect 4235 11757 4281 11770
rect 4011 10940 4057 10997
rect 4011 10837 4057 10894
rect 4011 10734 4057 10791
rect 4011 10631 4057 10688
rect 4011 10528 4057 10585
rect 4011 10425 4057 10482
rect 4011 10322 4057 10379
rect 4011 10219 4057 10276
rect 4011 10116 4057 10173
rect 3833 10070 3868 10109
rect 3753 10013 3868 10070
rect 3753 9967 3787 10013
rect 3833 9967 3868 10013
rect 3753 9863 3868 9967
rect 4235 10940 4281 10997
rect 4235 10837 4281 10894
rect 4235 10734 4281 10791
rect 4235 10631 4281 10688
rect 4235 10528 4281 10585
rect 4235 10425 4281 10482
rect 4235 10322 4281 10379
rect 4235 10219 4281 10276
rect 4235 10116 4281 10173
rect 4011 10013 4057 10070
rect 4011 9954 4057 9967
rect 4201 10070 4235 10109
rect 4459 11757 4505 11890
rect 5356 11859 5368 11911
rect 5420 11905 5506 11911
rect 5420 11859 5449 11905
rect 5495 11859 5506 11905
rect 5356 11840 5506 11859
rect 5579 11958 5625 12598
rect 5849 12824 5864 12836
rect 5803 12585 5849 12598
rect 6073 15474 6088 15486
rect 6251 16572 6297 16585
rect 6236 14996 6251 15008
rect 6460 16572 6536 16602
rect 7132 16654 7208 16682
rect 7132 16602 7144 16654
rect 7196 16602 7208 16654
rect 6460 16530 6475 16572
rect 6521 16530 6536 16572
rect 6460 16478 6472 16530
rect 6524 16478 6536 16530
rect 6460 16406 6475 16478
rect 6521 16406 6536 16478
rect 6460 16354 6472 16406
rect 6524 16354 6536 16406
rect 6460 16282 6475 16354
rect 6521 16282 6536 16354
rect 6460 16230 6472 16282
rect 6524 16230 6536 16282
rect 6460 16158 6475 16230
rect 6521 16158 6536 16230
rect 6460 16106 6472 16158
rect 6524 16106 6536 16158
rect 6460 16034 6475 16106
rect 6521 16034 6536 16106
rect 6460 15982 6472 16034
rect 6524 15982 6536 16034
rect 6460 15910 6475 15982
rect 6521 15910 6536 15982
rect 6460 15858 6472 15910
rect 6524 15858 6536 15910
rect 6460 15786 6475 15858
rect 6521 15786 6536 15858
rect 6460 15734 6472 15786
rect 6524 15734 6536 15786
rect 6460 15662 6475 15734
rect 6521 15662 6536 15734
rect 6460 15610 6472 15662
rect 6524 15610 6536 15662
rect 6460 15538 6475 15610
rect 6521 15538 6536 15610
rect 6460 15486 6472 15538
rect 6524 15486 6536 15538
rect 6460 15474 6475 15486
rect 6297 14996 6312 15008
rect 6236 14944 6248 14996
rect 6300 14944 6312 14996
rect 6236 14872 6251 14944
rect 6297 14872 6312 14944
rect 6236 14820 6248 14872
rect 6300 14820 6312 14872
rect 6236 14748 6251 14820
rect 6297 14748 6312 14820
rect 6236 14696 6248 14748
rect 6300 14696 6312 14748
rect 6236 14624 6251 14696
rect 6297 14624 6312 14696
rect 6236 14572 6248 14624
rect 6300 14572 6312 14624
rect 6236 14500 6251 14572
rect 6297 14500 6312 14572
rect 6236 14448 6248 14500
rect 6300 14448 6312 14500
rect 6236 14376 6251 14448
rect 6297 14376 6312 14448
rect 6236 14324 6248 14376
rect 6300 14324 6312 14376
rect 6236 14252 6251 14324
rect 6297 14252 6312 14324
rect 6236 14200 6248 14252
rect 6300 14200 6312 14252
rect 6236 14128 6251 14200
rect 6297 14128 6312 14200
rect 6236 14076 6248 14128
rect 6300 14076 6312 14128
rect 6236 14004 6251 14076
rect 6297 14004 6312 14076
rect 6236 13952 6248 14004
rect 6300 13952 6312 14004
rect 6236 13880 6251 13952
rect 6297 13880 6312 13952
rect 6236 13828 6248 13880
rect 6300 13828 6312 13880
rect 6236 13756 6251 13828
rect 6297 13756 6312 13828
rect 6236 13704 6248 13756
rect 6300 13704 6312 13756
rect 6236 13632 6251 13704
rect 6297 13632 6312 13704
rect 6236 13580 6248 13632
rect 6300 13580 6312 13632
rect 6236 13508 6251 13580
rect 6297 13508 6312 13580
rect 6236 13456 6248 13508
rect 6300 13456 6312 13508
rect 6236 13384 6251 13456
rect 6297 13384 6312 13456
rect 6236 13332 6248 13384
rect 6300 13332 6312 13384
rect 6236 13260 6251 13332
rect 6297 13260 6312 13332
rect 6236 13208 6248 13260
rect 6300 13208 6312 13260
rect 6236 13136 6251 13208
rect 6297 13136 6312 13208
rect 6236 13084 6248 13136
rect 6300 13084 6312 13136
rect 6236 13012 6251 13084
rect 6297 13012 6312 13084
rect 6236 12960 6248 13012
rect 6300 12960 6312 13012
rect 6236 12888 6251 12960
rect 6297 12888 6312 12960
rect 6236 12836 6248 12888
rect 6300 12836 6312 12888
rect 6236 12824 6251 12836
rect 6027 12274 6073 12598
rect 6297 12824 6312 12836
rect 6251 12585 6297 12598
rect 6521 15474 6536 15486
rect 6699 16572 6745 16585
rect 6475 12585 6521 12598
rect 6923 16572 6969 16585
rect 6908 14996 6923 15008
rect 7132 16572 7208 16602
rect 7580 16654 7656 16682
rect 7580 16602 7592 16654
rect 7644 16602 7656 16654
rect 7132 16530 7147 16572
rect 7193 16530 7208 16572
rect 7132 16478 7144 16530
rect 7196 16478 7208 16530
rect 7132 16406 7147 16478
rect 7193 16406 7208 16478
rect 7132 16354 7144 16406
rect 7196 16354 7208 16406
rect 7132 16282 7147 16354
rect 7193 16282 7208 16354
rect 7132 16230 7144 16282
rect 7196 16230 7208 16282
rect 7132 16158 7147 16230
rect 7193 16158 7208 16230
rect 7132 16106 7144 16158
rect 7196 16106 7208 16158
rect 7132 16034 7147 16106
rect 7193 16034 7208 16106
rect 7132 15982 7144 16034
rect 7196 15982 7208 16034
rect 7132 15910 7147 15982
rect 7193 15910 7208 15982
rect 7132 15858 7144 15910
rect 7196 15858 7208 15910
rect 7132 15786 7147 15858
rect 7193 15786 7208 15858
rect 7132 15734 7144 15786
rect 7196 15734 7208 15786
rect 7132 15662 7147 15734
rect 7193 15662 7208 15734
rect 7132 15610 7144 15662
rect 7196 15610 7208 15662
rect 7132 15538 7147 15610
rect 7193 15538 7208 15610
rect 7132 15486 7144 15538
rect 7196 15486 7208 15538
rect 7132 15474 7147 15486
rect 6969 14996 6984 15008
rect 6908 14944 6920 14996
rect 6972 14944 6984 14996
rect 6908 14872 6923 14944
rect 6969 14872 6984 14944
rect 6908 14820 6920 14872
rect 6972 14820 6984 14872
rect 6908 14748 6923 14820
rect 6969 14748 6984 14820
rect 6908 14696 6920 14748
rect 6972 14696 6984 14748
rect 6908 14624 6923 14696
rect 6969 14624 6984 14696
rect 6908 14572 6920 14624
rect 6972 14572 6984 14624
rect 6908 14500 6923 14572
rect 6969 14500 6984 14572
rect 6908 14448 6920 14500
rect 6972 14448 6984 14500
rect 6908 14376 6923 14448
rect 6969 14376 6984 14448
rect 6908 14324 6920 14376
rect 6972 14324 6984 14376
rect 6908 14252 6923 14324
rect 6969 14252 6984 14324
rect 6908 14200 6920 14252
rect 6972 14200 6984 14252
rect 6908 14128 6923 14200
rect 6969 14128 6984 14200
rect 6908 14076 6920 14128
rect 6972 14076 6984 14128
rect 6908 14004 6923 14076
rect 6969 14004 6984 14076
rect 6908 13952 6920 14004
rect 6972 13952 6984 14004
rect 6908 13880 6923 13952
rect 6969 13880 6984 13952
rect 6908 13828 6920 13880
rect 6972 13828 6984 13880
rect 6908 13756 6923 13828
rect 6969 13756 6984 13828
rect 6908 13704 6920 13756
rect 6972 13704 6984 13756
rect 6908 13632 6923 13704
rect 6969 13632 6984 13704
rect 6908 13580 6920 13632
rect 6972 13580 6984 13632
rect 6908 13508 6923 13580
rect 6969 13508 6984 13580
rect 6908 13456 6920 13508
rect 6972 13456 6984 13508
rect 6908 13384 6923 13456
rect 6969 13384 6984 13456
rect 6908 13332 6920 13384
rect 6972 13332 6984 13384
rect 6908 13260 6923 13332
rect 6969 13260 6984 13332
rect 6908 13208 6920 13260
rect 6972 13208 6984 13260
rect 6908 13136 6923 13208
rect 6969 13136 6984 13208
rect 6908 13084 6920 13136
rect 6972 13084 6984 13136
rect 6908 13012 6923 13084
rect 6969 13012 6984 13084
rect 6908 12960 6920 13012
rect 6972 12960 6984 13012
rect 6908 12888 6923 12960
rect 6969 12888 6984 12960
rect 6908 12836 6920 12888
rect 6972 12836 6984 12888
rect 6908 12824 6923 12836
rect 6265 12458 6427 12469
rect 6265 12412 6276 12458
rect 6416 12412 6427 12458
rect 6265 12401 6427 12412
rect 6558 12427 6626 12438
rect 5935 12263 6191 12274
rect 5935 12217 5946 12263
rect 6180 12217 6191 12263
rect 5935 12206 6191 12217
rect 6362 11958 6408 12401
rect 6558 12381 6569 12427
rect 6615 12381 6626 12427
rect 5579 11947 6427 11958
rect 5579 11901 6276 11947
rect 6416 11901 6427 11947
rect 6558 11923 6626 12381
rect 5579 11890 6427 11901
rect 6476 11911 6626 11923
rect 4668 11758 4744 11770
rect 4668 11706 4680 11758
rect 4732 11706 4744 11758
rect 4668 11634 4683 11706
rect 4729 11634 4744 11706
rect 4668 11582 4680 11634
rect 4732 11582 4744 11634
rect 4668 11510 4683 11582
rect 4729 11510 4744 11582
rect 4668 11458 4680 11510
rect 4732 11458 4744 11510
rect 4668 11446 4683 11458
rect 4459 10940 4505 10997
rect 4459 10837 4505 10894
rect 4459 10734 4505 10791
rect 4459 10631 4505 10688
rect 4459 10528 4505 10585
rect 4459 10425 4505 10482
rect 4459 10322 4505 10379
rect 4459 10219 4505 10276
rect 4459 10116 4505 10173
rect 4281 10070 4316 10109
rect 4201 10013 4316 10070
rect 4201 9967 4235 10013
rect 4281 9967 4316 10013
rect 4201 9863 4316 9967
rect 4459 10013 4505 10070
rect 4459 9954 4505 9967
rect 4729 11446 4744 11458
rect 4907 11757 4953 11770
rect 4683 10940 4729 10997
rect 4683 10837 4729 10894
rect 4683 10734 4729 10791
rect 4683 10631 4729 10688
rect 4683 10528 4729 10585
rect 4683 10425 4729 10482
rect 4683 10322 4729 10379
rect 4683 10219 4729 10276
rect 4683 10116 4729 10173
rect 5116 11758 5192 11770
rect 5116 11706 5128 11758
rect 5180 11706 5192 11758
rect 5116 11634 5131 11706
rect 5177 11634 5192 11706
rect 5116 11582 5128 11634
rect 5180 11582 5192 11634
rect 5116 11510 5131 11582
rect 5177 11510 5192 11582
rect 5116 11458 5128 11510
rect 5180 11458 5192 11510
rect 5116 11446 5131 11458
rect 4907 10940 4953 10997
rect 4907 10837 4953 10894
rect 4907 10734 4953 10791
rect 4907 10631 4953 10688
rect 4907 10528 4953 10585
rect 4907 10425 4953 10482
rect 4907 10322 4953 10379
rect 4907 10219 4953 10276
rect 4907 10116 4953 10173
rect 4683 10013 4729 10070
rect 4683 9954 4729 9967
rect 4873 10070 4907 10109
rect 5177 11446 5192 11458
rect 5355 11757 5401 11770
rect 5131 10940 5177 10997
rect 5131 10837 5177 10894
rect 5131 10734 5177 10791
rect 5131 10631 5177 10688
rect 5131 10528 5177 10585
rect 5131 10425 5177 10482
rect 5131 10322 5177 10379
rect 5131 10219 5177 10276
rect 5131 10116 5177 10173
rect 4953 10070 4988 10109
rect 4873 10013 4988 10070
rect 4873 9967 4907 10013
rect 4953 9967 4988 10013
rect 4873 9863 4988 9967
rect 5355 10940 5401 10997
rect 5355 10837 5401 10894
rect 5355 10734 5401 10791
rect 5355 10631 5401 10688
rect 5355 10528 5401 10585
rect 5355 10425 5401 10482
rect 5355 10322 5401 10379
rect 5355 10219 5401 10276
rect 5355 10116 5401 10173
rect 5131 10013 5177 10070
rect 5131 9954 5177 9967
rect 5321 10070 5355 10109
rect 5579 11757 5625 11890
rect 6476 11859 6488 11911
rect 6540 11905 6626 11911
rect 6540 11859 6569 11905
rect 6615 11859 6626 11905
rect 6476 11840 6626 11859
rect 6699 11958 6745 12598
rect 6969 12824 6984 12836
rect 6923 12585 6969 12598
rect 7193 15474 7208 15486
rect 7371 16572 7417 16585
rect 7356 14996 7371 15008
rect 7580 16572 7656 16602
rect 8252 16654 8328 16682
rect 8252 16602 8264 16654
rect 8316 16602 8328 16654
rect 7580 16530 7595 16572
rect 7641 16530 7656 16572
rect 7580 16478 7592 16530
rect 7644 16478 7656 16530
rect 7580 16406 7595 16478
rect 7641 16406 7656 16478
rect 7580 16354 7592 16406
rect 7644 16354 7656 16406
rect 7580 16282 7595 16354
rect 7641 16282 7656 16354
rect 7580 16230 7592 16282
rect 7644 16230 7656 16282
rect 7580 16158 7595 16230
rect 7641 16158 7656 16230
rect 7580 16106 7592 16158
rect 7644 16106 7656 16158
rect 7580 16034 7595 16106
rect 7641 16034 7656 16106
rect 7580 15982 7592 16034
rect 7644 15982 7656 16034
rect 7580 15910 7595 15982
rect 7641 15910 7656 15982
rect 7580 15858 7592 15910
rect 7644 15858 7656 15910
rect 7580 15786 7595 15858
rect 7641 15786 7656 15858
rect 7580 15734 7592 15786
rect 7644 15734 7656 15786
rect 7580 15662 7595 15734
rect 7641 15662 7656 15734
rect 7580 15610 7592 15662
rect 7644 15610 7656 15662
rect 7580 15538 7595 15610
rect 7641 15538 7656 15610
rect 7580 15486 7592 15538
rect 7644 15486 7656 15538
rect 7580 15474 7595 15486
rect 7417 14996 7432 15008
rect 7356 14944 7368 14996
rect 7420 14944 7432 14996
rect 7356 14872 7371 14944
rect 7417 14872 7432 14944
rect 7356 14820 7368 14872
rect 7420 14820 7432 14872
rect 7356 14748 7371 14820
rect 7417 14748 7432 14820
rect 7356 14696 7368 14748
rect 7420 14696 7432 14748
rect 7356 14624 7371 14696
rect 7417 14624 7432 14696
rect 7356 14572 7368 14624
rect 7420 14572 7432 14624
rect 7356 14500 7371 14572
rect 7417 14500 7432 14572
rect 7356 14448 7368 14500
rect 7420 14448 7432 14500
rect 7356 14376 7371 14448
rect 7417 14376 7432 14448
rect 7356 14324 7368 14376
rect 7420 14324 7432 14376
rect 7356 14252 7371 14324
rect 7417 14252 7432 14324
rect 7356 14200 7368 14252
rect 7420 14200 7432 14252
rect 7356 14128 7371 14200
rect 7417 14128 7432 14200
rect 7356 14076 7368 14128
rect 7420 14076 7432 14128
rect 7356 14004 7371 14076
rect 7417 14004 7432 14076
rect 7356 13952 7368 14004
rect 7420 13952 7432 14004
rect 7356 13880 7371 13952
rect 7417 13880 7432 13952
rect 7356 13828 7368 13880
rect 7420 13828 7432 13880
rect 7356 13756 7371 13828
rect 7417 13756 7432 13828
rect 7356 13704 7368 13756
rect 7420 13704 7432 13756
rect 7356 13632 7371 13704
rect 7417 13632 7432 13704
rect 7356 13580 7368 13632
rect 7420 13580 7432 13632
rect 7356 13508 7371 13580
rect 7417 13508 7432 13580
rect 7356 13456 7368 13508
rect 7420 13456 7432 13508
rect 7356 13384 7371 13456
rect 7417 13384 7432 13456
rect 7356 13332 7368 13384
rect 7420 13332 7432 13384
rect 7356 13260 7371 13332
rect 7417 13260 7432 13332
rect 7356 13208 7368 13260
rect 7420 13208 7432 13260
rect 7356 13136 7371 13208
rect 7417 13136 7432 13208
rect 7356 13084 7368 13136
rect 7420 13084 7432 13136
rect 7356 13012 7371 13084
rect 7417 13012 7432 13084
rect 7356 12960 7368 13012
rect 7420 12960 7432 13012
rect 7356 12888 7371 12960
rect 7417 12888 7432 12960
rect 7356 12836 7368 12888
rect 7420 12836 7432 12888
rect 7356 12824 7371 12836
rect 7147 12274 7193 12598
rect 7417 12824 7432 12836
rect 7371 12585 7417 12598
rect 7641 15474 7656 15486
rect 7819 16572 7865 16585
rect 7595 12585 7641 12598
rect 8043 16572 8089 16585
rect 8028 14996 8043 15008
rect 8252 16572 8328 16602
rect 8700 16654 8776 16682
rect 8700 16602 8712 16654
rect 8764 16602 8776 16654
rect 8252 16530 8267 16572
rect 8313 16530 8328 16572
rect 8252 16478 8264 16530
rect 8316 16478 8328 16530
rect 8252 16406 8267 16478
rect 8313 16406 8328 16478
rect 8252 16354 8264 16406
rect 8316 16354 8328 16406
rect 8252 16282 8267 16354
rect 8313 16282 8328 16354
rect 8252 16230 8264 16282
rect 8316 16230 8328 16282
rect 8252 16158 8267 16230
rect 8313 16158 8328 16230
rect 8252 16106 8264 16158
rect 8316 16106 8328 16158
rect 8252 16034 8267 16106
rect 8313 16034 8328 16106
rect 8252 15982 8264 16034
rect 8316 15982 8328 16034
rect 8252 15910 8267 15982
rect 8313 15910 8328 15982
rect 8252 15858 8264 15910
rect 8316 15858 8328 15910
rect 8252 15786 8267 15858
rect 8313 15786 8328 15858
rect 8252 15734 8264 15786
rect 8316 15734 8328 15786
rect 8252 15662 8267 15734
rect 8313 15662 8328 15734
rect 8252 15610 8264 15662
rect 8316 15610 8328 15662
rect 8252 15538 8267 15610
rect 8313 15538 8328 15610
rect 8252 15486 8264 15538
rect 8316 15486 8328 15538
rect 8252 15474 8267 15486
rect 8089 14996 8104 15008
rect 8028 14944 8040 14996
rect 8092 14944 8104 14996
rect 8028 14872 8043 14944
rect 8089 14872 8104 14944
rect 8028 14820 8040 14872
rect 8092 14820 8104 14872
rect 8028 14748 8043 14820
rect 8089 14748 8104 14820
rect 8028 14696 8040 14748
rect 8092 14696 8104 14748
rect 8028 14624 8043 14696
rect 8089 14624 8104 14696
rect 8028 14572 8040 14624
rect 8092 14572 8104 14624
rect 8028 14500 8043 14572
rect 8089 14500 8104 14572
rect 8028 14448 8040 14500
rect 8092 14448 8104 14500
rect 8028 14376 8043 14448
rect 8089 14376 8104 14448
rect 8028 14324 8040 14376
rect 8092 14324 8104 14376
rect 8028 14252 8043 14324
rect 8089 14252 8104 14324
rect 8028 14200 8040 14252
rect 8092 14200 8104 14252
rect 8028 14128 8043 14200
rect 8089 14128 8104 14200
rect 8028 14076 8040 14128
rect 8092 14076 8104 14128
rect 8028 14004 8043 14076
rect 8089 14004 8104 14076
rect 8028 13952 8040 14004
rect 8092 13952 8104 14004
rect 8028 13880 8043 13952
rect 8089 13880 8104 13952
rect 8028 13828 8040 13880
rect 8092 13828 8104 13880
rect 8028 13756 8043 13828
rect 8089 13756 8104 13828
rect 8028 13704 8040 13756
rect 8092 13704 8104 13756
rect 8028 13632 8043 13704
rect 8089 13632 8104 13704
rect 8028 13580 8040 13632
rect 8092 13580 8104 13632
rect 8028 13508 8043 13580
rect 8089 13508 8104 13580
rect 8028 13456 8040 13508
rect 8092 13456 8104 13508
rect 8028 13384 8043 13456
rect 8089 13384 8104 13456
rect 8028 13332 8040 13384
rect 8092 13332 8104 13384
rect 8028 13260 8043 13332
rect 8089 13260 8104 13332
rect 8028 13208 8040 13260
rect 8092 13208 8104 13260
rect 8028 13136 8043 13208
rect 8089 13136 8104 13208
rect 8028 13084 8040 13136
rect 8092 13084 8104 13136
rect 8028 13012 8043 13084
rect 8089 13012 8104 13084
rect 8028 12960 8040 13012
rect 8092 12960 8104 13012
rect 8028 12888 8043 12960
rect 8089 12888 8104 12960
rect 8028 12836 8040 12888
rect 8092 12836 8104 12888
rect 8028 12824 8043 12836
rect 7385 12458 7547 12469
rect 7385 12412 7396 12458
rect 7536 12412 7547 12458
rect 7385 12401 7547 12412
rect 7678 12427 7746 12438
rect 7055 12263 7311 12274
rect 7055 12217 7066 12263
rect 7300 12217 7311 12263
rect 7055 12206 7311 12217
rect 7482 11958 7528 12401
rect 7678 12381 7689 12427
rect 7735 12381 7746 12427
rect 6699 11947 7547 11958
rect 6699 11901 7396 11947
rect 7536 11901 7547 11947
rect 7678 11923 7746 12381
rect 6699 11890 7547 11901
rect 7596 11911 7746 11923
rect 5788 11758 5864 11770
rect 5788 11706 5800 11758
rect 5852 11706 5864 11758
rect 5788 11634 5803 11706
rect 5849 11634 5864 11706
rect 5788 11582 5800 11634
rect 5852 11582 5864 11634
rect 5788 11510 5803 11582
rect 5849 11510 5864 11582
rect 5788 11458 5800 11510
rect 5852 11458 5864 11510
rect 5788 11446 5803 11458
rect 5579 10940 5625 10997
rect 5579 10837 5625 10894
rect 5579 10734 5625 10791
rect 5579 10631 5625 10688
rect 5579 10528 5625 10585
rect 5579 10425 5625 10482
rect 5579 10322 5625 10379
rect 5579 10219 5625 10276
rect 5579 10116 5625 10173
rect 5401 10070 5436 10109
rect 5321 10013 5436 10070
rect 5321 9967 5355 10013
rect 5401 9967 5436 10013
rect 5321 9863 5436 9967
rect 5579 10013 5625 10070
rect 5579 9954 5625 9967
rect 5849 11446 5864 11458
rect 6027 11757 6073 11770
rect 5803 10940 5849 10997
rect 5803 10837 5849 10894
rect 5803 10734 5849 10791
rect 5803 10631 5849 10688
rect 5803 10528 5849 10585
rect 5803 10425 5849 10482
rect 5803 10322 5849 10379
rect 5803 10219 5849 10276
rect 5803 10116 5849 10173
rect 6236 11758 6312 11770
rect 6236 11706 6248 11758
rect 6300 11706 6312 11758
rect 6236 11634 6251 11706
rect 6297 11634 6312 11706
rect 6236 11582 6248 11634
rect 6300 11582 6312 11634
rect 6236 11510 6251 11582
rect 6297 11510 6312 11582
rect 6236 11458 6248 11510
rect 6300 11458 6312 11510
rect 6236 11446 6251 11458
rect 6027 10940 6073 10997
rect 6027 10837 6073 10894
rect 6027 10734 6073 10791
rect 6027 10631 6073 10688
rect 6027 10528 6073 10585
rect 6027 10425 6073 10482
rect 6027 10322 6073 10379
rect 6027 10219 6073 10276
rect 6027 10116 6073 10173
rect 5803 10013 5849 10070
rect 5803 9954 5849 9967
rect 5993 10070 6027 10109
rect 6297 11446 6312 11458
rect 6475 11757 6521 11770
rect 6251 10940 6297 10997
rect 6251 10837 6297 10894
rect 6251 10734 6297 10791
rect 6251 10631 6297 10688
rect 6251 10528 6297 10585
rect 6251 10425 6297 10482
rect 6251 10322 6297 10379
rect 6251 10219 6297 10276
rect 6251 10116 6297 10173
rect 6073 10070 6108 10109
rect 5993 10013 6108 10070
rect 5993 9967 6027 10013
rect 6073 9967 6108 10013
rect 5993 9863 6108 9967
rect 6475 10940 6521 10997
rect 6475 10837 6521 10894
rect 6475 10734 6521 10791
rect 6475 10631 6521 10688
rect 6475 10528 6521 10585
rect 6475 10425 6521 10482
rect 6475 10322 6521 10379
rect 6475 10219 6521 10276
rect 6475 10116 6521 10173
rect 6251 10013 6297 10070
rect 6251 9954 6297 9967
rect 6441 10070 6475 10109
rect 6699 11757 6745 11890
rect 7596 11859 7608 11911
rect 7660 11905 7746 11911
rect 7660 11859 7689 11905
rect 7735 11859 7746 11905
rect 7596 11840 7746 11859
rect 7819 11958 7865 12598
rect 8089 12824 8104 12836
rect 8043 12585 8089 12598
rect 8313 15474 8328 15486
rect 8491 16572 8537 16585
rect 8476 14996 8491 15008
rect 8700 16572 8776 16602
rect 9372 16654 9448 16682
rect 9372 16602 9384 16654
rect 9436 16602 9448 16654
rect 8700 16530 8715 16572
rect 8761 16530 8776 16572
rect 8700 16478 8712 16530
rect 8764 16478 8776 16530
rect 8700 16406 8715 16478
rect 8761 16406 8776 16478
rect 8700 16354 8712 16406
rect 8764 16354 8776 16406
rect 8700 16282 8715 16354
rect 8761 16282 8776 16354
rect 8700 16230 8712 16282
rect 8764 16230 8776 16282
rect 8700 16158 8715 16230
rect 8761 16158 8776 16230
rect 8700 16106 8712 16158
rect 8764 16106 8776 16158
rect 8700 16034 8715 16106
rect 8761 16034 8776 16106
rect 8700 15982 8712 16034
rect 8764 15982 8776 16034
rect 8700 15910 8715 15982
rect 8761 15910 8776 15982
rect 8700 15858 8712 15910
rect 8764 15858 8776 15910
rect 8700 15786 8715 15858
rect 8761 15786 8776 15858
rect 8700 15734 8712 15786
rect 8764 15734 8776 15786
rect 8700 15662 8715 15734
rect 8761 15662 8776 15734
rect 8700 15610 8712 15662
rect 8764 15610 8776 15662
rect 8700 15538 8715 15610
rect 8761 15538 8776 15610
rect 8700 15486 8712 15538
rect 8764 15486 8776 15538
rect 8700 15474 8715 15486
rect 8537 14996 8552 15008
rect 8476 14944 8488 14996
rect 8540 14944 8552 14996
rect 8476 14872 8491 14944
rect 8537 14872 8552 14944
rect 8476 14820 8488 14872
rect 8540 14820 8552 14872
rect 8476 14748 8491 14820
rect 8537 14748 8552 14820
rect 8476 14696 8488 14748
rect 8540 14696 8552 14748
rect 8476 14624 8491 14696
rect 8537 14624 8552 14696
rect 8476 14572 8488 14624
rect 8540 14572 8552 14624
rect 8476 14500 8491 14572
rect 8537 14500 8552 14572
rect 8476 14448 8488 14500
rect 8540 14448 8552 14500
rect 8476 14376 8491 14448
rect 8537 14376 8552 14448
rect 8476 14324 8488 14376
rect 8540 14324 8552 14376
rect 8476 14252 8491 14324
rect 8537 14252 8552 14324
rect 8476 14200 8488 14252
rect 8540 14200 8552 14252
rect 8476 14128 8491 14200
rect 8537 14128 8552 14200
rect 8476 14076 8488 14128
rect 8540 14076 8552 14128
rect 8476 14004 8491 14076
rect 8537 14004 8552 14076
rect 8476 13952 8488 14004
rect 8540 13952 8552 14004
rect 8476 13880 8491 13952
rect 8537 13880 8552 13952
rect 8476 13828 8488 13880
rect 8540 13828 8552 13880
rect 8476 13756 8491 13828
rect 8537 13756 8552 13828
rect 8476 13704 8488 13756
rect 8540 13704 8552 13756
rect 8476 13632 8491 13704
rect 8537 13632 8552 13704
rect 8476 13580 8488 13632
rect 8540 13580 8552 13632
rect 8476 13508 8491 13580
rect 8537 13508 8552 13580
rect 8476 13456 8488 13508
rect 8540 13456 8552 13508
rect 8476 13384 8491 13456
rect 8537 13384 8552 13456
rect 8476 13332 8488 13384
rect 8540 13332 8552 13384
rect 8476 13260 8491 13332
rect 8537 13260 8552 13332
rect 8476 13208 8488 13260
rect 8540 13208 8552 13260
rect 8476 13136 8491 13208
rect 8537 13136 8552 13208
rect 8476 13084 8488 13136
rect 8540 13084 8552 13136
rect 8476 13012 8491 13084
rect 8537 13012 8552 13084
rect 8476 12960 8488 13012
rect 8540 12960 8552 13012
rect 8476 12888 8491 12960
rect 8537 12888 8552 12960
rect 8476 12836 8488 12888
rect 8540 12836 8552 12888
rect 8476 12824 8491 12836
rect 8267 12274 8313 12598
rect 8537 12824 8552 12836
rect 8491 12585 8537 12598
rect 8761 15474 8776 15486
rect 8939 16572 8985 16585
rect 8715 12585 8761 12598
rect 9163 16572 9209 16585
rect 9148 14996 9163 15008
rect 9372 16572 9448 16602
rect 9820 16654 9896 16682
rect 9820 16602 9832 16654
rect 9884 16602 9896 16654
rect 9372 16530 9387 16572
rect 9433 16530 9448 16572
rect 9372 16478 9384 16530
rect 9436 16478 9448 16530
rect 9372 16406 9387 16478
rect 9433 16406 9448 16478
rect 9372 16354 9384 16406
rect 9436 16354 9448 16406
rect 9372 16282 9387 16354
rect 9433 16282 9448 16354
rect 9372 16230 9384 16282
rect 9436 16230 9448 16282
rect 9372 16158 9387 16230
rect 9433 16158 9448 16230
rect 9372 16106 9384 16158
rect 9436 16106 9448 16158
rect 9372 16034 9387 16106
rect 9433 16034 9448 16106
rect 9372 15982 9384 16034
rect 9436 15982 9448 16034
rect 9372 15910 9387 15982
rect 9433 15910 9448 15982
rect 9372 15858 9384 15910
rect 9436 15858 9448 15910
rect 9372 15786 9387 15858
rect 9433 15786 9448 15858
rect 9372 15734 9384 15786
rect 9436 15734 9448 15786
rect 9372 15662 9387 15734
rect 9433 15662 9448 15734
rect 9372 15610 9384 15662
rect 9436 15610 9448 15662
rect 9372 15538 9387 15610
rect 9433 15538 9448 15610
rect 9372 15486 9384 15538
rect 9436 15486 9448 15538
rect 9372 15474 9387 15486
rect 9209 14996 9224 15008
rect 9148 14944 9160 14996
rect 9212 14944 9224 14996
rect 9148 14872 9163 14944
rect 9209 14872 9224 14944
rect 9148 14820 9160 14872
rect 9212 14820 9224 14872
rect 9148 14748 9163 14820
rect 9209 14748 9224 14820
rect 9148 14696 9160 14748
rect 9212 14696 9224 14748
rect 9148 14624 9163 14696
rect 9209 14624 9224 14696
rect 9148 14572 9160 14624
rect 9212 14572 9224 14624
rect 9148 14500 9163 14572
rect 9209 14500 9224 14572
rect 9148 14448 9160 14500
rect 9212 14448 9224 14500
rect 9148 14376 9163 14448
rect 9209 14376 9224 14448
rect 9148 14324 9160 14376
rect 9212 14324 9224 14376
rect 9148 14252 9163 14324
rect 9209 14252 9224 14324
rect 9148 14200 9160 14252
rect 9212 14200 9224 14252
rect 9148 14128 9163 14200
rect 9209 14128 9224 14200
rect 9148 14076 9160 14128
rect 9212 14076 9224 14128
rect 9148 14004 9163 14076
rect 9209 14004 9224 14076
rect 9148 13952 9160 14004
rect 9212 13952 9224 14004
rect 9148 13880 9163 13952
rect 9209 13880 9224 13952
rect 9148 13828 9160 13880
rect 9212 13828 9224 13880
rect 9148 13756 9163 13828
rect 9209 13756 9224 13828
rect 9148 13704 9160 13756
rect 9212 13704 9224 13756
rect 9148 13632 9163 13704
rect 9209 13632 9224 13704
rect 9148 13580 9160 13632
rect 9212 13580 9224 13632
rect 9148 13508 9163 13580
rect 9209 13508 9224 13580
rect 9148 13456 9160 13508
rect 9212 13456 9224 13508
rect 9148 13384 9163 13456
rect 9209 13384 9224 13456
rect 9148 13332 9160 13384
rect 9212 13332 9224 13384
rect 9148 13260 9163 13332
rect 9209 13260 9224 13332
rect 9148 13208 9160 13260
rect 9212 13208 9224 13260
rect 9148 13136 9163 13208
rect 9209 13136 9224 13208
rect 9148 13084 9160 13136
rect 9212 13084 9224 13136
rect 9148 13012 9163 13084
rect 9209 13012 9224 13084
rect 9148 12960 9160 13012
rect 9212 12960 9224 13012
rect 9148 12888 9163 12960
rect 9209 12888 9224 12960
rect 9148 12836 9160 12888
rect 9212 12836 9224 12888
rect 9148 12824 9163 12836
rect 8505 12458 8667 12469
rect 8505 12412 8516 12458
rect 8656 12412 8667 12458
rect 8505 12401 8667 12412
rect 8798 12427 8866 12438
rect 8175 12263 8431 12274
rect 8175 12217 8186 12263
rect 8420 12217 8431 12263
rect 8175 12206 8431 12217
rect 8602 11958 8648 12401
rect 8798 12381 8809 12427
rect 8855 12381 8866 12427
rect 7819 11947 8667 11958
rect 7819 11901 8516 11947
rect 8656 11901 8667 11947
rect 8798 11923 8866 12381
rect 7819 11890 8667 11901
rect 8716 11911 8866 11923
rect 6908 11758 6984 11770
rect 6908 11706 6920 11758
rect 6972 11706 6984 11758
rect 6908 11634 6923 11706
rect 6969 11634 6984 11706
rect 6908 11582 6920 11634
rect 6972 11582 6984 11634
rect 6908 11510 6923 11582
rect 6969 11510 6984 11582
rect 6908 11458 6920 11510
rect 6972 11458 6984 11510
rect 6908 11446 6923 11458
rect 6699 10940 6745 10997
rect 6699 10837 6745 10894
rect 6699 10734 6745 10791
rect 6699 10631 6745 10688
rect 6699 10528 6745 10585
rect 6699 10425 6745 10482
rect 6699 10322 6745 10379
rect 6699 10219 6745 10276
rect 6699 10116 6745 10173
rect 6521 10070 6556 10109
rect 6441 10013 6556 10070
rect 6441 9967 6475 10013
rect 6521 9967 6556 10013
rect 6441 9863 6556 9967
rect 6699 10013 6745 10070
rect 6699 9954 6745 9967
rect 6969 11446 6984 11458
rect 7147 11757 7193 11770
rect 6923 10940 6969 10997
rect 6923 10837 6969 10894
rect 6923 10734 6969 10791
rect 6923 10631 6969 10688
rect 6923 10528 6969 10585
rect 6923 10425 6969 10482
rect 6923 10322 6969 10379
rect 6923 10219 6969 10276
rect 6923 10116 6969 10173
rect 7356 11758 7432 11770
rect 7356 11706 7368 11758
rect 7420 11706 7432 11758
rect 7356 11634 7371 11706
rect 7417 11634 7432 11706
rect 7356 11582 7368 11634
rect 7420 11582 7432 11634
rect 7356 11510 7371 11582
rect 7417 11510 7432 11582
rect 7356 11458 7368 11510
rect 7420 11458 7432 11510
rect 7356 11446 7371 11458
rect 7147 10940 7193 10997
rect 7147 10837 7193 10894
rect 7147 10734 7193 10791
rect 7147 10631 7193 10688
rect 7147 10528 7193 10585
rect 7147 10425 7193 10482
rect 7147 10322 7193 10379
rect 7147 10219 7193 10276
rect 7147 10116 7193 10173
rect 6923 10013 6969 10070
rect 6923 9954 6969 9967
rect 7113 10070 7147 10109
rect 7417 11446 7432 11458
rect 7595 11757 7641 11770
rect 7371 10940 7417 10997
rect 7371 10837 7417 10894
rect 7371 10734 7417 10791
rect 7371 10631 7417 10688
rect 7371 10528 7417 10585
rect 7371 10425 7417 10482
rect 7371 10322 7417 10379
rect 7371 10219 7417 10276
rect 7371 10116 7417 10173
rect 7193 10070 7228 10109
rect 7113 10013 7228 10070
rect 7113 9967 7147 10013
rect 7193 9967 7228 10013
rect 7113 9863 7228 9967
rect 7595 10940 7641 10997
rect 7595 10837 7641 10894
rect 7595 10734 7641 10791
rect 7595 10631 7641 10688
rect 7595 10528 7641 10585
rect 7595 10425 7641 10482
rect 7595 10322 7641 10379
rect 7595 10219 7641 10276
rect 7595 10116 7641 10173
rect 7371 10013 7417 10070
rect 7371 9954 7417 9967
rect 7561 10070 7595 10109
rect 7819 11757 7865 11890
rect 8716 11859 8728 11911
rect 8780 11905 8866 11911
rect 8780 11859 8809 11905
rect 8855 11859 8866 11905
rect 8716 11840 8866 11859
rect 8939 11958 8985 12598
rect 9209 12824 9224 12836
rect 9163 12585 9209 12598
rect 9433 15474 9448 15486
rect 9611 16572 9657 16585
rect 9596 14996 9611 15008
rect 9820 16572 9896 16602
rect 10492 16654 10568 16682
rect 10492 16602 10504 16654
rect 10556 16602 10568 16654
rect 9820 16530 9835 16572
rect 9881 16530 9896 16572
rect 9820 16478 9832 16530
rect 9884 16478 9896 16530
rect 9820 16406 9835 16478
rect 9881 16406 9896 16478
rect 9820 16354 9832 16406
rect 9884 16354 9896 16406
rect 9820 16282 9835 16354
rect 9881 16282 9896 16354
rect 9820 16230 9832 16282
rect 9884 16230 9896 16282
rect 9820 16158 9835 16230
rect 9881 16158 9896 16230
rect 9820 16106 9832 16158
rect 9884 16106 9896 16158
rect 9820 16034 9835 16106
rect 9881 16034 9896 16106
rect 9820 15982 9832 16034
rect 9884 15982 9896 16034
rect 9820 15910 9835 15982
rect 9881 15910 9896 15982
rect 9820 15858 9832 15910
rect 9884 15858 9896 15910
rect 9820 15786 9835 15858
rect 9881 15786 9896 15858
rect 9820 15734 9832 15786
rect 9884 15734 9896 15786
rect 9820 15662 9835 15734
rect 9881 15662 9896 15734
rect 9820 15610 9832 15662
rect 9884 15610 9896 15662
rect 9820 15538 9835 15610
rect 9881 15538 9896 15610
rect 9820 15486 9832 15538
rect 9884 15486 9896 15538
rect 9820 15474 9835 15486
rect 9657 14996 9672 15008
rect 9596 14944 9608 14996
rect 9660 14944 9672 14996
rect 9596 14872 9611 14944
rect 9657 14872 9672 14944
rect 9596 14820 9608 14872
rect 9660 14820 9672 14872
rect 9596 14748 9611 14820
rect 9657 14748 9672 14820
rect 9596 14696 9608 14748
rect 9660 14696 9672 14748
rect 9596 14624 9611 14696
rect 9657 14624 9672 14696
rect 9596 14572 9608 14624
rect 9660 14572 9672 14624
rect 9596 14500 9611 14572
rect 9657 14500 9672 14572
rect 9596 14448 9608 14500
rect 9660 14448 9672 14500
rect 9596 14376 9611 14448
rect 9657 14376 9672 14448
rect 9596 14324 9608 14376
rect 9660 14324 9672 14376
rect 9596 14252 9611 14324
rect 9657 14252 9672 14324
rect 9596 14200 9608 14252
rect 9660 14200 9672 14252
rect 9596 14128 9611 14200
rect 9657 14128 9672 14200
rect 9596 14076 9608 14128
rect 9660 14076 9672 14128
rect 9596 14004 9611 14076
rect 9657 14004 9672 14076
rect 9596 13952 9608 14004
rect 9660 13952 9672 14004
rect 9596 13880 9611 13952
rect 9657 13880 9672 13952
rect 9596 13828 9608 13880
rect 9660 13828 9672 13880
rect 9596 13756 9611 13828
rect 9657 13756 9672 13828
rect 9596 13704 9608 13756
rect 9660 13704 9672 13756
rect 9596 13632 9611 13704
rect 9657 13632 9672 13704
rect 9596 13580 9608 13632
rect 9660 13580 9672 13632
rect 9596 13508 9611 13580
rect 9657 13508 9672 13580
rect 9596 13456 9608 13508
rect 9660 13456 9672 13508
rect 9596 13384 9611 13456
rect 9657 13384 9672 13456
rect 9596 13332 9608 13384
rect 9660 13332 9672 13384
rect 9596 13260 9611 13332
rect 9657 13260 9672 13332
rect 9596 13208 9608 13260
rect 9660 13208 9672 13260
rect 9596 13136 9611 13208
rect 9657 13136 9672 13208
rect 9596 13084 9608 13136
rect 9660 13084 9672 13136
rect 9596 13012 9611 13084
rect 9657 13012 9672 13084
rect 9596 12960 9608 13012
rect 9660 12960 9672 13012
rect 9596 12888 9611 12960
rect 9657 12888 9672 12960
rect 9596 12836 9608 12888
rect 9660 12836 9672 12888
rect 9596 12824 9611 12836
rect 9387 12274 9433 12598
rect 9657 12824 9672 12836
rect 9611 12585 9657 12598
rect 9881 15474 9896 15486
rect 10059 16572 10105 16585
rect 9835 12585 9881 12598
rect 10283 16572 10329 16585
rect 10268 14996 10283 15008
rect 10492 16572 10568 16602
rect 10940 16654 11016 16682
rect 10940 16602 10952 16654
rect 11004 16602 11016 16654
rect 10492 16530 10507 16572
rect 10553 16530 10568 16572
rect 10492 16478 10504 16530
rect 10556 16478 10568 16530
rect 10492 16406 10507 16478
rect 10553 16406 10568 16478
rect 10492 16354 10504 16406
rect 10556 16354 10568 16406
rect 10492 16282 10507 16354
rect 10553 16282 10568 16354
rect 10492 16230 10504 16282
rect 10556 16230 10568 16282
rect 10492 16158 10507 16230
rect 10553 16158 10568 16230
rect 10492 16106 10504 16158
rect 10556 16106 10568 16158
rect 10492 16034 10507 16106
rect 10553 16034 10568 16106
rect 10492 15982 10504 16034
rect 10556 15982 10568 16034
rect 10492 15910 10507 15982
rect 10553 15910 10568 15982
rect 10492 15858 10504 15910
rect 10556 15858 10568 15910
rect 10492 15786 10507 15858
rect 10553 15786 10568 15858
rect 10492 15734 10504 15786
rect 10556 15734 10568 15786
rect 10492 15662 10507 15734
rect 10553 15662 10568 15734
rect 10492 15610 10504 15662
rect 10556 15610 10568 15662
rect 10492 15538 10507 15610
rect 10553 15538 10568 15610
rect 10492 15486 10504 15538
rect 10556 15486 10568 15538
rect 10492 15474 10507 15486
rect 10329 14996 10344 15008
rect 10268 14944 10280 14996
rect 10332 14944 10344 14996
rect 10268 14872 10283 14944
rect 10329 14872 10344 14944
rect 10268 14820 10280 14872
rect 10332 14820 10344 14872
rect 10268 14748 10283 14820
rect 10329 14748 10344 14820
rect 10268 14696 10280 14748
rect 10332 14696 10344 14748
rect 10268 14624 10283 14696
rect 10329 14624 10344 14696
rect 10268 14572 10280 14624
rect 10332 14572 10344 14624
rect 10268 14500 10283 14572
rect 10329 14500 10344 14572
rect 10268 14448 10280 14500
rect 10332 14448 10344 14500
rect 10268 14376 10283 14448
rect 10329 14376 10344 14448
rect 10268 14324 10280 14376
rect 10332 14324 10344 14376
rect 10268 14252 10283 14324
rect 10329 14252 10344 14324
rect 10268 14200 10280 14252
rect 10332 14200 10344 14252
rect 10268 14128 10283 14200
rect 10329 14128 10344 14200
rect 10268 14076 10280 14128
rect 10332 14076 10344 14128
rect 10268 14004 10283 14076
rect 10329 14004 10344 14076
rect 10268 13952 10280 14004
rect 10332 13952 10344 14004
rect 10268 13880 10283 13952
rect 10329 13880 10344 13952
rect 10268 13828 10280 13880
rect 10332 13828 10344 13880
rect 10268 13756 10283 13828
rect 10329 13756 10344 13828
rect 10268 13704 10280 13756
rect 10332 13704 10344 13756
rect 10268 13632 10283 13704
rect 10329 13632 10344 13704
rect 10268 13580 10280 13632
rect 10332 13580 10344 13632
rect 10268 13508 10283 13580
rect 10329 13508 10344 13580
rect 10268 13456 10280 13508
rect 10332 13456 10344 13508
rect 10268 13384 10283 13456
rect 10329 13384 10344 13456
rect 10268 13332 10280 13384
rect 10332 13332 10344 13384
rect 10268 13260 10283 13332
rect 10329 13260 10344 13332
rect 10268 13208 10280 13260
rect 10332 13208 10344 13260
rect 10268 13136 10283 13208
rect 10329 13136 10344 13208
rect 10268 13084 10280 13136
rect 10332 13084 10344 13136
rect 10268 13012 10283 13084
rect 10329 13012 10344 13084
rect 10268 12960 10280 13012
rect 10332 12960 10344 13012
rect 10268 12888 10283 12960
rect 10329 12888 10344 12960
rect 10268 12836 10280 12888
rect 10332 12836 10344 12888
rect 10268 12824 10283 12836
rect 9625 12458 9787 12469
rect 9625 12412 9636 12458
rect 9776 12412 9787 12458
rect 9625 12401 9787 12412
rect 9918 12427 9986 12438
rect 9295 12263 9551 12274
rect 9295 12217 9306 12263
rect 9540 12217 9551 12263
rect 9295 12206 9551 12217
rect 9722 11958 9768 12401
rect 9918 12381 9929 12427
rect 9975 12381 9986 12427
rect 8939 11947 9787 11958
rect 8939 11901 9636 11947
rect 9776 11901 9787 11947
rect 9918 11923 9986 12381
rect 8939 11890 9787 11901
rect 9836 11911 9986 11923
rect 8028 11758 8104 11770
rect 8028 11706 8040 11758
rect 8092 11706 8104 11758
rect 8028 11634 8043 11706
rect 8089 11634 8104 11706
rect 8028 11582 8040 11634
rect 8092 11582 8104 11634
rect 8028 11510 8043 11582
rect 8089 11510 8104 11582
rect 8028 11458 8040 11510
rect 8092 11458 8104 11510
rect 8028 11446 8043 11458
rect 7819 10940 7865 10997
rect 7819 10837 7865 10894
rect 7819 10734 7865 10791
rect 7819 10631 7865 10688
rect 7819 10528 7865 10585
rect 7819 10425 7865 10482
rect 7819 10322 7865 10379
rect 7819 10219 7865 10276
rect 7819 10116 7865 10173
rect 7641 10070 7676 10109
rect 7561 10013 7676 10070
rect 7561 9967 7595 10013
rect 7641 9967 7676 10013
rect 7561 9863 7676 9967
rect 7819 10013 7865 10070
rect 7819 9954 7865 9967
rect 8089 11446 8104 11458
rect 8267 11757 8313 11770
rect 8043 10940 8089 10997
rect 8043 10837 8089 10894
rect 8043 10734 8089 10791
rect 8043 10631 8089 10688
rect 8043 10528 8089 10585
rect 8043 10425 8089 10482
rect 8043 10322 8089 10379
rect 8043 10219 8089 10276
rect 8043 10116 8089 10173
rect 8476 11758 8552 11770
rect 8476 11706 8488 11758
rect 8540 11706 8552 11758
rect 8476 11634 8491 11706
rect 8537 11634 8552 11706
rect 8476 11582 8488 11634
rect 8540 11582 8552 11634
rect 8476 11510 8491 11582
rect 8537 11510 8552 11582
rect 8476 11458 8488 11510
rect 8540 11458 8552 11510
rect 8476 11446 8491 11458
rect 8267 10940 8313 10997
rect 8267 10837 8313 10894
rect 8267 10734 8313 10791
rect 8267 10631 8313 10688
rect 8267 10528 8313 10585
rect 8267 10425 8313 10482
rect 8267 10322 8313 10379
rect 8267 10219 8313 10276
rect 8267 10116 8313 10173
rect 8043 10013 8089 10070
rect 8043 9954 8089 9967
rect 8233 10070 8267 10109
rect 8537 11446 8552 11458
rect 8715 11757 8761 11770
rect 8491 10940 8537 10997
rect 8491 10837 8537 10894
rect 8491 10734 8537 10791
rect 8491 10631 8537 10688
rect 8491 10528 8537 10585
rect 8491 10425 8537 10482
rect 8491 10322 8537 10379
rect 8491 10219 8537 10276
rect 8491 10116 8537 10173
rect 8313 10070 8348 10109
rect 8233 10013 8348 10070
rect 8233 9967 8267 10013
rect 8313 9967 8348 10013
rect 8233 9863 8348 9967
rect 8715 10940 8761 10997
rect 8715 10837 8761 10894
rect 8715 10734 8761 10791
rect 8715 10631 8761 10688
rect 8715 10528 8761 10585
rect 8715 10425 8761 10482
rect 8715 10322 8761 10379
rect 8715 10219 8761 10276
rect 8715 10116 8761 10173
rect 8491 10013 8537 10070
rect 8491 9954 8537 9967
rect 8681 10070 8715 10109
rect 8939 11757 8985 11890
rect 9836 11859 9848 11911
rect 9900 11905 9986 11911
rect 9900 11859 9929 11905
rect 9975 11859 9986 11905
rect 9836 11840 9986 11859
rect 10059 11958 10105 12598
rect 10329 12824 10344 12836
rect 10283 12585 10329 12598
rect 10553 15474 10568 15486
rect 10731 16572 10777 16585
rect 10716 14996 10731 15008
rect 10940 16572 11016 16602
rect 11612 16654 11688 16682
rect 11612 16602 11624 16654
rect 11676 16602 11688 16654
rect 10940 16530 10955 16572
rect 11001 16530 11016 16572
rect 10940 16478 10952 16530
rect 11004 16478 11016 16530
rect 10940 16406 10955 16478
rect 11001 16406 11016 16478
rect 10940 16354 10952 16406
rect 11004 16354 11016 16406
rect 10940 16282 10955 16354
rect 11001 16282 11016 16354
rect 10940 16230 10952 16282
rect 11004 16230 11016 16282
rect 10940 16158 10955 16230
rect 11001 16158 11016 16230
rect 10940 16106 10952 16158
rect 11004 16106 11016 16158
rect 10940 16034 10955 16106
rect 11001 16034 11016 16106
rect 10940 15982 10952 16034
rect 11004 15982 11016 16034
rect 10940 15910 10955 15982
rect 11001 15910 11016 15982
rect 10940 15858 10952 15910
rect 11004 15858 11016 15910
rect 10940 15786 10955 15858
rect 11001 15786 11016 15858
rect 10940 15734 10952 15786
rect 11004 15734 11016 15786
rect 10940 15662 10955 15734
rect 11001 15662 11016 15734
rect 10940 15610 10952 15662
rect 11004 15610 11016 15662
rect 10940 15538 10955 15610
rect 11001 15538 11016 15610
rect 10940 15486 10952 15538
rect 11004 15486 11016 15538
rect 10940 15474 10955 15486
rect 10777 14996 10792 15008
rect 10716 14944 10728 14996
rect 10780 14944 10792 14996
rect 10716 14872 10731 14944
rect 10777 14872 10792 14944
rect 10716 14820 10728 14872
rect 10780 14820 10792 14872
rect 10716 14748 10731 14820
rect 10777 14748 10792 14820
rect 10716 14696 10728 14748
rect 10780 14696 10792 14748
rect 10716 14624 10731 14696
rect 10777 14624 10792 14696
rect 10716 14572 10728 14624
rect 10780 14572 10792 14624
rect 10716 14500 10731 14572
rect 10777 14500 10792 14572
rect 10716 14448 10728 14500
rect 10780 14448 10792 14500
rect 10716 14376 10731 14448
rect 10777 14376 10792 14448
rect 10716 14324 10728 14376
rect 10780 14324 10792 14376
rect 10716 14252 10731 14324
rect 10777 14252 10792 14324
rect 10716 14200 10728 14252
rect 10780 14200 10792 14252
rect 10716 14128 10731 14200
rect 10777 14128 10792 14200
rect 10716 14076 10728 14128
rect 10780 14076 10792 14128
rect 10716 14004 10731 14076
rect 10777 14004 10792 14076
rect 10716 13952 10728 14004
rect 10780 13952 10792 14004
rect 10716 13880 10731 13952
rect 10777 13880 10792 13952
rect 10716 13828 10728 13880
rect 10780 13828 10792 13880
rect 10716 13756 10731 13828
rect 10777 13756 10792 13828
rect 10716 13704 10728 13756
rect 10780 13704 10792 13756
rect 10716 13632 10731 13704
rect 10777 13632 10792 13704
rect 10716 13580 10728 13632
rect 10780 13580 10792 13632
rect 10716 13508 10731 13580
rect 10777 13508 10792 13580
rect 10716 13456 10728 13508
rect 10780 13456 10792 13508
rect 10716 13384 10731 13456
rect 10777 13384 10792 13456
rect 10716 13332 10728 13384
rect 10780 13332 10792 13384
rect 10716 13260 10731 13332
rect 10777 13260 10792 13332
rect 10716 13208 10728 13260
rect 10780 13208 10792 13260
rect 10716 13136 10731 13208
rect 10777 13136 10792 13208
rect 10716 13084 10728 13136
rect 10780 13084 10792 13136
rect 10716 13012 10731 13084
rect 10777 13012 10792 13084
rect 10716 12960 10728 13012
rect 10780 12960 10792 13012
rect 10716 12888 10731 12960
rect 10777 12888 10792 12960
rect 10716 12836 10728 12888
rect 10780 12836 10792 12888
rect 10716 12824 10731 12836
rect 10507 12274 10553 12598
rect 10777 12824 10792 12836
rect 10731 12585 10777 12598
rect 11001 15474 11016 15486
rect 11179 16572 11225 16585
rect 10955 12585 11001 12598
rect 11403 16572 11449 16585
rect 11388 14996 11403 15008
rect 11612 16572 11688 16602
rect 12060 16654 12136 16682
rect 12060 16602 12072 16654
rect 12124 16602 12136 16654
rect 11612 16530 11627 16572
rect 11673 16530 11688 16572
rect 11612 16478 11624 16530
rect 11676 16478 11688 16530
rect 11612 16406 11627 16478
rect 11673 16406 11688 16478
rect 11612 16354 11624 16406
rect 11676 16354 11688 16406
rect 11612 16282 11627 16354
rect 11673 16282 11688 16354
rect 11612 16230 11624 16282
rect 11676 16230 11688 16282
rect 11612 16158 11627 16230
rect 11673 16158 11688 16230
rect 11612 16106 11624 16158
rect 11676 16106 11688 16158
rect 11612 16034 11627 16106
rect 11673 16034 11688 16106
rect 11612 15982 11624 16034
rect 11676 15982 11688 16034
rect 11612 15910 11627 15982
rect 11673 15910 11688 15982
rect 11612 15858 11624 15910
rect 11676 15858 11688 15910
rect 11612 15786 11627 15858
rect 11673 15786 11688 15858
rect 11612 15734 11624 15786
rect 11676 15734 11688 15786
rect 11612 15662 11627 15734
rect 11673 15662 11688 15734
rect 11612 15610 11624 15662
rect 11676 15610 11688 15662
rect 11612 15538 11627 15610
rect 11673 15538 11688 15610
rect 11612 15486 11624 15538
rect 11676 15486 11688 15538
rect 11612 15474 11627 15486
rect 11449 14996 11464 15008
rect 11388 14944 11400 14996
rect 11452 14944 11464 14996
rect 11388 14872 11403 14944
rect 11449 14872 11464 14944
rect 11388 14820 11400 14872
rect 11452 14820 11464 14872
rect 11388 14748 11403 14820
rect 11449 14748 11464 14820
rect 11388 14696 11400 14748
rect 11452 14696 11464 14748
rect 11388 14624 11403 14696
rect 11449 14624 11464 14696
rect 11388 14572 11400 14624
rect 11452 14572 11464 14624
rect 11388 14500 11403 14572
rect 11449 14500 11464 14572
rect 11388 14448 11400 14500
rect 11452 14448 11464 14500
rect 11388 14376 11403 14448
rect 11449 14376 11464 14448
rect 11388 14324 11400 14376
rect 11452 14324 11464 14376
rect 11388 14252 11403 14324
rect 11449 14252 11464 14324
rect 11388 14200 11400 14252
rect 11452 14200 11464 14252
rect 11388 14128 11403 14200
rect 11449 14128 11464 14200
rect 11388 14076 11400 14128
rect 11452 14076 11464 14128
rect 11388 14004 11403 14076
rect 11449 14004 11464 14076
rect 11388 13952 11400 14004
rect 11452 13952 11464 14004
rect 11388 13880 11403 13952
rect 11449 13880 11464 13952
rect 11388 13828 11400 13880
rect 11452 13828 11464 13880
rect 11388 13756 11403 13828
rect 11449 13756 11464 13828
rect 11388 13704 11400 13756
rect 11452 13704 11464 13756
rect 11388 13632 11403 13704
rect 11449 13632 11464 13704
rect 11388 13580 11400 13632
rect 11452 13580 11464 13632
rect 11388 13508 11403 13580
rect 11449 13508 11464 13580
rect 11388 13456 11400 13508
rect 11452 13456 11464 13508
rect 11388 13384 11403 13456
rect 11449 13384 11464 13456
rect 11388 13332 11400 13384
rect 11452 13332 11464 13384
rect 11388 13260 11403 13332
rect 11449 13260 11464 13332
rect 11388 13208 11400 13260
rect 11452 13208 11464 13260
rect 11388 13136 11403 13208
rect 11449 13136 11464 13208
rect 11388 13084 11400 13136
rect 11452 13084 11464 13136
rect 11388 13012 11403 13084
rect 11449 13012 11464 13084
rect 11388 12960 11400 13012
rect 11452 12960 11464 13012
rect 11388 12888 11403 12960
rect 11449 12888 11464 12960
rect 11388 12836 11400 12888
rect 11452 12836 11464 12888
rect 11388 12824 11403 12836
rect 10745 12458 10907 12469
rect 10745 12412 10756 12458
rect 10896 12412 10907 12458
rect 10745 12401 10907 12412
rect 11038 12427 11106 12438
rect 10415 12263 10671 12274
rect 10415 12217 10426 12263
rect 10660 12217 10671 12263
rect 10415 12206 10671 12217
rect 10842 11958 10888 12401
rect 11038 12381 11049 12427
rect 11095 12381 11106 12427
rect 10059 11947 10907 11958
rect 10059 11901 10756 11947
rect 10896 11901 10907 11947
rect 11038 11923 11106 12381
rect 10059 11890 10907 11901
rect 10956 11911 11106 11923
rect 9148 11758 9224 11770
rect 9148 11706 9160 11758
rect 9212 11706 9224 11758
rect 9148 11634 9163 11706
rect 9209 11634 9224 11706
rect 9148 11582 9160 11634
rect 9212 11582 9224 11634
rect 9148 11510 9163 11582
rect 9209 11510 9224 11582
rect 9148 11458 9160 11510
rect 9212 11458 9224 11510
rect 9148 11446 9163 11458
rect 8939 10940 8985 10997
rect 8939 10837 8985 10894
rect 8939 10734 8985 10791
rect 8939 10631 8985 10688
rect 8939 10528 8985 10585
rect 8939 10425 8985 10482
rect 8939 10322 8985 10379
rect 8939 10219 8985 10276
rect 8939 10116 8985 10173
rect 8761 10070 8796 10109
rect 8681 10013 8796 10070
rect 8681 9967 8715 10013
rect 8761 9967 8796 10013
rect 8681 9863 8796 9967
rect 8939 10013 8985 10070
rect 8939 9954 8985 9967
rect 9209 11446 9224 11458
rect 9387 11757 9433 11770
rect 9163 10940 9209 10997
rect 9163 10837 9209 10894
rect 9163 10734 9209 10791
rect 9163 10631 9209 10688
rect 9163 10528 9209 10585
rect 9163 10425 9209 10482
rect 9163 10322 9209 10379
rect 9163 10219 9209 10276
rect 9163 10116 9209 10173
rect 9596 11758 9672 11770
rect 9596 11706 9608 11758
rect 9660 11706 9672 11758
rect 9596 11634 9611 11706
rect 9657 11634 9672 11706
rect 9596 11582 9608 11634
rect 9660 11582 9672 11634
rect 9596 11510 9611 11582
rect 9657 11510 9672 11582
rect 9596 11458 9608 11510
rect 9660 11458 9672 11510
rect 9596 11446 9611 11458
rect 9387 10940 9433 10997
rect 9387 10837 9433 10894
rect 9387 10734 9433 10791
rect 9387 10631 9433 10688
rect 9387 10528 9433 10585
rect 9387 10425 9433 10482
rect 9387 10322 9433 10379
rect 9387 10219 9433 10276
rect 9387 10116 9433 10173
rect 9163 10013 9209 10070
rect 9163 9954 9209 9967
rect 9353 10070 9387 10109
rect 9657 11446 9672 11458
rect 9835 11757 9881 11770
rect 9611 10940 9657 10997
rect 9611 10837 9657 10894
rect 9611 10734 9657 10791
rect 9611 10631 9657 10688
rect 9611 10528 9657 10585
rect 9611 10425 9657 10482
rect 9611 10322 9657 10379
rect 9611 10219 9657 10276
rect 9611 10116 9657 10173
rect 9433 10070 9468 10109
rect 9353 10013 9468 10070
rect 9353 9967 9387 10013
rect 9433 9967 9468 10013
rect 9353 9863 9468 9967
rect 9835 10940 9881 10997
rect 9835 10837 9881 10894
rect 9835 10734 9881 10791
rect 9835 10631 9881 10688
rect 9835 10528 9881 10585
rect 9835 10425 9881 10482
rect 9835 10322 9881 10379
rect 9835 10219 9881 10276
rect 9835 10116 9881 10173
rect 9611 10013 9657 10070
rect 9611 9954 9657 9967
rect 9801 10070 9835 10109
rect 10059 11757 10105 11890
rect 10956 11859 10968 11911
rect 11020 11905 11106 11911
rect 11020 11859 11049 11905
rect 11095 11859 11106 11905
rect 10956 11840 11106 11859
rect 11179 11958 11225 12598
rect 11449 12824 11464 12836
rect 11403 12585 11449 12598
rect 11673 15474 11688 15486
rect 11851 16572 11897 16585
rect 11836 14996 11851 15008
rect 12060 16572 12136 16602
rect 12732 16654 12808 16682
rect 12732 16602 12744 16654
rect 12796 16602 12808 16654
rect 12060 16530 12075 16572
rect 12121 16530 12136 16572
rect 12060 16478 12072 16530
rect 12124 16478 12136 16530
rect 12060 16406 12075 16478
rect 12121 16406 12136 16478
rect 12060 16354 12072 16406
rect 12124 16354 12136 16406
rect 12060 16282 12075 16354
rect 12121 16282 12136 16354
rect 12060 16230 12072 16282
rect 12124 16230 12136 16282
rect 12060 16158 12075 16230
rect 12121 16158 12136 16230
rect 12060 16106 12072 16158
rect 12124 16106 12136 16158
rect 12060 16034 12075 16106
rect 12121 16034 12136 16106
rect 12060 15982 12072 16034
rect 12124 15982 12136 16034
rect 12060 15910 12075 15982
rect 12121 15910 12136 15982
rect 12060 15858 12072 15910
rect 12124 15858 12136 15910
rect 12060 15786 12075 15858
rect 12121 15786 12136 15858
rect 12060 15734 12072 15786
rect 12124 15734 12136 15786
rect 12060 15662 12075 15734
rect 12121 15662 12136 15734
rect 12060 15610 12072 15662
rect 12124 15610 12136 15662
rect 12060 15538 12075 15610
rect 12121 15538 12136 15610
rect 12060 15486 12072 15538
rect 12124 15486 12136 15538
rect 12060 15474 12075 15486
rect 11897 14996 11912 15008
rect 11836 14944 11848 14996
rect 11900 14944 11912 14996
rect 11836 14872 11851 14944
rect 11897 14872 11912 14944
rect 11836 14820 11848 14872
rect 11900 14820 11912 14872
rect 11836 14748 11851 14820
rect 11897 14748 11912 14820
rect 11836 14696 11848 14748
rect 11900 14696 11912 14748
rect 11836 14624 11851 14696
rect 11897 14624 11912 14696
rect 11836 14572 11848 14624
rect 11900 14572 11912 14624
rect 11836 14500 11851 14572
rect 11897 14500 11912 14572
rect 11836 14448 11848 14500
rect 11900 14448 11912 14500
rect 11836 14376 11851 14448
rect 11897 14376 11912 14448
rect 11836 14324 11848 14376
rect 11900 14324 11912 14376
rect 11836 14252 11851 14324
rect 11897 14252 11912 14324
rect 11836 14200 11848 14252
rect 11900 14200 11912 14252
rect 11836 14128 11851 14200
rect 11897 14128 11912 14200
rect 11836 14076 11848 14128
rect 11900 14076 11912 14128
rect 11836 14004 11851 14076
rect 11897 14004 11912 14076
rect 11836 13952 11848 14004
rect 11900 13952 11912 14004
rect 11836 13880 11851 13952
rect 11897 13880 11912 13952
rect 11836 13828 11848 13880
rect 11900 13828 11912 13880
rect 11836 13756 11851 13828
rect 11897 13756 11912 13828
rect 11836 13704 11848 13756
rect 11900 13704 11912 13756
rect 11836 13632 11851 13704
rect 11897 13632 11912 13704
rect 11836 13580 11848 13632
rect 11900 13580 11912 13632
rect 11836 13508 11851 13580
rect 11897 13508 11912 13580
rect 11836 13456 11848 13508
rect 11900 13456 11912 13508
rect 11836 13384 11851 13456
rect 11897 13384 11912 13456
rect 11836 13332 11848 13384
rect 11900 13332 11912 13384
rect 11836 13260 11851 13332
rect 11897 13260 11912 13332
rect 11836 13208 11848 13260
rect 11900 13208 11912 13260
rect 11836 13136 11851 13208
rect 11897 13136 11912 13208
rect 11836 13084 11848 13136
rect 11900 13084 11912 13136
rect 11836 13012 11851 13084
rect 11897 13012 11912 13084
rect 11836 12960 11848 13012
rect 11900 12960 11912 13012
rect 11836 12888 11851 12960
rect 11897 12888 11912 12960
rect 11836 12836 11848 12888
rect 11900 12836 11912 12888
rect 11836 12824 11851 12836
rect 11627 12274 11673 12598
rect 11897 12824 11912 12836
rect 11851 12585 11897 12598
rect 12121 15474 12136 15486
rect 12299 16572 12345 16585
rect 12075 12585 12121 12598
rect 12523 16572 12569 16585
rect 12508 14996 12523 15008
rect 12732 16572 12808 16602
rect 13180 16654 13256 16682
rect 13180 16602 13192 16654
rect 13244 16602 13256 16654
rect 12732 16530 12747 16572
rect 12793 16530 12808 16572
rect 12732 16478 12744 16530
rect 12796 16478 12808 16530
rect 12732 16406 12747 16478
rect 12793 16406 12808 16478
rect 12732 16354 12744 16406
rect 12796 16354 12808 16406
rect 12732 16282 12747 16354
rect 12793 16282 12808 16354
rect 12732 16230 12744 16282
rect 12796 16230 12808 16282
rect 12732 16158 12747 16230
rect 12793 16158 12808 16230
rect 12732 16106 12744 16158
rect 12796 16106 12808 16158
rect 12732 16034 12747 16106
rect 12793 16034 12808 16106
rect 12732 15982 12744 16034
rect 12796 15982 12808 16034
rect 12732 15910 12747 15982
rect 12793 15910 12808 15982
rect 12732 15858 12744 15910
rect 12796 15858 12808 15910
rect 12732 15786 12747 15858
rect 12793 15786 12808 15858
rect 12732 15734 12744 15786
rect 12796 15734 12808 15786
rect 12732 15662 12747 15734
rect 12793 15662 12808 15734
rect 12732 15610 12744 15662
rect 12796 15610 12808 15662
rect 12732 15538 12747 15610
rect 12793 15538 12808 15610
rect 12732 15486 12744 15538
rect 12796 15486 12808 15538
rect 12732 15474 12747 15486
rect 12569 14996 12584 15008
rect 12508 14944 12520 14996
rect 12572 14944 12584 14996
rect 12508 14872 12523 14944
rect 12569 14872 12584 14944
rect 12508 14820 12520 14872
rect 12572 14820 12584 14872
rect 12508 14748 12523 14820
rect 12569 14748 12584 14820
rect 12508 14696 12520 14748
rect 12572 14696 12584 14748
rect 12508 14624 12523 14696
rect 12569 14624 12584 14696
rect 12508 14572 12520 14624
rect 12572 14572 12584 14624
rect 12508 14500 12523 14572
rect 12569 14500 12584 14572
rect 12508 14448 12520 14500
rect 12572 14448 12584 14500
rect 12508 14376 12523 14448
rect 12569 14376 12584 14448
rect 12508 14324 12520 14376
rect 12572 14324 12584 14376
rect 12508 14252 12523 14324
rect 12569 14252 12584 14324
rect 12508 14200 12520 14252
rect 12572 14200 12584 14252
rect 12508 14128 12523 14200
rect 12569 14128 12584 14200
rect 12508 14076 12520 14128
rect 12572 14076 12584 14128
rect 12508 14004 12523 14076
rect 12569 14004 12584 14076
rect 12508 13952 12520 14004
rect 12572 13952 12584 14004
rect 12508 13880 12523 13952
rect 12569 13880 12584 13952
rect 12508 13828 12520 13880
rect 12572 13828 12584 13880
rect 12508 13756 12523 13828
rect 12569 13756 12584 13828
rect 12508 13704 12520 13756
rect 12572 13704 12584 13756
rect 12508 13632 12523 13704
rect 12569 13632 12584 13704
rect 12508 13580 12520 13632
rect 12572 13580 12584 13632
rect 12508 13508 12523 13580
rect 12569 13508 12584 13580
rect 12508 13456 12520 13508
rect 12572 13456 12584 13508
rect 12508 13384 12523 13456
rect 12569 13384 12584 13456
rect 12508 13332 12520 13384
rect 12572 13332 12584 13384
rect 12508 13260 12523 13332
rect 12569 13260 12584 13332
rect 12508 13208 12520 13260
rect 12572 13208 12584 13260
rect 12508 13136 12523 13208
rect 12569 13136 12584 13208
rect 12508 13084 12520 13136
rect 12572 13084 12584 13136
rect 12508 13012 12523 13084
rect 12569 13012 12584 13084
rect 12508 12960 12520 13012
rect 12572 12960 12584 13012
rect 12508 12888 12523 12960
rect 12569 12888 12584 12960
rect 12508 12836 12520 12888
rect 12572 12836 12584 12888
rect 12508 12824 12523 12836
rect 11865 12458 12027 12469
rect 11865 12412 11876 12458
rect 12016 12412 12027 12458
rect 11865 12401 12027 12412
rect 12158 12427 12226 12438
rect 11535 12263 11791 12274
rect 11535 12217 11546 12263
rect 11780 12217 11791 12263
rect 11535 12206 11791 12217
rect 11962 11958 12008 12401
rect 12158 12381 12169 12427
rect 12215 12381 12226 12427
rect 11179 11947 12027 11958
rect 11179 11901 11876 11947
rect 12016 11901 12027 11947
rect 12158 11923 12226 12381
rect 11179 11890 12027 11901
rect 12076 11911 12226 11923
rect 10268 11758 10344 11770
rect 10268 11706 10280 11758
rect 10332 11706 10344 11758
rect 10268 11634 10283 11706
rect 10329 11634 10344 11706
rect 10268 11582 10280 11634
rect 10332 11582 10344 11634
rect 10268 11510 10283 11582
rect 10329 11510 10344 11582
rect 10268 11458 10280 11510
rect 10332 11458 10344 11510
rect 10268 11446 10283 11458
rect 10059 10940 10105 10997
rect 10059 10837 10105 10894
rect 10059 10734 10105 10791
rect 10059 10631 10105 10688
rect 10059 10528 10105 10585
rect 10059 10425 10105 10482
rect 10059 10322 10105 10379
rect 10059 10219 10105 10276
rect 10059 10116 10105 10173
rect 9881 10070 9916 10109
rect 9801 10013 9916 10070
rect 9801 9967 9835 10013
rect 9881 9967 9916 10013
rect 9801 9863 9916 9967
rect 10059 10013 10105 10070
rect 10059 9954 10105 9967
rect 10329 11446 10344 11458
rect 10507 11757 10553 11770
rect 10283 10940 10329 10997
rect 10283 10837 10329 10894
rect 10283 10734 10329 10791
rect 10283 10631 10329 10688
rect 10283 10528 10329 10585
rect 10283 10425 10329 10482
rect 10283 10322 10329 10379
rect 10283 10219 10329 10276
rect 10283 10116 10329 10173
rect 10716 11758 10792 11770
rect 10716 11706 10728 11758
rect 10780 11706 10792 11758
rect 10716 11634 10731 11706
rect 10777 11634 10792 11706
rect 10716 11582 10728 11634
rect 10780 11582 10792 11634
rect 10716 11510 10731 11582
rect 10777 11510 10792 11582
rect 10716 11458 10728 11510
rect 10780 11458 10792 11510
rect 10716 11446 10731 11458
rect 10507 10940 10553 10997
rect 10507 10837 10553 10894
rect 10507 10734 10553 10791
rect 10507 10631 10553 10688
rect 10507 10528 10553 10585
rect 10507 10425 10553 10482
rect 10507 10322 10553 10379
rect 10507 10219 10553 10276
rect 10507 10116 10553 10173
rect 10283 10013 10329 10070
rect 10283 9954 10329 9967
rect 10473 10070 10507 10109
rect 10777 11446 10792 11458
rect 10955 11757 11001 11770
rect 10731 10940 10777 10997
rect 10731 10837 10777 10894
rect 10731 10734 10777 10791
rect 10731 10631 10777 10688
rect 10731 10528 10777 10585
rect 10731 10425 10777 10482
rect 10731 10322 10777 10379
rect 10731 10219 10777 10276
rect 10731 10116 10777 10173
rect 10553 10070 10588 10109
rect 10473 10013 10588 10070
rect 10473 9967 10507 10013
rect 10553 9967 10588 10013
rect 10473 9863 10588 9967
rect 10955 10940 11001 10997
rect 10955 10837 11001 10894
rect 10955 10734 11001 10791
rect 10955 10631 11001 10688
rect 10955 10528 11001 10585
rect 10955 10425 11001 10482
rect 10955 10322 11001 10379
rect 10955 10219 11001 10276
rect 10955 10116 11001 10173
rect 10731 10013 10777 10070
rect 10731 9954 10777 9967
rect 10921 10070 10955 10109
rect 11179 11757 11225 11890
rect 12076 11859 12088 11911
rect 12140 11905 12226 11911
rect 12140 11859 12169 11905
rect 12215 11859 12226 11905
rect 12076 11840 12226 11859
rect 12299 11958 12345 12598
rect 12569 12824 12584 12836
rect 12523 12585 12569 12598
rect 12793 15474 12808 15486
rect 12971 16572 13017 16585
rect 12956 14996 12971 15008
rect 13180 16572 13256 16602
rect 13852 16654 13928 16682
rect 13852 16602 13864 16654
rect 13916 16602 13928 16654
rect 13180 16530 13195 16572
rect 13241 16530 13256 16572
rect 13180 16478 13192 16530
rect 13244 16478 13256 16530
rect 13180 16406 13195 16478
rect 13241 16406 13256 16478
rect 13180 16354 13192 16406
rect 13244 16354 13256 16406
rect 13180 16282 13195 16354
rect 13241 16282 13256 16354
rect 13180 16230 13192 16282
rect 13244 16230 13256 16282
rect 13180 16158 13195 16230
rect 13241 16158 13256 16230
rect 13180 16106 13192 16158
rect 13244 16106 13256 16158
rect 13180 16034 13195 16106
rect 13241 16034 13256 16106
rect 13180 15982 13192 16034
rect 13244 15982 13256 16034
rect 13180 15910 13195 15982
rect 13241 15910 13256 15982
rect 13180 15858 13192 15910
rect 13244 15858 13256 15910
rect 13180 15786 13195 15858
rect 13241 15786 13256 15858
rect 13180 15734 13192 15786
rect 13244 15734 13256 15786
rect 13180 15662 13195 15734
rect 13241 15662 13256 15734
rect 13180 15610 13192 15662
rect 13244 15610 13256 15662
rect 13180 15538 13195 15610
rect 13241 15538 13256 15610
rect 13180 15486 13192 15538
rect 13244 15486 13256 15538
rect 13180 15474 13195 15486
rect 13017 14996 13032 15008
rect 12956 14944 12968 14996
rect 13020 14944 13032 14996
rect 12956 14872 12971 14944
rect 13017 14872 13032 14944
rect 12956 14820 12968 14872
rect 13020 14820 13032 14872
rect 12956 14748 12971 14820
rect 13017 14748 13032 14820
rect 12956 14696 12968 14748
rect 13020 14696 13032 14748
rect 12956 14624 12971 14696
rect 13017 14624 13032 14696
rect 12956 14572 12968 14624
rect 13020 14572 13032 14624
rect 12956 14500 12971 14572
rect 13017 14500 13032 14572
rect 12956 14448 12968 14500
rect 13020 14448 13032 14500
rect 12956 14376 12971 14448
rect 13017 14376 13032 14448
rect 12956 14324 12968 14376
rect 13020 14324 13032 14376
rect 12956 14252 12971 14324
rect 13017 14252 13032 14324
rect 12956 14200 12968 14252
rect 13020 14200 13032 14252
rect 12956 14128 12971 14200
rect 13017 14128 13032 14200
rect 12956 14076 12968 14128
rect 13020 14076 13032 14128
rect 12956 14004 12971 14076
rect 13017 14004 13032 14076
rect 12956 13952 12968 14004
rect 13020 13952 13032 14004
rect 12956 13880 12971 13952
rect 13017 13880 13032 13952
rect 12956 13828 12968 13880
rect 13020 13828 13032 13880
rect 12956 13756 12971 13828
rect 13017 13756 13032 13828
rect 12956 13704 12968 13756
rect 13020 13704 13032 13756
rect 12956 13632 12971 13704
rect 13017 13632 13032 13704
rect 12956 13580 12968 13632
rect 13020 13580 13032 13632
rect 12956 13508 12971 13580
rect 13017 13508 13032 13580
rect 12956 13456 12968 13508
rect 13020 13456 13032 13508
rect 12956 13384 12971 13456
rect 13017 13384 13032 13456
rect 12956 13332 12968 13384
rect 13020 13332 13032 13384
rect 12956 13260 12971 13332
rect 13017 13260 13032 13332
rect 12956 13208 12968 13260
rect 13020 13208 13032 13260
rect 12956 13136 12971 13208
rect 13017 13136 13032 13208
rect 12956 13084 12968 13136
rect 13020 13084 13032 13136
rect 12956 13012 12971 13084
rect 13017 13012 13032 13084
rect 12956 12960 12968 13012
rect 13020 12960 13032 13012
rect 12956 12888 12971 12960
rect 13017 12888 13032 12960
rect 12956 12836 12968 12888
rect 13020 12836 13032 12888
rect 12956 12824 12971 12836
rect 12747 12274 12793 12598
rect 13017 12824 13032 12836
rect 12971 12585 13017 12598
rect 13241 15474 13256 15486
rect 13419 16572 13465 16585
rect 13195 12585 13241 12598
rect 13643 16572 13689 16585
rect 13628 14996 13643 15008
rect 13852 16572 13928 16602
rect 14300 16654 14376 16682
rect 14300 16602 14312 16654
rect 14364 16602 14376 16654
rect 13852 16530 13867 16572
rect 13913 16530 13928 16572
rect 13852 16478 13864 16530
rect 13916 16478 13928 16530
rect 13852 16406 13867 16478
rect 13913 16406 13928 16478
rect 13852 16354 13864 16406
rect 13916 16354 13928 16406
rect 13852 16282 13867 16354
rect 13913 16282 13928 16354
rect 13852 16230 13864 16282
rect 13916 16230 13928 16282
rect 13852 16158 13867 16230
rect 13913 16158 13928 16230
rect 13852 16106 13864 16158
rect 13916 16106 13928 16158
rect 13852 16034 13867 16106
rect 13913 16034 13928 16106
rect 13852 15982 13864 16034
rect 13916 15982 13928 16034
rect 13852 15910 13867 15982
rect 13913 15910 13928 15982
rect 13852 15858 13864 15910
rect 13916 15858 13928 15910
rect 13852 15786 13867 15858
rect 13913 15786 13928 15858
rect 13852 15734 13864 15786
rect 13916 15734 13928 15786
rect 13852 15662 13867 15734
rect 13913 15662 13928 15734
rect 13852 15610 13864 15662
rect 13916 15610 13928 15662
rect 13852 15538 13867 15610
rect 13913 15538 13928 15610
rect 13852 15486 13864 15538
rect 13916 15486 13928 15538
rect 13852 15474 13867 15486
rect 13689 14996 13704 15008
rect 13628 14944 13640 14996
rect 13692 14944 13704 14996
rect 13628 14872 13643 14944
rect 13689 14872 13704 14944
rect 13628 14820 13640 14872
rect 13692 14820 13704 14872
rect 13628 14748 13643 14820
rect 13689 14748 13704 14820
rect 13628 14696 13640 14748
rect 13692 14696 13704 14748
rect 13628 14624 13643 14696
rect 13689 14624 13704 14696
rect 13628 14572 13640 14624
rect 13692 14572 13704 14624
rect 13628 14500 13643 14572
rect 13689 14500 13704 14572
rect 13628 14448 13640 14500
rect 13692 14448 13704 14500
rect 13628 14376 13643 14448
rect 13689 14376 13704 14448
rect 13628 14324 13640 14376
rect 13692 14324 13704 14376
rect 13628 14252 13643 14324
rect 13689 14252 13704 14324
rect 13628 14200 13640 14252
rect 13692 14200 13704 14252
rect 13628 14128 13643 14200
rect 13689 14128 13704 14200
rect 13628 14076 13640 14128
rect 13692 14076 13704 14128
rect 13628 14004 13643 14076
rect 13689 14004 13704 14076
rect 13628 13952 13640 14004
rect 13692 13952 13704 14004
rect 13628 13880 13643 13952
rect 13689 13880 13704 13952
rect 13628 13828 13640 13880
rect 13692 13828 13704 13880
rect 13628 13756 13643 13828
rect 13689 13756 13704 13828
rect 13628 13704 13640 13756
rect 13692 13704 13704 13756
rect 13628 13632 13643 13704
rect 13689 13632 13704 13704
rect 13628 13580 13640 13632
rect 13692 13580 13704 13632
rect 13628 13508 13643 13580
rect 13689 13508 13704 13580
rect 13628 13456 13640 13508
rect 13692 13456 13704 13508
rect 13628 13384 13643 13456
rect 13689 13384 13704 13456
rect 13628 13332 13640 13384
rect 13692 13332 13704 13384
rect 13628 13260 13643 13332
rect 13689 13260 13704 13332
rect 13628 13208 13640 13260
rect 13692 13208 13704 13260
rect 13628 13136 13643 13208
rect 13689 13136 13704 13208
rect 13628 13084 13640 13136
rect 13692 13084 13704 13136
rect 13628 13012 13643 13084
rect 13689 13012 13704 13084
rect 13628 12960 13640 13012
rect 13692 12960 13704 13012
rect 13628 12888 13643 12960
rect 13689 12888 13704 12960
rect 13628 12836 13640 12888
rect 13692 12836 13704 12888
rect 13628 12824 13643 12836
rect 12985 12458 13147 12469
rect 12985 12412 12996 12458
rect 13136 12412 13147 12458
rect 12985 12401 13147 12412
rect 13278 12427 13346 12438
rect 12655 12263 12911 12274
rect 12655 12217 12666 12263
rect 12900 12217 12911 12263
rect 12655 12206 12911 12217
rect 13082 11958 13128 12401
rect 13278 12381 13289 12427
rect 13335 12381 13346 12427
rect 12299 11947 13147 11958
rect 12299 11901 12996 11947
rect 13136 11901 13147 11947
rect 13278 11923 13346 12381
rect 12299 11890 13147 11901
rect 13196 11911 13346 11923
rect 11388 11758 11464 11770
rect 11388 11706 11400 11758
rect 11452 11706 11464 11758
rect 11388 11634 11403 11706
rect 11449 11634 11464 11706
rect 11388 11582 11400 11634
rect 11452 11582 11464 11634
rect 11388 11510 11403 11582
rect 11449 11510 11464 11582
rect 11388 11458 11400 11510
rect 11452 11458 11464 11510
rect 11388 11446 11403 11458
rect 11179 10940 11225 10997
rect 11179 10837 11225 10894
rect 11179 10734 11225 10791
rect 11179 10631 11225 10688
rect 11179 10528 11225 10585
rect 11179 10425 11225 10482
rect 11179 10322 11225 10379
rect 11179 10219 11225 10276
rect 11179 10116 11225 10173
rect 11001 10070 11036 10109
rect 10921 10013 11036 10070
rect 10921 9967 10955 10013
rect 11001 9967 11036 10013
rect 10921 9863 11036 9967
rect 11179 10013 11225 10070
rect 11179 9954 11225 9967
rect 11449 11446 11464 11458
rect 11627 11757 11673 11770
rect 11403 10940 11449 10997
rect 11403 10837 11449 10894
rect 11403 10734 11449 10791
rect 11403 10631 11449 10688
rect 11403 10528 11449 10585
rect 11403 10425 11449 10482
rect 11403 10322 11449 10379
rect 11403 10219 11449 10276
rect 11403 10116 11449 10173
rect 11836 11758 11912 11770
rect 11836 11706 11848 11758
rect 11900 11706 11912 11758
rect 11836 11634 11851 11706
rect 11897 11634 11912 11706
rect 11836 11582 11848 11634
rect 11900 11582 11912 11634
rect 11836 11510 11851 11582
rect 11897 11510 11912 11582
rect 11836 11458 11848 11510
rect 11900 11458 11912 11510
rect 11836 11446 11851 11458
rect 11627 10940 11673 10997
rect 11627 10837 11673 10894
rect 11627 10734 11673 10791
rect 11627 10631 11673 10688
rect 11627 10528 11673 10585
rect 11627 10425 11673 10482
rect 11627 10322 11673 10379
rect 11627 10219 11673 10276
rect 11627 10116 11673 10173
rect 11403 10013 11449 10070
rect 11403 9954 11449 9967
rect 11593 10070 11627 10109
rect 11897 11446 11912 11458
rect 12075 11757 12121 11770
rect 11851 10940 11897 10997
rect 11851 10837 11897 10894
rect 11851 10734 11897 10791
rect 11851 10631 11897 10688
rect 11851 10528 11897 10585
rect 11851 10425 11897 10482
rect 11851 10322 11897 10379
rect 11851 10219 11897 10276
rect 11851 10116 11897 10173
rect 11673 10070 11708 10109
rect 11593 10013 11708 10070
rect 11593 9967 11627 10013
rect 11673 9967 11708 10013
rect 11593 9863 11708 9967
rect 12075 10940 12121 10997
rect 12075 10837 12121 10894
rect 12075 10734 12121 10791
rect 12075 10631 12121 10688
rect 12075 10528 12121 10585
rect 12075 10425 12121 10482
rect 12075 10322 12121 10379
rect 12075 10219 12121 10276
rect 12075 10116 12121 10173
rect 11851 10013 11897 10070
rect 11851 9954 11897 9967
rect 12041 10070 12075 10109
rect 12299 11757 12345 11890
rect 13196 11859 13208 11911
rect 13260 11905 13346 11911
rect 13260 11859 13289 11905
rect 13335 11859 13346 11905
rect 13196 11840 13346 11859
rect 13419 11958 13465 12598
rect 13689 12824 13704 12836
rect 13643 12585 13689 12598
rect 13913 15474 13928 15486
rect 14091 16572 14137 16585
rect 14076 14996 14091 15008
rect 14300 16572 14376 16602
rect 14972 16654 15048 16682
rect 14972 16602 14984 16654
rect 15036 16602 15048 16654
rect 14300 16530 14315 16572
rect 14361 16530 14376 16572
rect 14300 16478 14312 16530
rect 14364 16478 14376 16530
rect 14300 16406 14315 16478
rect 14361 16406 14376 16478
rect 14300 16354 14312 16406
rect 14364 16354 14376 16406
rect 14300 16282 14315 16354
rect 14361 16282 14376 16354
rect 14300 16230 14312 16282
rect 14364 16230 14376 16282
rect 14300 16158 14315 16230
rect 14361 16158 14376 16230
rect 14300 16106 14312 16158
rect 14364 16106 14376 16158
rect 14300 16034 14315 16106
rect 14361 16034 14376 16106
rect 14300 15982 14312 16034
rect 14364 15982 14376 16034
rect 14300 15910 14315 15982
rect 14361 15910 14376 15982
rect 14300 15858 14312 15910
rect 14364 15858 14376 15910
rect 14300 15786 14315 15858
rect 14361 15786 14376 15858
rect 14300 15734 14312 15786
rect 14364 15734 14376 15786
rect 14300 15662 14315 15734
rect 14361 15662 14376 15734
rect 14300 15610 14312 15662
rect 14364 15610 14376 15662
rect 14300 15538 14315 15610
rect 14361 15538 14376 15610
rect 14300 15486 14312 15538
rect 14364 15486 14376 15538
rect 14300 15474 14315 15486
rect 14137 14996 14152 15008
rect 14076 14944 14088 14996
rect 14140 14944 14152 14996
rect 14076 14872 14091 14944
rect 14137 14872 14152 14944
rect 14076 14820 14088 14872
rect 14140 14820 14152 14872
rect 14076 14748 14091 14820
rect 14137 14748 14152 14820
rect 14076 14696 14088 14748
rect 14140 14696 14152 14748
rect 14076 14624 14091 14696
rect 14137 14624 14152 14696
rect 14076 14572 14088 14624
rect 14140 14572 14152 14624
rect 14076 14500 14091 14572
rect 14137 14500 14152 14572
rect 14076 14448 14088 14500
rect 14140 14448 14152 14500
rect 14076 14376 14091 14448
rect 14137 14376 14152 14448
rect 14076 14324 14088 14376
rect 14140 14324 14152 14376
rect 14076 14252 14091 14324
rect 14137 14252 14152 14324
rect 14076 14200 14088 14252
rect 14140 14200 14152 14252
rect 14076 14128 14091 14200
rect 14137 14128 14152 14200
rect 14076 14076 14088 14128
rect 14140 14076 14152 14128
rect 14076 14004 14091 14076
rect 14137 14004 14152 14076
rect 14076 13952 14088 14004
rect 14140 13952 14152 14004
rect 14076 13880 14091 13952
rect 14137 13880 14152 13952
rect 14076 13828 14088 13880
rect 14140 13828 14152 13880
rect 14076 13756 14091 13828
rect 14137 13756 14152 13828
rect 14076 13704 14088 13756
rect 14140 13704 14152 13756
rect 14076 13632 14091 13704
rect 14137 13632 14152 13704
rect 14076 13580 14088 13632
rect 14140 13580 14152 13632
rect 14076 13508 14091 13580
rect 14137 13508 14152 13580
rect 14076 13456 14088 13508
rect 14140 13456 14152 13508
rect 14076 13384 14091 13456
rect 14137 13384 14152 13456
rect 14076 13332 14088 13384
rect 14140 13332 14152 13384
rect 14076 13260 14091 13332
rect 14137 13260 14152 13332
rect 14076 13208 14088 13260
rect 14140 13208 14152 13260
rect 14076 13136 14091 13208
rect 14137 13136 14152 13208
rect 14076 13084 14088 13136
rect 14140 13084 14152 13136
rect 14076 13012 14091 13084
rect 14137 13012 14152 13084
rect 14076 12960 14088 13012
rect 14140 12960 14152 13012
rect 14076 12888 14091 12960
rect 14137 12888 14152 12960
rect 14076 12836 14088 12888
rect 14140 12836 14152 12888
rect 14076 12824 14091 12836
rect 13867 12274 13913 12598
rect 14137 12824 14152 12836
rect 14091 12585 14137 12598
rect 14361 15474 14376 15486
rect 14539 16572 14585 16585
rect 14315 12585 14361 12598
rect 14763 16572 14809 16585
rect 14748 14996 14763 15008
rect 14972 16572 15048 16602
rect 15420 16654 15496 16682
rect 15420 16602 15432 16654
rect 15484 16602 15496 16654
rect 14972 16530 14987 16572
rect 15033 16530 15048 16572
rect 14972 16478 14984 16530
rect 15036 16478 15048 16530
rect 14972 16406 14987 16478
rect 15033 16406 15048 16478
rect 14972 16354 14984 16406
rect 15036 16354 15048 16406
rect 14972 16282 14987 16354
rect 15033 16282 15048 16354
rect 14972 16230 14984 16282
rect 15036 16230 15048 16282
rect 14972 16158 14987 16230
rect 15033 16158 15048 16230
rect 14972 16106 14984 16158
rect 15036 16106 15048 16158
rect 14972 16034 14987 16106
rect 15033 16034 15048 16106
rect 14972 15982 14984 16034
rect 15036 15982 15048 16034
rect 14972 15910 14987 15982
rect 15033 15910 15048 15982
rect 14972 15858 14984 15910
rect 15036 15858 15048 15910
rect 14972 15786 14987 15858
rect 15033 15786 15048 15858
rect 14972 15734 14984 15786
rect 15036 15734 15048 15786
rect 14972 15662 14987 15734
rect 15033 15662 15048 15734
rect 14972 15610 14984 15662
rect 15036 15610 15048 15662
rect 14972 15538 14987 15610
rect 15033 15538 15048 15610
rect 14972 15486 14984 15538
rect 15036 15486 15048 15538
rect 14972 15474 14987 15486
rect 14809 14996 14824 15008
rect 14748 14944 14760 14996
rect 14812 14944 14824 14996
rect 14748 14872 14763 14944
rect 14809 14872 14824 14944
rect 14748 14820 14760 14872
rect 14812 14820 14824 14872
rect 14748 14748 14763 14820
rect 14809 14748 14824 14820
rect 14748 14696 14760 14748
rect 14812 14696 14824 14748
rect 14748 14624 14763 14696
rect 14809 14624 14824 14696
rect 14748 14572 14760 14624
rect 14812 14572 14824 14624
rect 14748 14500 14763 14572
rect 14809 14500 14824 14572
rect 14748 14448 14760 14500
rect 14812 14448 14824 14500
rect 14748 14376 14763 14448
rect 14809 14376 14824 14448
rect 14748 14324 14760 14376
rect 14812 14324 14824 14376
rect 14748 14252 14763 14324
rect 14809 14252 14824 14324
rect 14748 14200 14760 14252
rect 14812 14200 14824 14252
rect 14748 14128 14763 14200
rect 14809 14128 14824 14200
rect 14748 14076 14760 14128
rect 14812 14076 14824 14128
rect 14748 14004 14763 14076
rect 14809 14004 14824 14076
rect 14748 13952 14760 14004
rect 14812 13952 14824 14004
rect 14748 13880 14763 13952
rect 14809 13880 14824 13952
rect 14748 13828 14760 13880
rect 14812 13828 14824 13880
rect 14748 13756 14763 13828
rect 14809 13756 14824 13828
rect 14748 13704 14760 13756
rect 14812 13704 14824 13756
rect 14748 13632 14763 13704
rect 14809 13632 14824 13704
rect 14748 13580 14760 13632
rect 14812 13580 14824 13632
rect 14748 13508 14763 13580
rect 14809 13508 14824 13580
rect 14748 13456 14760 13508
rect 14812 13456 14824 13508
rect 14748 13384 14763 13456
rect 14809 13384 14824 13456
rect 14748 13332 14760 13384
rect 14812 13332 14824 13384
rect 14748 13260 14763 13332
rect 14809 13260 14824 13332
rect 14748 13208 14760 13260
rect 14812 13208 14824 13260
rect 14748 13136 14763 13208
rect 14809 13136 14824 13208
rect 14748 13084 14760 13136
rect 14812 13084 14824 13136
rect 14748 13012 14763 13084
rect 14809 13012 14824 13084
rect 14748 12960 14760 13012
rect 14812 12960 14824 13012
rect 14748 12888 14763 12960
rect 14809 12888 14824 12960
rect 14748 12836 14760 12888
rect 14812 12836 14824 12888
rect 14748 12824 14763 12836
rect 14105 12458 14267 12469
rect 14105 12412 14116 12458
rect 14256 12412 14267 12458
rect 14105 12401 14267 12412
rect 14398 12427 14466 12438
rect 13775 12263 14031 12274
rect 13775 12217 13786 12263
rect 14020 12217 14031 12263
rect 13775 12206 14031 12217
rect 14202 11958 14248 12401
rect 14398 12381 14409 12427
rect 14455 12381 14466 12427
rect 13419 11947 14267 11958
rect 13419 11901 14116 11947
rect 14256 11901 14267 11947
rect 14398 11923 14466 12381
rect 13419 11890 14267 11901
rect 14316 11911 14466 11923
rect 12508 11758 12584 11770
rect 12508 11706 12520 11758
rect 12572 11706 12584 11758
rect 12508 11634 12523 11706
rect 12569 11634 12584 11706
rect 12508 11582 12520 11634
rect 12572 11582 12584 11634
rect 12508 11510 12523 11582
rect 12569 11510 12584 11582
rect 12508 11458 12520 11510
rect 12572 11458 12584 11510
rect 12508 11446 12523 11458
rect 12299 10940 12345 10997
rect 12299 10837 12345 10894
rect 12299 10734 12345 10791
rect 12299 10631 12345 10688
rect 12299 10528 12345 10585
rect 12299 10425 12345 10482
rect 12299 10322 12345 10379
rect 12299 10219 12345 10276
rect 12299 10116 12345 10173
rect 12121 10070 12156 10109
rect 12041 10013 12156 10070
rect 12041 9967 12075 10013
rect 12121 9967 12156 10013
rect 12041 9863 12156 9967
rect 12299 10013 12345 10070
rect 12299 9954 12345 9967
rect 12569 11446 12584 11458
rect 12747 11757 12793 11770
rect 12523 10940 12569 10997
rect 12523 10837 12569 10894
rect 12523 10734 12569 10791
rect 12523 10631 12569 10688
rect 12523 10528 12569 10585
rect 12523 10425 12569 10482
rect 12523 10322 12569 10379
rect 12523 10219 12569 10276
rect 12523 10116 12569 10173
rect 12956 11758 13032 11770
rect 12956 11706 12968 11758
rect 13020 11706 13032 11758
rect 12956 11634 12971 11706
rect 13017 11634 13032 11706
rect 12956 11582 12968 11634
rect 13020 11582 13032 11634
rect 12956 11510 12971 11582
rect 13017 11510 13032 11582
rect 12956 11458 12968 11510
rect 13020 11458 13032 11510
rect 12956 11446 12971 11458
rect 12747 10940 12793 10997
rect 12747 10837 12793 10894
rect 12747 10734 12793 10791
rect 12747 10631 12793 10688
rect 12747 10528 12793 10585
rect 12747 10425 12793 10482
rect 12747 10322 12793 10379
rect 12747 10219 12793 10276
rect 12747 10116 12793 10173
rect 12523 10013 12569 10070
rect 12523 9954 12569 9967
rect 12713 10070 12747 10109
rect 13017 11446 13032 11458
rect 13195 11757 13241 11770
rect 12971 10940 13017 10997
rect 12971 10837 13017 10894
rect 12971 10734 13017 10791
rect 12971 10631 13017 10688
rect 12971 10528 13017 10585
rect 12971 10425 13017 10482
rect 12971 10322 13017 10379
rect 12971 10219 13017 10276
rect 12971 10116 13017 10173
rect 12793 10070 12828 10109
rect 12713 10013 12828 10070
rect 12713 9967 12747 10013
rect 12793 9967 12828 10013
rect 12713 9863 12828 9967
rect 13195 10940 13241 10997
rect 13195 10837 13241 10894
rect 13195 10734 13241 10791
rect 13195 10631 13241 10688
rect 13195 10528 13241 10585
rect 13195 10425 13241 10482
rect 13195 10322 13241 10379
rect 13195 10219 13241 10276
rect 13195 10116 13241 10173
rect 12971 10013 13017 10070
rect 12971 9954 13017 9967
rect 13161 10070 13195 10109
rect 13419 11757 13465 11890
rect 14316 11859 14328 11911
rect 14380 11905 14466 11911
rect 14380 11859 14409 11905
rect 14455 11859 14466 11905
rect 14316 11840 14466 11859
rect 14539 11958 14585 12598
rect 14809 12824 14824 12836
rect 14763 12585 14809 12598
rect 15033 15474 15048 15486
rect 15211 16572 15257 16585
rect 15196 14996 15211 15008
rect 15420 16572 15496 16602
rect 16092 16654 16168 16682
rect 16092 16602 16104 16654
rect 16156 16602 16168 16654
rect 15420 16530 15435 16572
rect 15481 16530 15496 16572
rect 15420 16478 15432 16530
rect 15484 16478 15496 16530
rect 15420 16406 15435 16478
rect 15481 16406 15496 16478
rect 15420 16354 15432 16406
rect 15484 16354 15496 16406
rect 15420 16282 15435 16354
rect 15481 16282 15496 16354
rect 15420 16230 15432 16282
rect 15484 16230 15496 16282
rect 15420 16158 15435 16230
rect 15481 16158 15496 16230
rect 15420 16106 15432 16158
rect 15484 16106 15496 16158
rect 15420 16034 15435 16106
rect 15481 16034 15496 16106
rect 15420 15982 15432 16034
rect 15484 15982 15496 16034
rect 15420 15910 15435 15982
rect 15481 15910 15496 15982
rect 15420 15858 15432 15910
rect 15484 15858 15496 15910
rect 15420 15786 15435 15858
rect 15481 15786 15496 15858
rect 15420 15734 15432 15786
rect 15484 15734 15496 15786
rect 15420 15662 15435 15734
rect 15481 15662 15496 15734
rect 15420 15610 15432 15662
rect 15484 15610 15496 15662
rect 15420 15538 15435 15610
rect 15481 15538 15496 15610
rect 15420 15486 15432 15538
rect 15484 15486 15496 15538
rect 15420 15474 15435 15486
rect 15257 14996 15272 15008
rect 15196 14944 15208 14996
rect 15260 14944 15272 14996
rect 15196 14872 15211 14944
rect 15257 14872 15272 14944
rect 15196 14820 15208 14872
rect 15260 14820 15272 14872
rect 15196 14748 15211 14820
rect 15257 14748 15272 14820
rect 15196 14696 15208 14748
rect 15260 14696 15272 14748
rect 15196 14624 15211 14696
rect 15257 14624 15272 14696
rect 15196 14572 15208 14624
rect 15260 14572 15272 14624
rect 15196 14500 15211 14572
rect 15257 14500 15272 14572
rect 15196 14448 15208 14500
rect 15260 14448 15272 14500
rect 15196 14376 15211 14448
rect 15257 14376 15272 14448
rect 15196 14324 15208 14376
rect 15260 14324 15272 14376
rect 15196 14252 15211 14324
rect 15257 14252 15272 14324
rect 15196 14200 15208 14252
rect 15260 14200 15272 14252
rect 15196 14128 15211 14200
rect 15257 14128 15272 14200
rect 15196 14076 15208 14128
rect 15260 14076 15272 14128
rect 15196 14004 15211 14076
rect 15257 14004 15272 14076
rect 15196 13952 15208 14004
rect 15260 13952 15272 14004
rect 15196 13880 15211 13952
rect 15257 13880 15272 13952
rect 15196 13828 15208 13880
rect 15260 13828 15272 13880
rect 15196 13756 15211 13828
rect 15257 13756 15272 13828
rect 15196 13704 15208 13756
rect 15260 13704 15272 13756
rect 15196 13632 15211 13704
rect 15257 13632 15272 13704
rect 15196 13580 15208 13632
rect 15260 13580 15272 13632
rect 15196 13508 15211 13580
rect 15257 13508 15272 13580
rect 15196 13456 15208 13508
rect 15260 13456 15272 13508
rect 15196 13384 15211 13456
rect 15257 13384 15272 13456
rect 15196 13332 15208 13384
rect 15260 13332 15272 13384
rect 15196 13260 15211 13332
rect 15257 13260 15272 13332
rect 15196 13208 15208 13260
rect 15260 13208 15272 13260
rect 15196 13136 15211 13208
rect 15257 13136 15272 13208
rect 15196 13084 15208 13136
rect 15260 13084 15272 13136
rect 15196 13012 15211 13084
rect 15257 13012 15272 13084
rect 15196 12960 15208 13012
rect 15260 12960 15272 13012
rect 15196 12888 15211 12960
rect 15257 12888 15272 12960
rect 15196 12836 15208 12888
rect 15260 12836 15272 12888
rect 15196 12824 15211 12836
rect 14987 12274 15033 12598
rect 15257 12824 15272 12836
rect 15211 12585 15257 12598
rect 15481 15474 15496 15486
rect 15659 16572 15705 16585
rect 15435 12585 15481 12598
rect 15883 16572 15929 16585
rect 15868 14996 15883 15008
rect 16092 16572 16168 16602
rect 16540 16654 16616 16682
rect 16540 16602 16552 16654
rect 16604 16602 16616 16654
rect 16092 16530 16107 16572
rect 16153 16530 16168 16572
rect 16092 16478 16104 16530
rect 16156 16478 16168 16530
rect 16092 16406 16107 16478
rect 16153 16406 16168 16478
rect 16092 16354 16104 16406
rect 16156 16354 16168 16406
rect 16092 16282 16107 16354
rect 16153 16282 16168 16354
rect 16092 16230 16104 16282
rect 16156 16230 16168 16282
rect 16092 16158 16107 16230
rect 16153 16158 16168 16230
rect 16092 16106 16104 16158
rect 16156 16106 16168 16158
rect 16092 16034 16107 16106
rect 16153 16034 16168 16106
rect 16092 15982 16104 16034
rect 16156 15982 16168 16034
rect 16092 15910 16107 15982
rect 16153 15910 16168 15982
rect 16092 15858 16104 15910
rect 16156 15858 16168 15910
rect 16092 15786 16107 15858
rect 16153 15786 16168 15858
rect 16092 15734 16104 15786
rect 16156 15734 16168 15786
rect 16092 15662 16107 15734
rect 16153 15662 16168 15734
rect 16092 15610 16104 15662
rect 16156 15610 16168 15662
rect 16092 15538 16107 15610
rect 16153 15538 16168 15610
rect 16092 15486 16104 15538
rect 16156 15486 16168 15538
rect 16092 15474 16107 15486
rect 15929 14996 15944 15008
rect 15868 14944 15880 14996
rect 15932 14944 15944 14996
rect 15868 14872 15883 14944
rect 15929 14872 15944 14944
rect 15868 14820 15880 14872
rect 15932 14820 15944 14872
rect 15868 14748 15883 14820
rect 15929 14748 15944 14820
rect 15868 14696 15880 14748
rect 15932 14696 15944 14748
rect 15868 14624 15883 14696
rect 15929 14624 15944 14696
rect 15868 14572 15880 14624
rect 15932 14572 15944 14624
rect 15868 14500 15883 14572
rect 15929 14500 15944 14572
rect 15868 14448 15880 14500
rect 15932 14448 15944 14500
rect 15868 14376 15883 14448
rect 15929 14376 15944 14448
rect 15868 14324 15880 14376
rect 15932 14324 15944 14376
rect 15868 14252 15883 14324
rect 15929 14252 15944 14324
rect 15868 14200 15880 14252
rect 15932 14200 15944 14252
rect 15868 14128 15883 14200
rect 15929 14128 15944 14200
rect 15868 14076 15880 14128
rect 15932 14076 15944 14128
rect 15868 14004 15883 14076
rect 15929 14004 15944 14076
rect 15868 13952 15880 14004
rect 15932 13952 15944 14004
rect 15868 13880 15883 13952
rect 15929 13880 15944 13952
rect 15868 13828 15880 13880
rect 15932 13828 15944 13880
rect 15868 13756 15883 13828
rect 15929 13756 15944 13828
rect 15868 13704 15880 13756
rect 15932 13704 15944 13756
rect 15868 13632 15883 13704
rect 15929 13632 15944 13704
rect 15868 13580 15880 13632
rect 15932 13580 15944 13632
rect 15868 13508 15883 13580
rect 15929 13508 15944 13580
rect 15868 13456 15880 13508
rect 15932 13456 15944 13508
rect 15868 13384 15883 13456
rect 15929 13384 15944 13456
rect 15868 13332 15880 13384
rect 15932 13332 15944 13384
rect 15868 13260 15883 13332
rect 15929 13260 15944 13332
rect 15868 13208 15880 13260
rect 15932 13208 15944 13260
rect 15868 13136 15883 13208
rect 15929 13136 15944 13208
rect 15868 13084 15880 13136
rect 15932 13084 15944 13136
rect 15868 13012 15883 13084
rect 15929 13012 15944 13084
rect 15868 12960 15880 13012
rect 15932 12960 15944 13012
rect 15868 12888 15883 12960
rect 15929 12888 15944 12960
rect 15868 12836 15880 12888
rect 15932 12836 15944 12888
rect 15868 12824 15883 12836
rect 15225 12458 15387 12469
rect 15225 12412 15236 12458
rect 15376 12412 15387 12458
rect 15225 12401 15387 12412
rect 15518 12427 15586 12438
rect 14895 12263 15151 12274
rect 14895 12217 14906 12263
rect 15140 12217 15151 12263
rect 14895 12206 15151 12217
rect 15322 11958 15368 12401
rect 15518 12381 15529 12427
rect 15575 12381 15586 12427
rect 14539 11947 15387 11958
rect 14539 11901 15236 11947
rect 15376 11901 15387 11947
rect 15518 11923 15586 12381
rect 14539 11890 15387 11901
rect 15436 11911 15586 11923
rect 13628 11758 13704 11770
rect 13628 11706 13640 11758
rect 13692 11706 13704 11758
rect 13628 11634 13643 11706
rect 13689 11634 13704 11706
rect 13628 11582 13640 11634
rect 13692 11582 13704 11634
rect 13628 11510 13643 11582
rect 13689 11510 13704 11582
rect 13628 11458 13640 11510
rect 13692 11458 13704 11510
rect 13628 11446 13643 11458
rect 13419 10940 13465 10997
rect 13419 10837 13465 10894
rect 13419 10734 13465 10791
rect 13419 10631 13465 10688
rect 13419 10528 13465 10585
rect 13419 10425 13465 10482
rect 13419 10322 13465 10379
rect 13419 10219 13465 10276
rect 13419 10116 13465 10173
rect 13241 10070 13276 10109
rect 13161 10013 13276 10070
rect 13161 9967 13195 10013
rect 13241 9967 13276 10013
rect 13161 9863 13276 9967
rect 13419 10013 13465 10070
rect 13419 9954 13465 9967
rect 13689 11446 13704 11458
rect 13867 11757 13913 11770
rect 13643 10940 13689 10997
rect 13643 10837 13689 10894
rect 13643 10734 13689 10791
rect 13643 10631 13689 10688
rect 13643 10528 13689 10585
rect 13643 10425 13689 10482
rect 13643 10322 13689 10379
rect 13643 10219 13689 10276
rect 13643 10116 13689 10173
rect 14076 11758 14152 11770
rect 14076 11706 14088 11758
rect 14140 11706 14152 11758
rect 14076 11634 14091 11706
rect 14137 11634 14152 11706
rect 14076 11582 14088 11634
rect 14140 11582 14152 11634
rect 14076 11510 14091 11582
rect 14137 11510 14152 11582
rect 14076 11458 14088 11510
rect 14140 11458 14152 11510
rect 14076 11446 14091 11458
rect 13867 10940 13913 10997
rect 13867 10837 13913 10894
rect 13867 10734 13913 10791
rect 13867 10631 13913 10688
rect 13867 10528 13913 10585
rect 13867 10425 13913 10482
rect 13867 10322 13913 10379
rect 13867 10219 13913 10276
rect 13867 10116 13913 10173
rect 13643 10013 13689 10070
rect 13643 9954 13689 9967
rect 13833 10070 13867 10109
rect 14137 11446 14152 11458
rect 14315 11757 14361 11770
rect 14091 10940 14137 10997
rect 14091 10837 14137 10894
rect 14091 10734 14137 10791
rect 14091 10631 14137 10688
rect 14091 10528 14137 10585
rect 14091 10425 14137 10482
rect 14091 10322 14137 10379
rect 14091 10219 14137 10276
rect 14091 10116 14137 10173
rect 13913 10070 13948 10109
rect 13833 10013 13948 10070
rect 13833 9967 13867 10013
rect 13913 9967 13948 10013
rect 13833 9863 13948 9967
rect 14315 10940 14361 10997
rect 14315 10837 14361 10894
rect 14315 10734 14361 10791
rect 14315 10631 14361 10688
rect 14315 10528 14361 10585
rect 14315 10425 14361 10482
rect 14315 10322 14361 10379
rect 14315 10219 14361 10276
rect 14315 10116 14361 10173
rect 14091 10013 14137 10070
rect 14091 9954 14137 9967
rect 14281 10070 14315 10109
rect 14539 11757 14585 11890
rect 15436 11859 15448 11911
rect 15500 11905 15586 11911
rect 15500 11859 15529 11905
rect 15575 11859 15586 11905
rect 15436 11840 15586 11859
rect 15659 11958 15705 12598
rect 15929 12824 15944 12836
rect 15883 12585 15929 12598
rect 16153 15474 16168 15486
rect 16331 16572 16377 16585
rect 16316 14996 16331 15008
rect 16540 16572 16616 16602
rect 17212 16654 17288 16682
rect 17212 16602 17224 16654
rect 17276 16602 17288 16654
rect 16540 16530 16555 16572
rect 16601 16530 16616 16572
rect 16540 16478 16552 16530
rect 16604 16478 16616 16530
rect 16540 16406 16555 16478
rect 16601 16406 16616 16478
rect 16540 16354 16552 16406
rect 16604 16354 16616 16406
rect 16540 16282 16555 16354
rect 16601 16282 16616 16354
rect 16540 16230 16552 16282
rect 16604 16230 16616 16282
rect 16540 16158 16555 16230
rect 16601 16158 16616 16230
rect 16540 16106 16552 16158
rect 16604 16106 16616 16158
rect 16540 16034 16555 16106
rect 16601 16034 16616 16106
rect 16540 15982 16552 16034
rect 16604 15982 16616 16034
rect 16540 15910 16555 15982
rect 16601 15910 16616 15982
rect 16540 15858 16552 15910
rect 16604 15858 16616 15910
rect 16540 15786 16555 15858
rect 16601 15786 16616 15858
rect 16540 15734 16552 15786
rect 16604 15734 16616 15786
rect 16540 15662 16555 15734
rect 16601 15662 16616 15734
rect 16540 15610 16552 15662
rect 16604 15610 16616 15662
rect 16540 15538 16555 15610
rect 16601 15538 16616 15610
rect 16540 15486 16552 15538
rect 16604 15486 16616 15538
rect 16540 15474 16555 15486
rect 16377 14996 16392 15008
rect 16316 14944 16328 14996
rect 16380 14944 16392 14996
rect 16316 14872 16331 14944
rect 16377 14872 16392 14944
rect 16316 14820 16328 14872
rect 16380 14820 16392 14872
rect 16316 14748 16331 14820
rect 16377 14748 16392 14820
rect 16316 14696 16328 14748
rect 16380 14696 16392 14748
rect 16316 14624 16331 14696
rect 16377 14624 16392 14696
rect 16316 14572 16328 14624
rect 16380 14572 16392 14624
rect 16316 14500 16331 14572
rect 16377 14500 16392 14572
rect 16316 14448 16328 14500
rect 16380 14448 16392 14500
rect 16316 14376 16331 14448
rect 16377 14376 16392 14448
rect 16316 14324 16328 14376
rect 16380 14324 16392 14376
rect 16316 14252 16331 14324
rect 16377 14252 16392 14324
rect 16316 14200 16328 14252
rect 16380 14200 16392 14252
rect 16316 14128 16331 14200
rect 16377 14128 16392 14200
rect 16316 14076 16328 14128
rect 16380 14076 16392 14128
rect 16316 14004 16331 14076
rect 16377 14004 16392 14076
rect 16316 13952 16328 14004
rect 16380 13952 16392 14004
rect 16316 13880 16331 13952
rect 16377 13880 16392 13952
rect 16316 13828 16328 13880
rect 16380 13828 16392 13880
rect 16316 13756 16331 13828
rect 16377 13756 16392 13828
rect 16316 13704 16328 13756
rect 16380 13704 16392 13756
rect 16316 13632 16331 13704
rect 16377 13632 16392 13704
rect 16316 13580 16328 13632
rect 16380 13580 16392 13632
rect 16316 13508 16331 13580
rect 16377 13508 16392 13580
rect 16316 13456 16328 13508
rect 16380 13456 16392 13508
rect 16316 13384 16331 13456
rect 16377 13384 16392 13456
rect 16316 13332 16328 13384
rect 16380 13332 16392 13384
rect 16316 13260 16331 13332
rect 16377 13260 16392 13332
rect 16316 13208 16328 13260
rect 16380 13208 16392 13260
rect 16316 13136 16331 13208
rect 16377 13136 16392 13208
rect 16316 13084 16328 13136
rect 16380 13084 16392 13136
rect 16316 13012 16331 13084
rect 16377 13012 16392 13084
rect 16316 12960 16328 13012
rect 16380 12960 16392 13012
rect 16316 12888 16331 12960
rect 16377 12888 16392 12960
rect 16316 12836 16328 12888
rect 16380 12836 16392 12888
rect 16316 12824 16331 12836
rect 16107 12274 16153 12598
rect 16377 12824 16392 12836
rect 16331 12585 16377 12598
rect 16601 15474 16616 15486
rect 16779 16572 16825 16585
rect 16555 12585 16601 12598
rect 17003 16572 17049 16585
rect 16988 14996 17003 15008
rect 17212 16572 17288 16602
rect 17660 16654 17736 16682
rect 17660 16602 17672 16654
rect 17724 16602 17736 16654
rect 17212 16530 17227 16572
rect 17273 16530 17288 16572
rect 17212 16478 17224 16530
rect 17276 16478 17288 16530
rect 17212 16406 17227 16478
rect 17273 16406 17288 16478
rect 17212 16354 17224 16406
rect 17276 16354 17288 16406
rect 17212 16282 17227 16354
rect 17273 16282 17288 16354
rect 17212 16230 17224 16282
rect 17276 16230 17288 16282
rect 17212 16158 17227 16230
rect 17273 16158 17288 16230
rect 17212 16106 17224 16158
rect 17276 16106 17288 16158
rect 17212 16034 17227 16106
rect 17273 16034 17288 16106
rect 17212 15982 17224 16034
rect 17276 15982 17288 16034
rect 17212 15910 17227 15982
rect 17273 15910 17288 15982
rect 17212 15858 17224 15910
rect 17276 15858 17288 15910
rect 17212 15786 17227 15858
rect 17273 15786 17288 15858
rect 17212 15734 17224 15786
rect 17276 15734 17288 15786
rect 17212 15662 17227 15734
rect 17273 15662 17288 15734
rect 17212 15610 17224 15662
rect 17276 15610 17288 15662
rect 17212 15538 17227 15610
rect 17273 15538 17288 15610
rect 17212 15486 17224 15538
rect 17276 15486 17288 15538
rect 17212 15474 17227 15486
rect 17049 14996 17064 15008
rect 16988 14944 17000 14996
rect 17052 14944 17064 14996
rect 16988 14872 17003 14944
rect 17049 14872 17064 14944
rect 16988 14820 17000 14872
rect 17052 14820 17064 14872
rect 16988 14748 17003 14820
rect 17049 14748 17064 14820
rect 16988 14696 17000 14748
rect 17052 14696 17064 14748
rect 16988 14624 17003 14696
rect 17049 14624 17064 14696
rect 16988 14572 17000 14624
rect 17052 14572 17064 14624
rect 16988 14500 17003 14572
rect 17049 14500 17064 14572
rect 16988 14448 17000 14500
rect 17052 14448 17064 14500
rect 16988 14376 17003 14448
rect 17049 14376 17064 14448
rect 16988 14324 17000 14376
rect 17052 14324 17064 14376
rect 16988 14252 17003 14324
rect 17049 14252 17064 14324
rect 16988 14200 17000 14252
rect 17052 14200 17064 14252
rect 16988 14128 17003 14200
rect 17049 14128 17064 14200
rect 16988 14076 17000 14128
rect 17052 14076 17064 14128
rect 16988 14004 17003 14076
rect 17049 14004 17064 14076
rect 16988 13952 17000 14004
rect 17052 13952 17064 14004
rect 16988 13880 17003 13952
rect 17049 13880 17064 13952
rect 16988 13828 17000 13880
rect 17052 13828 17064 13880
rect 16988 13756 17003 13828
rect 17049 13756 17064 13828
rect 16988 13704 17000 13756
rect 17052 13704 17064 13756
rect 16988 13632 17003 13704
rect 17049 13632 17064 13704
rect 16988 13580 17000 13632
rect 17052 13580 17064 13632
rect 16988 13508 17003 13580
rect 17049 13508 17064 13580
rect 16988 13456 17000 13508
rect 17052 13456 17064 13508
rect 16988 13384 17003 13456
rect 17049 13384 17064 13456
rect 16988 13332 17000 13384
rect 17052 13332 17064 13384
rect 16988 13260 17003 13332
rect 17049 13260 17064 13332
rect 16988 13208 17000 13260
rect 17052 13208 17064 13260
rect 16988 13136 17003 13208
rect 17049 13136 17064 13208
rect 16988 13084 17000 13136
rect 17052 13084 17064 13136
rect 16988 13012 17003 13084
rect 17049 13012 17064 13084
rect 16988 12960 17000 13012
rect 17052 12960 17064 13012
rect 16988 12888 17003 12960
rect 17049 12888 17064 12960
rect 16988 12836 17000 12888
rect 17052 12836 17064 12888
rect 16988 12824 17003 12836
rect 16345 12458 16507 12469
rect 16345 12412 16356 12458
rect 16496 12412 16507 12458
rect 16345 12401 16507 12412
rect 16638 12427 16706 12438
rect 16015 12263 16271 12274
rect 16015 12217 16026 12263
rect 16260 12217 16271 12263
rect 16015 12206 16271 12217
rect 16442 11958 16488 12401
rect 16638 12381 16649 12427
rect 16695 12381 16706 12427
rect 15659 11947 16507 11958
rect 15659 11901 16356 11947
rect 16496 11901 16507 11947
rect 16638 11923 16706 12381
rect 15659 11890 16507 11901
rect 16556 11911 16706 11923
rect 14748 11758 14824 11770
rect 14748 11706 14760 11758
rect 14812 11706 14824 11758
rect 14748 11634 14763 11706
rect 14809 11634 14824 11706
rect 14748 11582 14760 11634
rect 14812 11582 14824 11634
rect 14748 11510 14763 11582
rect 14809 11510 14824 11582
rect 14748 11458 14760 11510
rect 14812 11458 14824 11510
rect 14748 11446 14763 11458
rect 14539 10940 14585 10997
rect 14539 10837 14585 10894
rect 14539 10734 14585 10791
rect 14539 10631 14585 10688
rect 14539 10528 14585 10585
rect 14539 10425 14585 10482
rect 14539 10322 14585 10379
rect 14539 10219 14585 10276
rect 14539 10116 14585 10173
rect 14361 10070 14396 10109
rect 14281 10013 14396 10070
rect 14281 9967 14315 10013
rect 14361 9967 14396 10013
rect 14281 9863 14396 9967
rect 14539 10013 14585 10070
rect 14539 9954 14585 9967
rect 14809 11446 14824 11458
rect 14987 11757 15033 11770
rect 14763 10940 14809 10997
rect 14763 10837 14809 10894
rect 14763 10734 14809 10791
rect 14763 10631 14809 10688
rect 14763 10528 14809 10585
rect 14763 10425 14809 10482
rect 14763 10322 14809 10379
rect 14763 10219 14809 10276
rect 14763 10116 14809 10173
rect 15196 11758 15272 11770
rect 15196 11706 15208 11758
rect 15260 11706 15272 11758
rect 15196 11634 15211 11706
rect 15257 11634 15272 11706
rect 15196 11582 15208 11634
rect 15260 11582 15272 11634
rect 15196 11510 15211 11582
rect 15257 11510 15272 11582
rect 15196 11458 15208 11510
rect 15260 11458 15272 11510
rect 15196 11446 15211 11458
rect 14987 10940 15033 10997
rect 14987 10837 15033 10894
rect 14987 10734 15033 10791
rect 14987 10631 15033 10688
rect 14987 10528 15033 10585
rect 14987 10425 15033 10482
rect 14987 10322 15033 10379
rect 14987 10219 15033 10276
rect 14987 10116 15033 10173
rect 14763 10013 14809 10070
rect 14763 9954 14809 9967
rect 14953 10070 14987 10109
rect 15257 11446 15272 11458
rect 15435 11757 15481 11770
rect 15211 10940 15257 10997
rect 15211 10837 15257 10894
rect 15211 10734 15257 10791
rect 15211 10631 15257 10688
rect 15211 10528 15257 10585
rect 15211 10425 15257 10482
rect 15211 10322 15257 10379
rect 15211 10219 15257 10276
rect 15211 10116 15257 10173
rect 15033 10070 15068 10109
rect 14953 10013 15068 10070
rect 14953 9967 14987 10013
rect 15033 9967 15068 10013
rect 14953 9863 15068 9967
rect 15435 10940 15481 10997
rect 15435 10837 15481 10894
rect 15435 10734 15481 10791
rect 15435 10631 15481 10688
rect 15435 10528 15481 10585
rect 15435 10425 15481 10482
rect 15435 10322 15481 10379
rect 15435 10219 15481 10276
rect 15435 10116 15481 10173
rect 15211 10013 15257 10070
rect 15211 9954 15257 9967
rect 15401 10070 15435 10109
rect 15659 11757 15705 11890
rect 16556 11859 16568 11911
rect 16620 11905 16706 11911
rect 16620 11859 16649 11905
rect 16695 11859 16706 11905
rect 16556 11840 16706 11859
rect 16779 11958 16825 12598
rect 17049 12824 17064 12836
rect 17003 12585 17049 12598
rect 17273 15474 17288 15486
rect 17451 16572 17497 16585
rect 17436 14996 17451 15008
rect 17660 16572 17736 16602
rect 18332 16654 18408 16682
rect 18332 16602 18344 16654
rect 18396 16602 18408 16654
rect 17660 16530 17675 16572
rect 17721 16530 17736 16572
rect 17660 16478 17672 16530
rect 17724 16478 17736 16530
rect 17660 16406 17675 16478
rect 17721 16406 17736 16478
rect 17660 16354 17672 16406
rect 17724 16354 17736 16406
rect 17660 16282 17675 16354
rect 17721 16282 17736 16354
rect 17660 16230 17672 16282
rect 17724 16230 17736 16282
rect 17660 16158 17675 16230
rect 17721 16158 17736 16230
rect 17660 16106 17672 16158
rect 17724 16106 17736 16158
rect 17660 16034 17675 16106
rect 17721 16034 17736 16106
rect 17660 15982 17672 16034
rect 17724 15982 17736 16034
rect 17660 15910 17675 15982
rect 17721 15910 17736 15982
rect 17660 15858 17672 15910
rect 17724 15858 17736 15910
rect 17660 15786 17675 15858
rect 17721 15786 17736 15858
rect 17660 15734 17672 15786
rect 17724 15734 17736 15786
rect 17660 15662 17675 15734
rect 17721 15662 17736 15734
rect 17660 15610 17672 15662
rect 17724 15610 17736 15662
rect 17660 15538 17675 15610
rect 17721 15538 17736 15610
rect 17660 15486 17672 15538
rect 17724 15486 17736 15538
rect 17660 15474 17675 15486
rect 17497 14996 17512 15008
rect 17436 14944 17448 14996
rect 17500 14944 17512 14996
rect 17436 14872 17451 14944
rect 17497 14872 17512 14944
rect 17436 14820 17448 14872
rect 17500 14820 17512 14872
rect 17436 14748 17451 14820
rect 17497 14748 17512 14820
rect 17436 14696 17448 14748
rect 17500 14696 17512 14748
rect 17436 14624 17451 14696
rect 17497 14624 17512 14696
rect 17436 14572 17448 14624
rect 17500 14572 17512 14624
rect 17436 14500 17451 14572
rect 17497 14500 17512 14572
rect 17436 14448 17448 14500
rect 17500 14448 17512 14500
rect 17436 14376 17451 14448
rect 17497 14376 17512 14448
rect 17436 14324 17448 14376
rect 17500 14324 17512 14376
rect 17436 14252 17451 14324
rect 17497 14252 17512 14324
rect 17436 14200 17448 14252
rect 17500 14200 17512 14252
rect 17436 14128 17451 14200
rect 17497 14128 17512 14200
rect 17436 14076 17448 14128
rect 17500 14076 17512 14128
rect 17436 14004 17451 14076
rect 17497 14004 17512 14076
rect 17436 13952 17448 14004
rect 17500 13952 17512 14004
rect 17436 13880 17451 13952
rect 17497 13880 17512 13952
rect 17436 13828 17448 13880
rect 17500 13828 17512 13880
rect 17436 13756 17451 13828
rect 17497 13756 17512 13828
rect 17436 13704 17448 13756
rect 17500 13704 17512 13756
rect 17436 13632 17451 13704
rect 17497 13632 17512 13704
rect 17436 13580 17448 13632
rect 17500 13580 17512 13632
rect 17436 13508 17451 13580
rect 17497 13508 17512 13580
rect 17436 13456 17448 13508
rect 17500 13456 17512 13508
rect 17436 13384 17451 13456
rect 17497 13384 17512 13456
rect 17436 13332 17448 13384
rect 17500 13332 17512 13384
rect 17436 13260 17451 13332
rect 17497 13260 17512 13332
rect 17436 13208 17448 13260
rect 17500 13208 17512 13260
rect 17436 13136 17451 13208
rect 17497 13136 17512 13208
rect 17436 13084 17448 13136
rect 17500 13084 17512 13136
rect 17436 13012 17451 13084
rect 17497 13012 17512 13084
rect 17436 12960 17448 13012
rect 17500 12960 17512 13012
rect 17436 12888 17451 12960
rect 17497 12888 17512 12960
rect 17436 12836 17448 12888
rect 17500 12836 17512 12888
rect 17436 12824 17451 12836
rect 17227 12274 17273 12598
rect 17497 12824 17512 12836
rect 17451 12585 17497 12598
rect 17721 15474 17736 15486
rect 17899 16572 17945 16585
rect 17675 12585 17721 12598
rect 18123 16572 18169 16585
rect 18108 14996 18123 15008
rect 18332 16572 18408 16602
rect 18780 16654 18856 16682
rect 18780 16602 18792 16654
rect 18844 16602 18856 16654
rect 18332 16530 18347 16572
rect 18393 16530 18408 16572
rect 18332 16478 18344 16530
rect 18396 16478 18408 16530
rect 18332 16406 18347 16478
rect 18393 16406 18408 16478
rect 18332 16354 18344 16406
rect 18396 16354 18408 16406
rect 18332 16282 18347 16354
rect 18393 16282 18408 16354
rect 18332 16230 18344 16282
rect 18396 16230 18408 16282
rect 18332 16158 18347 16230
rect 18393 16158 18408 16230
rect 18332 16106 18344 16158
rect 18396 16106 18408 16158
rect 18332 16034 18347 16106
rect 18393 16034 18408 16106
rect 18332 15982 18344 16034
rect 18396 15982 18408 16034
rect 18332 15910 18347 15982
rect 18393 15910 18408 15982
rect 18332 15858 18344 15910
rect 18396 15858 18408 15910
rect 18332 15786 18347 15858
rect 18393 15786 18408 15858
rect 18332 15734 18344 15786
rect 18396 15734 18408 15786
rect 18332 15662 18347 15734
rect 18393 15662 18408 15734
rect 18332 15610 18344 15662
rect 18396 15610 18408 15662
rect 18332 15538 18347 15610
rect 18393 15538 18408 15610
rect 18332 15486 18344 15538
rect 18396 15486 18408 15538
rect 18332 15474 18347 15486
rect 18169 14996 18184 15008
rect 18108 14944 18120 14996
rect 18172 14944 18184 14996
rect 18108 14872 18123 14944
rect 18169 14872 18184 14944
rect 18108 14820 18120 14872
rect 18172 14820 18184 14872
rect 18108 14748 18123 14820
rect 18169 14748 18184 14820
rect 18108 14696 18120 14748
rect 18172 14696 18184 14748
rect 18108 14624 18123 14696
rect 18169 14624 18184 14696
rect 18108 14572 18120 14624
rect 18172 14572 18184 14624
rect 18108 14500 18123 14572
rect 18169 14500 18184 14572
rect 18108 14448 18120 14500
rect 18172 14448 18184 14500
rect 18108 14376 18123 14448
rect 18169 14376 18184 14448
rect 18108 14324 18120 14376
rect 18172 14324 18184 14376
rect 18108 14252 18123 14324
rect 18169 14252 18184 14324
rect 18108 14200 18120 14252
rect 18172 14200 18184 14252
rect 18108 14128 18123 14200
rect 18169 14128 18184 14200
rect 18108 14076 18120 14128
rect 18172 14076 18184 14128
rect 18108 14004 18123 14076
rect 18169 14004 18184 14076
rect 18108 13952 18120 14004
rect 18172 13952 18184 14004
rect 18108 13880 18123 13952
rect 18169 13880 18184 13952
rect 18108 13828 18120 13880
rect 18172 13828 18184 13880
rect 18108 13756 18123 13828
rect 18169 13756 18184 13828
rect 18108 13704 18120 13756
rect 18172 13704 18184 13756
rect 18108 13632 18123 13704
rect 18169 13632 18184 13704
rect 18108 13580 18120 13632
rect 18172 13580 18184 13632
rect 18108 13508 18123 13580
rect 18169 13508 18184 13580
rect 18108 13456 18120 13508
rect 18172 13456 18184 13508
rect 18108 13384 18123 13456
rect 18169 13384 18184 13456
rect 18108 13332 18120 13384
rect 18172 13332 18184 13384
rect 18108 13260 18123 13332
rect 18169 13260 18184 13332
rect 18108 13208 18120 13260
rect 18172 13208 18184 13260
rect 18108 13136 18123 13208
rect 18169 13136 18184 13208
rect 18108 13084 18120 13136
rect 18172 13084 18184 13136
rect 18108 13012 18123 13084
rect 18169 13012 18184 13084
rect 18108 12960 18120 13012
rect 18172 12960 18184 13012
rect 18108 12888 18123 12960
rect 18169 12888 18184 12960
rect 18108 12836 18120 12888
rect 18172 12836 18184 12888
rect 18108 12824 18123 12836
rect 17465 12458 17627 12469
rect 17465 12412 17476 12458
rect 17616 12412 17627 12458
rect 17465 12401 17627 12412
rect 17758 12427 17826 12438
rect 17135 12263 17391 12274
rect 17135 12217 17146 12263
rect 17380 12217 17391 12263
rect 17135 12206 17391 12217
rect 17562 11958 17608 12401
rect 17758 12381 17769 12427
rect 17815 12381 17826 12427
rect 16779 11947 17627 11958
rect 16779 11901 17476 11947
rect 17616 11901 17627 11947
rect 17758 11923 17826 12381
rect 16779 11890 17627 11901
rect 17676 11911 17826 11923
rect 15868 11758 15944 11770
rect 15868 11706 15880 11758
rect 15932 11706 15944 11758
rect 15868 11634 15883 11706
rect 15929 11634 15944 11706
rect 15868 11582 15880 11634
rect 15932 11582 15944 11634
rect 15868 11510 15883 11582
rect 15929 11510 15944 11582
rect 15868 11458 15880 11510
rect 15932 11458 15944 11510
rect 15868 11446 15883 11458
rect 15659 10940 15705 10997
rect 15659 10837 15705 10894
rect 15659 10734 15705 10791
rect 15659 10631 15705 10688
rect 15659 10528 15705 10585
rect 15659 10425 15705 10482
rect 15659 10322 15705 10379
rect 15659 10219 15705 10276
rect 15659 10116 15705 10173
rect 15481 10070 15516 10109
rect 15401 10013 15516 10070
rect 15401 9967 15435 10013
rect 15481 9967 15516 10013
rect 15401 9863 15516 9967
rect 15659 10013 15705 10070
rect 15659 9954 15705 9967
rect 15929 11446 15944 11458
rect 16107 11757 16153 11770
rect 15883 10940 15929 10997
rect 15883 10837 15929 10894
rect 15883 10734 15929 10791
rect 15883 10631 15929 10688
rect 15883 10528 15929 10585
rect 15883 10425 15929 10482
rect 15883 10322 15929 10379
rect 15883 10219 15929 10276
rect 15883 10116 15929 10173
rect 16316 11758 16392 11770
rect 16316 11706 16328 11758
rect 16380 11706 16392 11758
rect 16316 11634 16331 11706
rect 16377 11634 16392 11706
rect 16316 11582 16328 11634
rect 16380 11582 16392 11634
rect 16316 11510 16331 11582
rect 16377 11510 16392 11582
rect 16316 11458 16328 11510
rect 16380 11458 16392 11510
rect 16316 11446 16331 11458
rect 16107 10940 16153 10997
rect 16107 10837 16153 10894
rect 16107 10734 16153 10791
rect 16107 10631 16153 10688
rect 16107 10528 16153 10585
rect 16107 10425 16153 10482
rect 16107 10322 16153 10379
rect 16107 10219 16153 10276
rect 16107 10116 16153 10173
rect 15883 10013 15929 10070
rect 15883 9954 15929 9967
rect 16073 10070 16107 10109
rect 16377 11446 16392 11458
rect 16555 11757 16601 11770
rect 16331 10940 16377 10997
rect 16331 10837 16377 10894
rect 16331 10734 16377 10791
rect 16331 10631 16377 10688
rect 16331 10528 16377 10585
rect 16331 10425 16377 10482
rect 16331 10322 16377 10379
rect 16331 10219 16377 10276
rect 16331 10116 16377 10173
rect 16153 10070 16188 10109
rect 16073 10013 16188 10070
rect 16073 9967 16107 10013
rect 16153 9967 16188 10013
rect 16073 9863 16188 9967
rect 16555 10940 16601 10997
rect 16555 10837 16601 10894
rect 16555 10734 16601 10791
rect 16555 10631 16601 10688
rect 16555 10528 16601 10585
rect 16555 10425 16601 10482
rect 16555 10322 16601 10379
rect 16555 10219 16601 10276
rect 16555 10116 16601 10173
rect 16331 10013 16377 10070
rect 16331 9954 16377 9967
rect 16521 10070 16555 10109
rect 16779 11757 16825 11890
rect 17676 11859 17688 11911
rect 17740 11905 17826 11911
rect 17740 11859 17769 11905
rect 17815 11859 17826 11905
rect 17676 11840 17826 11859
rect 17899 11958 17945 12598
rect 18169 12824 18184 12836
rect 18123 12585 18169 12598
rect 18393 15474 18408 15486
rect 18571 16572 18617 16585
rect 18556 14996 18571 15008
rect 18780 16572 18856 16602
rect 19452 16654 19528 16682
rect 19452 16602 19464 16654
rect 19516 16602 19528 16654
rect 18780 16530 18795 16572
rect 18841 16530 18856 16572
rect 18780 16478 18792 16530
rect 18844 16478 18856 16530
rect 18780 16406 18795 16478
rect 18841 16406 18856 16478
rect 18780 16354 18792 16406
rect 18844 16354 18856 16406
rect 18780 16282 18795 16354
rect 18841 16282 18856 16354
rect 18780 16230 18792 16282
rect 18844 16230 18856 16282
rect 18780 16158 18795 16230
rect 18841 16158 18856 16230
rect 18780 16106 18792 16158
rect 18844 16106 18856 16158
rect 18780 16034 18795 16106
rect 18841 16034 18856 16106
rect 18780 15982 18792 16034
rect 18844 15982 18856 16034
rect 18780 15910 18795 15982
rect 18841 15910 18856 15982
rect 18780 15858 18792 15910
rect 18844 15858 18856 15910
rect 18780 15786 18795 15858
rect 18841 15786 18856 15858
rect 18780 15734 18792 15786
rect 18844 15734 18856 15786
rect 18780 15662 18795 15734
rect 18841 15662 18856 15734
rect 18780 15610 18792 15662
rect 18844 15610 18856 15662
rect 18780 15538 18795 15610
rect 18841 15538 18856 15610
rect 18780 15486 18792 15538
rect 18844 15486 18856 15538
rect 18780 15474 18795 15486
rect 18617 14996 18632 15008
rect 18556 14944 18568 14996
rect 18620 14944 18632 14996
rect 18556 14872 18571 14944
rect 18617 14872 18632 14944
rect 18556 14820 18568 14872
rect 18620 14820 18632 14872
rect 18556 14748 18571 14820
rect 18617 14748 18632 14820
rect 18556 14696 18568 14748
rect 18620 14696 18632 14748
rect 18556 14624 18571 14696
rect 18617 14624 18632 14696
rect 18556 14572 18568 14624
rect 18620 14572 18632 14624
rect 18556 14500 18571 14572
rect 18617 14500 18632 14572
rect 18556 14448 18568 14500
rect 18620 14448 18632 14500
rect 18556 14376 18571 14448
rect 18617 14376 18632 14448
rect 18556 14324 18568 14376
rect 18620 14324 18632 14376
rect 18556 14252 18571 14324
rect 18617 14252 18632 14324
rect 18556 14200 18568 14252
rect 18620 14200 18632 14252
rect 18556 14128 18571 14200
rect 18617 14128 18632 14200
rect 18556 14076 18568 14128
rect 18620 14076 18632 14128
rect 18556 14004 18571 14076
rect 18617 14004 18632 14076
rect 18556 13952 18568 14004
rect 18620 13952 18632 14004
rect 18556 13880 18571 13952
rect 18617 13880 18632 13952
rect 18556 13828 18568 13880
rect 18620 13828 18632 13880
rect 18556 13756 18571 13828
rect 18617 13756 18632 13828
rect 18556 13704 18568 13756
rect 18620 13704 18632 13756
rect 18556 13632 18571 13704
rect 18617 13632 18632 13704
rect 18556 13580 18568 13632
rect 18620 13580 18632 13632
rect 18556 13508 18571 13580
rect 18617 13508 18632 13580
rect 18556 13456 18568 13508
rect 18620 13456 18632 13508
rect 18556 13384 18571 13456
rect 18617 13384 18632 13456
rect 18556 13332 18568 13384
rect 18620 13332 18632 13384
rect 18556 13260 18571 13332
rect 18617 13260 18632 13332
rect 18556 13208 18568 13260
rect 18620 13208 18632 13260
rect 18556 13136 18571 13208
rect 18617 13136 18632 13208
rect 18556 13084 18568 13136
rect 18620 13084 18632 13136
rect 18556 13012 18571 13084
rect 18617 13012 18632 13084
rect 18556 12960 18568 13012
rect 18620 12960 18632 13012
rect 18556 12888 18571 12960
rect 18617 12888 18632 12960
rect 18556 12836 18568 12888
rect 18620 12836 18632 12888
rect 18556 12824 18571 12836
rect 18347 12274 18393 12598
rect 18617 12824 18632 12836
rect 18571 12585 18617 12598
rect 18841 15474 18856 15486
rect 19019 16572 19065 16585
rect 18795 12585 18841 12598
rect 19243 16572 19289 16585
rect 19228 14996 19243 15008
rect 19452 16572 19528 16602
rect 19900 16654 19976 16682
rect 19900 16602 19912 16654
rect 19964 16602 19976 16654
rect 19452 16530 19467 16572
rect 19513 16530 19528 16572
rect 19452 16478 19464 16530
rect 19516 16478 19528 16530
rect 19452 16406 19467 16478
rect 19513 16406 19528 16478
rect 19452 16354 19464 16406
rect 19516 16354 19528 16406
rect 19452 16282 19467 16354
rect 19513 16282 19528 16354
rect 19452 16230 19464 16282
rect 19516 16230 19528 16282
rect 19452 16158 19467 16230
rect 19513 16158 19528 16230
rect 19452 16106 19464 16158
rect 19516 16106 19528 16158
rect 19452 16034 19467 16106
rect 19513 16034 19528 16106
rect 19452 15982 19464 16034
rect 19516 15982 19528 16034
rect 19452 15910 19467 15982
rect 19513 15910 19528 15982
rect 19452 15858 19464 15910
rect 19516 15858 19528 15910
rect 19452 15786 19467 15858
rect 19513 15786 19528 15858
rect 19452 15734 19464 15786
rect 19516 15734 19528 15786
rect 19452 15662 19467 15734
rect 19513 15662 19528 15734
rect 19452 15610 19464 15662
rect 19516 15610 19528 15662
rect 19452 15538 19467 15610
rect 19513 15538 19528 15610
rect 19452 15486 19464 15538
rect 19516 15486 19528 15538
rect 19452 15474 19467 15486
rect 19289 14996 19304 15008
rect 19228 14944 19240 14996
rect 19292 14944 19304 14996
rect 19228 14872 19243 14944
rect 19289 14872 19304 14944
rect 19228 14820 19240 14872
rect 19292 14820 19304 14872
rect 19228 14748 19243 14820
rect 19289 14748 19304 14820
rect 19228 14696 19240 14748
rect 19292 14696 19304 14748
rect 19228 14624 19243 14696
rect 19289 14624 19304 14696
rect 19228 14572 19240 14624
rect 19292 14572 19304 14624
rect 19228 14500 19243 14572
rect 19289 14500 19304 14572
rect 19228 14448 19240 14500
rect 19292 14448 19304 14500
rect 19228 14376 19243 14448
rect 19289 14376 19304 14448
rect 19228 14324 19240 14376
rect 19292 14324 19304 14376
rect 19228 14252 19243 14324
rect 19289 14252 19304 14324
rect 19228 14200 19240 14252
rect 19292 14200 19304 14252
rect 19228 14128 19243 14200
rect 19289 14128 19304 14200
rect 19228 14076 19240 14128
rect 19292 14076 19304 14128
rect 19228 14004 19243 14076
rect 19289 14004 19304 14076
rect 19228 13952 19240 14004
rect 19292 13952 19304 14004
rect 19228 13880 19243 13952
rect 19289 13880 19304 13952
rect 19228 13828 19240 13880
rect 19292 13828 19304 13880
rect 19228 13756 19243 13828
rect 19289 13756 19304 13828
rect 19228 13704 19240 13756
rect 19292 13704 19304 13756
rect 19228 13632 19243 13704
rect 19289 13632 19304 13704
rect 19228 13580 19240 13632
rect 19292 13580 19304 13632
rect 19228 13508 19243 13580
rect 19289 13508 19304 13580
rect 19228 13456 19240 13508
rect 19292 13456 19304 13508
rect 19228 13384 19243 13456
rect 19289 13384 19304 13456
rect 19228 13332 19240 13384
rect 19292 13332 19304 13384
rect 19228 13260 19243 13332
rect 19289 13260 19304 13332
rect 19228 13208 19240 13260
rect 19292 13208 19304 13260
rect 19228 13136 19243 13208
rect 19289 13136 19304 13208
rect 19228 13084 19240 13136
rect 19292 13084 19304 13136
rect 19228 13012 19243 13084
rect 19289 13012 19304 13084
rect 19228 12960 19240 13012
rect 19292 12960 19304 13012
rect 19228 12888 19243 12960
rect 19289 12888 19304 12960
rect 19228 12836 19240 12888
rect 19292 12836 19304 12888
rect 19228 12824 19243 12836
rect 18585 12458 18747 12469
rect 18585 12412 18596 12458
rect 18736 12412 18747 12458
rect 18585 12401 18747 12412
rect 18878 12427 18946 12438
rect 18255 12263 18511 12274
rect 18255 12217 18266 12263
rect 18500 12217 18511 12263
rect 18255 12206 18511 12217
rect 18682 11958 18728 12401
rect 18878 12381 18889 12427
rect 18935 12381 18946 12427
rect 17899 11947 18747 11958
rect 17899 11901 18596 11947
rect 18736 11901 18747 11947
rect 18878 11923 18946 12381
rect 17899 11890 18747 11901
rect 18796 11911 18946 11923
rect 16988 11758 17064 11770
rect 16988 11706 17000 11758
rect 17052 11706 17064 11758
rect 16988 11634 17003 11706
rect 17049 11634 17064 11706
rect 16988 11582 17000 11634
rect 17052 11582 17064 11634
rect 16988 11510 17003 11582
rect 17049 11510 17064 11582
rect 16988 11458 17000 11510
rect 17052 11458 17064 11510
rect 16988 11446 17003 11458
rect 16779 10940 16825 10997
rect 16779 10837 16825 10894
rect 16779 10734 16825 10791
rect 16779 10631 16825 10688
rect 16779 10528 16825 10585
rect 16779 10425 16825 10482
rect 16779 10322 16825 10379
rect 16779 10219 16825 10276
rect 16779 10116 16825 10173
rect 16601 10070 16636 10109
rect 16521 10013 16636 10070
rect 16521 9967 16555 10013
rect 16601 9967 16636 10013
rect 16521 9863 16636 9967
rect 16779 10013 16825 10070
rect 16779 9954 16825 9967
rect 17049 11446 17064 11458
rect 17227 11757 17273 11770
rect 17003 10940 17049 10997
rect 17003 10837 17049 10894
rect 17003 10734 17049 10791
rect 17003 10631 17049 10688
rect 17003 10528 17049 10585
rect 17003 10425 17049 10482
rect 17003 10322 17049 10379
rect 17003 10219 17049 10276
rect 17003 10116 17049 10173
rect 17436 11758 17512 11770
rect 17436 11706 17448 11758
rect 17500 11706 17512 11758
rect 17436 11634 17451 11706
rect 17497 11634 17512 11706
rect 17436 11582 17448 11634
rect 17500 11582 17512 11634
rect 17436 11510 17451 11582
rect 17497 11510 17512 11582
rect 17436 11458 17448 11510
rect 17500 11458 17512 11510
rect 17436 11446 17451 11458
rect 17227 10940 17273 10997
rect 17227 10837 17273 10894
rect 17227 10734 17273 10791
rect 17227 10631 17273 10688
rect 17227 10528 17273 10585
rect 17227 10425 17273 10482
rect 17227 10322 17273 10379
rect 17227 10219 17273 10276
rect 17227 10116 17273 10173
rect 17003 10013 17049 10070
rect 17003 9954 17049 9967
rect 17193 10070 17227 10109
rect 17497 11446 17512 11458
rect 17675 11757 17721 11770
rect 17451 10940 17497 10997
rect 17451 10837 17497 10894
rect 17451 10734 17497 10791
rect 17451 10631 17497 10688
rect 17451 10528 17497 10585
rect 17451 10425 17497 10482
rect 17451 10322 17497 10379
rect 17451 10219 17497 10276
rect 17451 10116 17497 10173
rect 17273 10070 17308 10109
rect 17193 10013 17308 10070
rect 17193 9967 17227 10013
rect 17273 9967 17308 10013
rect 17193 9863 17308 9967
rect 17675 10940 17721 10997
rect 17675 10837 17721 10894
rect 17675 10734 17721 10791
rect 17675 10631 17721 10688
rect 17675 10528 17721 10585
rect 17675 10425 17721 10482
rect 17675 10322 17721 10379
rect 17675 10219 17721 10276
rect 17675 10116 17721 10173
rect 17451 10013 17497 10070
rect 17451 9954 17497 9967
rect 17641 10070 17675 10109
rect 17899 11757 17945 11890
rect 18796 11859 18808 11911
rect 18860 11905 18946 11911
rect 18860 11859 18889 11905
rect 18935 11859 18946 11905
rect 18796 11840 18946 11859
rect 19019 11958 19065 12598
rect 19289 12824 19304 12836
rect 19243 12585 19289 12598
rect 19513 15474 19528 15486
rect 19691 16572 19737 16585
rect 19676 14996 19691 15008
rect 19900 16572 19976 16602
rect 19900 16530 19915 16572
rect 19961 16530 19976 16572
rect 19900 16478 19912 16530
rect 19964 16478 19976 16530
rect 19900 16406 19915 16478
rect 19961 16406 19976 16478
rect 19900 16354 19912 16406
rect 19964 16354 19976 16406
rect 19900 16282 19915 16354
rect 19961 16282 19976 16354
rect 19900 16230 19912 16282
rect 19964 16230 19976 16282
rect 19900 16158 19915 16230
rect 19961 16158 19976 16230
rect 19900 16106 19912 16158
rect 19964 16106 19976 16158
rect 19900 16034 19915 16106
rect 19961 16034 19976 16106
rect 19900 15982 19912 16034
rect 19964 15982 19976 16034
rect 19900 15910 19915 15982
rect 19961 15910 19976 15982
rect 19900 15858 19912 15910
rect 19964 15858 19976 15910
rect 19900 15786 19915 15858
rect 19961 15786 19976 15858
rect 19900 15734 19912 15786
rect 19964 15734 19976 15786
rect 19900 15662 19915 15734
rect 19961 15662 19976 15734
rect 19900 15610 19912 15662
rect 19964 15610 19976 15662
rect 19900 15538 19915 15610
rect 19961 15538 19976 15610
rect 19900 15486 19912 15538
rect 19964 15486 19976 15538
rect 19900 15474 19915 15486
rect 19737 14996 19752 15008
rect 19676 14944 19688 14996
rect 19740 14944 19752 14996
rect 19676 14872 19691 14944
rect 19737 14872 19752 14944
rect 19676 14820 19688 14872
rect 19740 14820 19752 14872
rect 19676 14748 19691 14820
rect 19737 14748 19752 14820
rect 19676 14696 19688 14748
rect 19740 14696 19752 14748
rect 19676 14624 19691 14696
rect 19737 14624 19752 14696
rect 19676 14572 19688 14624
rect 19740 14572 19752 14624
rect 19676 14500 19691 14572
rect 19737 14500 19752 14572
rect 19676 14448 19688 14500
rect 19740 14448 19752 14500
rect 19676 14376 19691 14448
rect 19737 14376 19752 14448
rect 19676 14324 19688 14376
rect 19740 14324 19752 14376
rect 19676 14252 19691 14324
rect 19737 14252 19752 14324
rect 19676 14200 19688 14252
rect 19740 14200 19752 14252
rect 19676 14128 19691 14200
rect 19737 14128 19752 14200
rect 19676 14076 19688 14128
rect 19740 14076 19752 14128
rect 19676 14004 19691 14076
rect 19737 14004 19752 14076
rect 19676 13952 19688 14004
rect 19740 13952 19752 14004
rect 19676 13880 19691 13952
rect 19737 13880 19752 13952
rect 19676 13828 19688 13880
rect 19740 13828 19752 13880
rect 19676 13756 19691 13828
rect 19737 13756 19752 13828
rect 19676 13704 19688 13756
rect 19740 13704 19752 13756
rect 19676 13632 19691 13704
rect 19737 13632 19752 13704
rect 19676 13580 19688 13632
rect 19740 13580 19752 13632
rect 19676 13508 19691 13580
rect 19737 13508 19752 13580
rect 19676 13456 19688 13508
rect 19740 13456 19752 13508
rect 19676 13384 19691 13456
rect 19737 13384 19752 13456
rect 19676 13332 19688 13384
rect 19740 13332 19752 13384
rect 19676 13260 19691 13332
rect 19737 13260 19752 13332
rect 19676 13208 19688 13260
rect 19740 13208 19752 13260
rect 19676 13136 19691 13208
rect 19737 13136 19752 13208
rect 19676 13084 19688 13136
rect 19740 13084 19752 13136
rect 19676 13012 19691 13084
rect 19737 13012 19752 13084
rect 19676 12960 19688 13012
rect 19740 12960 19752 13012
rect 19676 12888 19691 12960
rect 19737 12888 19752 12960
rect 19676 12836 19688 12888
rect 19740 12836 19752 12888
rect 19676 12824 19691 12836
rect 19467 12274 19513 12598
rect 19737 12824 19752 12836
rect 19691 12585 19737 12598
rect 19961 15474 19976 15486
rect 19915 12585 19961 12598
rect 19705 12458 19867 12469
rect 19705 12412 19716 12458
rect 19856 12412 19867 12458
rect 19705 12401 19867 12412
rect 19375 12263 19631 12274
rect 19375 12217 19386 12263
rect 19620 12217 19631 12263
rect 19375 12206 19631 12217
rect 19802 11958 19848 12401
rect 19019 11947 19867 11958
rect 19019 11901 19716 11947
rect 19856 11901 19867 11947
rect 19019 11890 19867 11901
rect 18108 11758 18184 11770
rect 18108 11706 18120 11758
rect 18172 11706 18184 11758
rect 18108 11634 18123 11706
rect 18169 11634 18184 11706
rect 18108 11582 18120 11634
rect 18172 11582 18184 11634
rect 18108 11510 18123 11582
rect 18169 11510 18184 11582
rect 18108 11458 18120 11510
rect 18172 11458 18184 11510
rect 18108 11446 18123 11458
rect 17899 10940 17945 10997
rect 17899 10837 17945 10894
rect 17899 10734 17945 10791
rect 17899 10631 17945 10688
rect 17899 10528 17945 10585
rect 17899 10425 17945 10482
rect 17899 10322 17945 10379
rect 17899 10219 17945 10276
rect 17899 10116 17945 10173
rect 17721 10070 17756 10109
rect 17641 10013 17756 10070
rect 17641 9967 17675 10013
rect 17721 9967 17756 10013
rect 17641 9863 17756 9967
rect 17899 10013 17945 10070
rect 17899 9954 17945 9967
rect 18169 11446 18184 11458
rect 18347 11757 18393 11770
rect 18123 10940 18169 10997
rect 18123 10837 18169 10894
rect 18123 10734 18169 10791
rect 18123 10631 18169 10688
rect 18123 10528 18169 10585
rect 18123 10425 18169 10482
rect 18123 10322 18169 10379
rect 18123 10219 18169 10276
rect 18123 10116 18169 10173
rect 18556 11758 18632 11770
rect 18556 11706 18568 11758
rect 18620 11706 18632 11758
rect 18556 11634 18571 11706
rect 18617 11634 18632 11706
rect 18556 11582 18568 11634
rect 18620 11582 18632 11634
rect 18556 11510 18571 11582
rect 18617 11510 18632 11582
rect 18556 11458 18568 11510
rect 18620 11458 18632 11510
rect 18556 11446 18571 11458
rect 18347 10940 18393 10997
rect 18347 10837 18393 10894
rect 18347 10734 18393 10791
rect 18347 10631 18393 10688
rect 18347 10528 18393 10585
rect 18347 10425 18393 10482
rect 18347 10322 18393 10379
rect 18347 10219 18393 10276
rect 18347 10116 18393 10173
rect 18123 10013 18169 10070
rect 18123 9954 18169 9967
rect 18313 10070 18347 10109
rect 18617 11446 18632 11458
rect 18795 11757 18841 11770
rect 18571 10940 18617 10997
rect 18571 10837 18617 10894
rect 18571 10734 18617 10791
rect 18571 10631 18617 10688
rect 18571 10528 18617 10585
rect 18571 10425 18617 10482
rect 18571 10322 18617 10379
rect 18571 10219 18617 10276
rect 18571 10116 18617 10173
rect 18393 10070 18428 10109
rect 18313 10013 18428 10070
rect 18313 9967 18347 10013
rect 18393 9967 18428 10013
rect 18313 9863 18428 9967
rect 18795 10940 18841 10997
rect 18795 10837 18841 10894
rect 18795 10734 18841 10791
rect 18795 10631 18841 10688
rect 18795 10528 18841 10585
rect 18795 10425 18841 10482
rect 18795 10322 18841 10379
rect 18795 10219 18841 10276
rect 18795 10116 18841 10173
rect 18571 10013 18617 10070
rect 18571 9954 18617 9967
rect 18761 10070 18795 10109
rect 19019 11757 19065 11890
rect 19228 11758 19304 11770
rect 19228 11706 19240 11758
rect 19292 11706 19304 11758
rect 19228 11634 19243 11706
rect 19289 11634 19304 11706
rect 19228 11582 19240 11634
rect 19292 11582 19304 11634
rect 19228 11510 19243 11582
rect 19289 11510 19304 11582
rect 19228 11458 19240 11510
rect 19292 11458 19304 11510
rect 19228 11446 19243 11458
rect 19019 10940 19065 10997
rect 19019 10837 19065 10894
rect 19019 10734 19065 10791
rect 19019 10631 19065 10688
rect 19019 10528 19065 10585
rect 19019 10425 19065 10482
rect 19019 10322 19065 10379
rect 19019 10219 19065 10276
rect 19019 10116 19065 10173
rect 18841 10070 18876 10109
rect 18761 10013 18876 10070
rect 18761 9967 18795 10013
rect 18841 9967 18876 10013
rect 18761 9863 18876 9967
rect 19019 10013 19065 10070
rect 19019 9954 19065 9967
rect 19289 11446 19304 11458
rect 19467 11757 19513 11770
rect 19243 10940 19289 10997
rect 19243 10837 19289 10894
rect 19243 10734 19289 10791
rect 19243 10631 19289 10688
rect 19243 10528 19289 10585
rect 19243 10425 19289 10482
rect 19243 10322 19289 10379
rect 19243 10219 19289 10276
rect 19243 10116 19289 10173
rect 19676 11758 19752 11770
rect 19676 11706 19688 11758
rect 19740 11706 19752 11758
rect 19676 11634 19691 11706
rect 19737 11634 19752 11706
rect 19676 11582 19688 11634
rect 19740 11582 19752 11634
rect 19676 11510 19691 11582
rect 19737 11510 19752 11582
rect 19676 11458 19688 11510
rect 19740 11458 19752 11510
rect 19676 11446 19691 11458
rect 19467 10940 19513 10997
rect 19467 10837 19513 10894
rect 19467 10734 19513 10791
rect 19467 10631 19513 10688
rect 19467 10528 19513 10585
rect 19467 10425 19513 10482
rect 19467 10322 19513 10379
rect 19467 10219 19513 10276
rect 19467 10116 19513 10173
rect 19243 10013 19289 10070
rect 19243 9954 19289 9967
rect 19433 10070 19467 10109
rect 19737 11446 19752 11458
rect 19915 11757 19961 11770
rect 19691 10940 19737 10997
rect 19691 10837 19737 10894
rect 19691 10734 19737 10791
rect 19691 10631 19737 10688
rect 19691 10528 19737 10585
rect 19691 10425 19737 10482
rect 19691 10322 19737 10379
rect 19691 10219 19737 10276
rect 19691 10116 19737 10173
rect 19513 10070 19548 10109
rect 19433 10013 19548 10070
rect 19433 9967 19467 10013
rect 19513 9967 19548 10013
rect 19433 9863 19548 9967
rect 19915 10940 19961 10997
rect 19915 10837 19961 10894
rect 19915 10734 19961 10791
rect 19915 10631 19961 10688
rect 19915 10528 19961 10585
rect 19915 10425 19961 10482
rect 19915 10322 19961 10379
rect 19915 10219 19961 10276
rect 19915 10116 19961 10173
rect 19691 10013 19737 10070
rect 19691 9954 19737 9967
rect 19881 10070 19915 10109
rect 19961 10070 19996 10109
rect 19881 10013 19996 10070
rect 19881 9967 19915 10013
rect 19961 9967 19996 10013
rect 19881 9863 19996 9967
rect 1960 9862 2076 9863
rect 2632 9862 2748 9863
rect 3080 9862 3196 9863
rect 3752 9862 3868 9863
rect 4200 9862 4316 9863
rect 4872 9862 4988 9863
rect 5320 9862 5436 9863
rect 5992 9862 6108 9863
rect 6440 9862 6556 9863
rect 7112 9862 7228 9863
rect 7560 9862 7676 9863
rect 8232 9862 8348 9863
rect 8680 9862 8796 9863
rect 9352 9862 9468 9863
rect 9800 9862 9916 9863
rect 10472 9862 10588 9863
rect 10920 9862 11036 9863
rect 11592 9862 11708 9863
rect 12040 9862 12156 9863
rect 12712 9862 12828 9863
rect 13160 9862 13276 9863
rect 13832 9862 13948 9863
rect 14280 9862 14396 9863
rect 14952 9862 15068 9863
rect 15400 9862 15516 9863
rect 16072 9862 16188 9863
rect 16520 9862 16636 9863
rect 17191 9862 17308 9863
rect 17639 9862 17756 9863
rect 18311 9862 18428 9863
rect 18759 9862 18876 9863
rect 19431 9862 19548 9863
rect 19879 9862 19996 9863
rect 1934 9669 19996 9862
rect 1934 9623 2443 9669
rect 2489 9623 2601 9669
rect 2647 9623 2759 9669
rect 2805 9623 2917 9669
rect 2963 9623 3075 9669
rect 3121 9623 3233 9669
rect 3279 9623 3392 9669
rect 3438 9623 3550 9669
rect 3596 9623 3708 9669
rect 3754 9623 3866 9669
rect 3912 9623 4024 9669
rect 4070 9623 4182 9669
rect 4228 9623 4340 9669
rect 4386 9623 4498 9669
rect 4544 9623 4656 9669
rect 4702 9623 4815 9669
rect 4861 9623 4973 9669
rect 5019 9623 5131 9669
rect 5177 9623 5289 9669
rect 5335 9623 5447 9669
rect 5493 9623 5605 9669
rect 5651 9623 5763 9669
rect 5809 9623 5921 9669
rect 5967 9623 6079 9669
rect 6125 9623 6238 9669
rect 6284 9623 6396 9669
rect 6442 9623 6554 9669
rect 6600 9623 6712 9669
rect 6758 9623 6870 9669
rect 6916 9623 7028 9669
rect 7074 9623 7186 9669
rect 7232 9623 7344 9669
rect 7390 9623 7502 9669
rect 7548 9623 7661 9669
rect 7707 9623 7819 9669
rect 7865 9623 7977 9669
rect 8023 9623 8135 9669
rect 8181 9623 8293 9669
rect 8339 9623 8451 9669
rect 8497 9623 8609 9669
rect 8655 9623 8767 9669
rect 8813 9623 8925 9669
rect 8971 9623 9084 9669
rect 9130 9623 9242 9669
rect 9288 9623 9400 9669
rect 9446 9623 9558 9669
rect 9604 9623 9716 9669
rect 9762 9623 9874 9669
rect 9920 9623 10032 9669
rect 10078 9623 10190 9669
rect 10236 9623 10348 9669
rect 10394 9623 10507 9669
rect 10553 9623 10665 9669
rect 10711 9623 10823 9669
rect 10869 9623 10981 9669
rect 11027 9623 11139 9669
rect 11185 9623 11297 9669
rect 11343 9623 11455 9669
rect 11501 9623 11613 9669
rect 11659 9623 11771 9669
rect 11817 9623 11930 9669
rect 11976 9623 12088 9669
rect 12134 9623 12246 9669
rect 12292 9623 12404 9669
rect 12450 9623 12562 9669
rect 12608 9623 12720 9669
rect 12766 9623 12878 9669
rect 12924 9623 13036 9669
rect 13082 9623 13195 9669
rect 13241 9623 13353 9669
rect 13399 9623 13511 9669
rect 13557 9623 13669 9669
rect 13715 9623 13827 9669
rect 13873 9623 13985 9669
rect 14031 9623 14143 9669
rect 14189 9623 14301 9669
rect 14347 9623 14459 9669
rect 14505 9623 14618 9669
rect 14664 9623 14776 9669
rect 14822 9623 14934 9669
rect 14980 9623 15092 9669
rect 15138 9623 15250 9669
rect 15296 9623 15408 9669
rect 15454 9623 15566 9669
rect 15612 9623 15724 9669
rect 15770 9623 15882 9669
rect 15928 9623 16041 9669
rect 16087 9623 16199 9669
rect 16245 9623 16357 9669
rect 16403 9623 16515 9669
rect 16561 9623 16673 9669
rect 16719 9623 16831 9669
rect 16877 9623 16989 9669
rect 17035 9623 17147 9669
rect 17193 9623 17305 9669
rect 17351 9623 17464 9669
rect 17510 9623 17622 9669
rect 17668 9623 17780 9669
rect 17826 9623 17938 9669
rect 17984 9623 18096 9669
rect 18142 9623 18254 9669
rect 18300 9623 18412 9669
rect 18458 9623 18570 9669
rect 18616 9623 18728 9669
rect 18774 9623 18887 9669
rect 18933 9623 19045 9669
rect 19091 9623 19203 9669
rect 19249 9623 19361 9669
rect 19407 9623 19519 9669
rect 19565 9623 19677 9669
rect 19723 9623 19835 9669
rect 19881 9623 19996 9669
rect 1934 9613 19996 9623
rect 1934 9364 19995 9613
rect 21015 9604 21061 9788
rect 21463 9604 21509 9789
rect 21911 9604 21957 9796
rect 21015 9558 21957 9604
rect 1934 9312 2404 9364
rect 2456 9312 2611 9364
rect 2663 9312 3131 9364
rect 3183 9312 4095 9364
rect 4147 9312 4302 9364
rect 4354 9312 4822 9364
rect 4874 9312 5786 9364
rect 5838 9312 5993 9364
rect 6045 9312 6513 9364
rect 6565 9343 19995 9364
rect 6565 9312 7558 9343
rect 1934 9297 7558 9312
rect 7604 9324 7716 9343
rect 7604 9297 7671 9324
rect 7762 9297 7874 9343
rect 7920 9297 8032 9343
rect 8078 9324 8212 9343
rect 8078 9297 8119 9324
rect 1934 9272 7671 9297
rect 7723 9272 8119 9297
rect 8171 9297 8212 9324
rect 8258 9297 8370 9343
rect 8416 9297 8528 9343
rect 8574 9324 8686 9343
rect 8619 9297 8686 9324
rect 8732 9297 9191 9343
rect 9237 9324 9349 9343
rect 9237 9297 9304 9324
rect 9395 9297 9507 9343
rect 9553 9297 9665 9343
rect 9711 9324 9845 9343
rect 9711 9297 9752 9324
rect 8171 9272 8567 9297
rect 8619 9272 9304 9297
rect 9356 9272 9752 9297
rect 9804 9297 9845 9324
rect 9891 9297 10003 9343
rect 10049 9297 10161 9343
rect 10207 9324 10319 9343
rect 10252 9297 10319 9324
rect 10365 9297 10825 9343
rect 10871 9324 10983 9343
rect 10871 9297 10938 9324
rect 11029 9297 11141 9343
rect 11187 9297 11299 9343
rect 11345 9324 11479 9343
rect 11345 9297 11386 9324
rect 9804 9272 10200 9297
rect 10252 9272 10938 9297
rect 10990 9272 11386 9297
rect 11438 9297 11479 9324
rect 11525 9297 11637 9343
rect 11683 9297 11795 9343
rect 11841 9324 11953 9343
rect 11886 9297 11953 9324
rect 11999 9297 12459 9343
rect 12505 9324 12617 9343
rect 12505 9297 12572 9324
rect 12663 9297 12775 9343
rect 12821 9297 12933 9343
rect 12979 9324 13113 9343
rect 12979 9297 13020 9324
rect 11438 9272 11834 9297
rect 11886 9272 12572 9297
rect 12624 9272 13020 9297
rect 13072 9297 13113 9324
rect 13159 9297 13271 9343
rect 13317 9297 13429 9343
rect 13475 9324 13587 9343
rect 13520 9297 13587 9324
rect 13633 9297 19995 9343
rect 13072 9272 13468 9297
rect 13520 9272 19995 9297
rect 1934 9257 19995 9272
rect 2270 9152 2701 9257
rect 2270 9146 2621 9152
rect 2270 9107 2404 9146
rect 2270 9061 2317 9107
rect 2363 9094 2404 9107
rect 2456 9094 2611 9146
rect 2667 9106 2701 9152
rect 2663 9094 2701 9106
rect 2363 9061 2701 9094
rect 2270 9048 2701 9061
rect 2270 9002 2621 9048
rect 2667 9002 2701 9048
rect 2270 8944 2701 9002
rect 2270 8898 2317 8944
rect 2363 8928 2621 8944
rect 2363 8898 2404 8928
rect 2270 8876 2404 8898
rect 2456 8876 2611 8928
rect 2667 8898 2701 8944
rect 2663 8876 2701 8898
rect 2270 8840 2701 8876
rect 2270 8794 2621 8840
rect 2667 8794 2701 8840
rect 2270 8780 2701 8794
rect 2270 8734 2317 8780
rect 2363 8736 2701 8780
rect 2363 8734 2621 8736
rect 2270 8710 2621 8734
rect 2270 8658 2404 8710
rect 2456 8658 2611 8710
rect 2667 8690 2701 8736
rect 2663 8658 2701 8690
rect 2270 8631 2701 8658
rect 2270 8617 2621 8631
rect 2270 8571 2317 8617
rect 2363 8585 2621 8617
rect 2667 8585 2701 8631
rect 2363 8571 2701 8585
rect 2270 8526 2701 8571
rect 2270 8480 2621 8526
rect 2667 8480 2701 8526
rect 2270 8421 2701 8480
rect 2270 8375 2621 8421
rect 2667 8375 2701 8421
rect 2270 8316 2701 8375
rect 2845 9152 2891 9165
rect 2845 9048 2891 9106
rect 2845 8944 2891 9002
rect 2845 8840 2891 8898
rect 2845 8736 2891 8794
rect 2845 8631 2891 8690
rect 3093 9152 3221 9257
rect 3093 9146 3135 9152
rect 3181 9146 3221 9152
rect 3093 9094 3131 9146
rect 3183 9094 3221 9146
rect 3093 9048 3221 9094
rect 3093 9002 3135 9048
rect 3181 9002 3221 9048
rect 3093 8944 3221 9002
rect 3093 8928 3135 8944
rect 3181 8928 3221 8944
rect 3093 8876 3131 8928
rect 3183 8876 3221 8928
rect 3093 8840 3221 8876
rect 3093 8794 3135 8840
rect 3181 8794 3221 8840
rect 3093 8736 3221 8794
rect 3093 8710 3135 8736
rect 3181 8710 3221 8736
rect 3093 8658 3131 8710
rect 3183 8658 3221 8710
rect 3093 8631 3221 8658
rect 3093 8618 3135 8631
rect 2845 8526 2891 8585
rect 2845 8421 2891 8480
rect 2845 8326 2891 8375
rect 3181 8618 3221 8631
rect 3359 9152 3405 9165
rect 3359 9048 3405 9106
rect 3359 8944 3405 9002
rect 3359 8840 3405 8898
rect 3359 8736 3405 8794
rect 3359 8631 3405 8690
rect 3135 8526 3181 8585
rect 3135 8421 3181 8480
rect 2270 8270 2621 8316
rect 2667 8270 2701 8316
rect 2270 8265 2701 8270
rect 2810 8316 2925 8326
rect 2810 8270 2845 8316
rect 2891 8270 2925 8316
rect 2621 8257 2667 8265
rect 2366 8176 2706 8183
rect 2810 8176 2925 8270
rect 3135 8316 3181 8375
rect 3359 8526 3405 8585
rect 3359 8421 3405 8480
rect 3359 8326 3405 8375
rect 3961 9152 4392 9257
rect 3961 9146 4312 9152
rect 3961 9107 4095 9146
rect 3961 9061 4008 9107
rect 4054 9094 4095 9107
rect 4147 9094 4302 9146
rect 4358 9106 4392 9152
rect 4354 9094 4392 9106
rect 4054 9061 4392 9094
rect 3961 9048 4392 9061
rect 3961 9002 4312 9048
rect 4358 9002 4392 9048
rect 3961 8944 4392 9002
rect 3961 8898 4008 8944
rect 4054 8928 4312 8944
rect 4054 8898 4095 8928
rect 3961 8876 4095 8898
rect 4147 8876 4302 8928
rect 4358 8898 4392 8944
rect 4354 8876 4392 8898
rect 3961 8840 4392 8876
rect 3961 8794 4312 8840
rect 4358 8794 4392 8840
rect 3961 8780 4392 8794
rect 3961 8734 4008 8780
rect 4054 8736 4392 8780
rect 4054 8734 4312 8736
rect 3961 8710 4312 8734
rect 3961 8658 4095 8710
rect 4147 8658 4302 8710
rect 4358 8690 4392 8736
rect 4354 8658 4392 8690
rect 3961 8631 4392 8658
rect 3961 8617 4312 8631
rect 3961 8571 4008 8617
rect 4054 8585 4312 8617
rect 4358 8585 4392 8631
rect 4054 8571 4392 8585
rect 3961 8526 4392 8571
rect 3961 8480 4312 8526
rect 4358 8480 4392 8526
rect 3961 8421 4392 8480
rect 3961 8375 4312 8421
rect 4358 8375 4392 8421
rect 3135 8257 3181 8270
rect 3324 8316 3439 8326
rect 3324 8270 3359 8316
rect 3405 8270 3439 8316
rect 2366 8142 2723 8176
rect 2366 8090 2404 8142
rect 2456 8139 2616 8142
rect 2668 8139 2723 8142
rect 2456 8093 2484 8139
rect 2530 8093 2616 8139
rect 2688 8093 2723 8139
rect 2456 8090 2616 8093
rect 2668 8090 2723 8093
rect 2366 8056 2723 8090
rect 2810 8139 3233 8176
rect 2810 8093 2994 8139
rect 3040 8093 3152 8139
rect 3198 8093 3233 8139
rect 2810 8056 3233 8093
rect 2366 8050 2706 8056
rect 2621 7967 2667 7977
rect 2296 7964 2701 7967
rect 2296 7931 2621 7964
rect 2221 7894 2621 7931
rect 2221 7848 2256 7894
rect 2302 7848 2621 7894
rect 2667 7920 2701 7964
rect 2810 7964 2925 8056
rect 2667 7879 2714 7920
rect 2810 7902 2845 7964
rect 2221 7731 2621 7848
rect 2676 7827 2714 7879
rect 2221 7685 2256 7731
rect 2302 7685 2621 7731
rect 2221 7568 2621 7685
rect 2667 7662 2714 7827
rect 2676 7610 2714 7662
rect 2221 7522 2256 7568
rect 2302 7522 2621 7568
rect 2221 7405 2621 7522
rect 2667 7444 2714 7610
rect 2221 7359 2256 7405
rect 2302 7359 2621 7405
rect 2676 7392 2714 7444
rect 2221 7242 2621 7359
rect 2221 7196 2256 7242
rect 2302 7196 2621 7242
rect 2667 7226 2714 7392
rect 2221 7078 2621 7196
rect 2676 7174 2714 7226
rect 2221 7032 2256 7078
rect 2302 7032 2621 7078
rect 2221 6915 2621 7032
rect 2667 7008 2714 7174
rect 2676 6956 2714 7008
rect 2221 6869 2256 6915
rect 2302 6869 2621 6915
rect 2221 6752 2621 6869
rect 2667 6791 2714 6956
rect 2221 6706 2256 6752
rect 2302 6706 2621 6752
rect 2676 6739 2714 6791
rect 2221 6588 2621 6706
rect 2221 6542 2256 6588
rect 2302 6542 2621 6588
rect 2221 6425 2621 6542
rect 2221 6379 2256 6425
rect 2302 6379 2621 6425
rect 2221 6262 2621 6379
rect 2221 6216 2256 6262
rect 2302 6216 2621 6262
rect 2221 6098 2621 6216
rect 2221 6052 2256 6098
rect 2302 6052 2621 6098
rect 2221 5935 2621 6052
rect 2221 5889 2256 5935
rect 2302 5889 2621 5935
rect 2221 5772 2621 5889
rect 2221 5726 2256 5772
rect 2302 5726 2621 5772
rect 2221 5609 2621 5726
rect 2221 5563 2256 5609
rect 2302 5563 2621 5609
rect 2221 5446 2621 5563
rect 2221 5400 2256 5446
rect 2302 5400 2621 5446
rect 2221 5363 2621 5400
rect 2296 5268 2621 5363
rect 2667 6699 2714 6739
rect 2667 6698 2708 6699
rect 2667 5268 2701 6698
rect 2296 5263 2701 5268
rect 2803 5574 2845 5614
rect 2891 7902 2925 7964
rect 3135 7964 3181 7977
rect 3100 6699 3135 7920
rect 3324 7964 3439 8270
rect 3961 8316 4392 8375
rect 4536 9152 4582 9165
rect 4536 9048 4582 9106
rect 4536 8944 4582 9002
rect 4536 8840 4582 8898
rect 4536 8736 4582 8794
rect 4536 8631 4582 8690
rect 4784 9152 4912 9257
rect 4784 9146 4826 9152
rect 4872 9146 4912 9152
rect 4784 9094 4822 9146
rect 4874 9094 4912 9146
rect 4784 9048 4912 9094
rect 4784 9002 4826 9048
rect 4872 9002 4912 9048
rect 4784 8944 4912 9002
rect 4784 8928 4826 8944
rect 4872 8928 4912 8944
rect 4784 8876 4822 8928
rect 4874 8876 4912 8928
rect 4784 8840 4912 8876
rect 4784 8794 4826 8840
rect 4872 8794 4912 8840
rect 4784 8736 4912 8794
rect 4784 8710 4826 8736
rect 4872 8710 4912 8736
rect 4784 8658 4822 8710
rect 4874 8658 4912 8710
rect 4784 8631 4912 8658
rect 4784 8618 4826 8631
rect 4536 8526 4582 8585
rect 4536 8421 4582 8480
rect 4536 8326 4582 8375
rect 4872 8618 4912 8631
rect 5050 9152 5096 9165
rect 5050 9048 5096 9106
rect 5050 8944 5096 9002
rect 5050 8840 5096 8898
rect 5050 8736 5096 8794
rect 5050 8631 5096 8690
rect 4826 8526 4872 8585
rect 4826 8421 4872 8480
rect 3961 8270 4312 8316
rect 4358 8270 4392 8316
rect 3961 8265 4392 8270
rect 4501 8316 4616 8326
rect 4501 8270 4536 8316
rect 4582 8270 4616 8316
rect 4312 8257 4358 8265
rect 4057 8176 4397 8183
rect 4501 8176 4616 8270
rect 4826 8316 4872 8375
rect 5050 8526 5096 8585
rect 5050 8421 5096 8480
rect 5050 8326 5096 8375
rect 5652 9152 6083 9257
rect 5652 9146 6003 9152
rect 5652 9107 5786 9146
rect 5652 9061 5699 9107
rect 5745 9094 5786 9107
rect 5838 9094 5993 9146
rect 6049 9106 6083 9152
rect 6045 9094 6083 9106
rect 5745 9061 6083 9094
rect 5652 9048 6083 9061
rect 5652 9002 6003 9048
rect 6049 9002 6083 9048
rect 5652 8944 6083 9002
rect 5652 8898 5699 8944
rect 5745 8928 6003 8944
rect 5745 8898 5786 8928
rect 5652 8876 5786 8898
rect 5838 8876 5993 8928
rect 6049 8898 6083 8944
rect 6045 8876 6083 8898
rect 5652 8840 6083 8876
rect 5652 8794 6003 8840
rect 6049 8794 6083 8840
rect 5652 8780 6083 8794
rect 5652 8734 5699 8780
rect 5745 8736 6083 8780
rect 5745 8734 6003 8736
rect 5652 8710 6003 8734
rect 5652 8658 5786 8710
rect 5838 8658 5993 8710
rect 6049 8690 6083 8736
rect 6045 8658 6083 8690
rect 5652 8631 6083 8658
rect 5652 8617 6003 8631
rect 5652 8571 5699 8617
rect 5745 8585 6003 8617
rect 6049 8585 6083 8631
rect 5745 8571 6083 8585
rect 5652 8526 6083 8571
rect 5652 8480 6003 8526
rect 6049 8480 6083 8526
rect 5652 8421 6083 8480
rect 5652 8375 6003 8421
rect 6049 8375 6083 8421
rect 4826 8257 4872 8270
rect 5015 8316 5130 8326
rect 5015 8270 5050 8316
rect 5096 8270 5130 8316
rect 4057 8142 4414 8176
rect 4057 8090 4095 8142
rect 4147 8139 4307 8142
rect 4359 8139 4414 8142
rect 4147 8093 4175 8139
rect 4221 8093 4307 8139
rect 4379 8093 4414 8139
rect 4147 8090 4307 8093
rect 4359 8090 4414 8093
rect 4057 8056 4414 8090
rect 4501 8139 4924 8176
rect 4501 8093 4685 8139
rect 4731 8093 4843 8139
rect 4889 8093 4924 8139
rect 4501 8056 4924 8093
rect 4057 8050 4397 8056
rect 4312 7967 4358 7977
rect 3181 7879 3228 7920
rect 3324 7902 3359 7964
rect 3190 7827 3228 7879
rect 3181 7662 3228 7827
rect 3190 7610 3228 7662
rect 3181 7444 3228 7610
rect 3190 7392 3228 7444
rect 3181 7226 3228 7392
rect 3190 7174 3228 7226
rect 3181 7008 3228 7174
rect 3190 6956 3228 7008
rect 3181 6791 3228 6956
rect 3190 6739 3228 6791
rect 3106 6698 3135 6699
rect 2891 5574 2932 5614
rect 2803 5522 2841 5574
rect 2893 5522 2932 5574
rect 2803 5356 2845 5522
rect 2891 5356 2932 5522
rect 2803 5304 2841 5356
rect 2893 5304 2932 5356
rect 2803 5268 2845 5304
rect 2891 5268 2932 5304
rect 2621 5255 2667 5263
rect 2803 5161 2932 5268
rect 3181 6699 3228 6739
rect 3181 6698 3222 6699
rect 3135 5255 3181 5268
rect 3319 5574 3359 5614
rect 3405 7902 3439 7964
rect 3987 7964 4392 7967
rect 3987 7931 4312 7964
rect 3912 7894 4312 7931
rect 3912 7848 3947 7894
rect 3993 7848 4312 7894
rect 4358 7920 4392 7964
rect 4501 7964 4616 8056
rect 4358 7879 4405 7920
rect 4501 7902 4536 7964
rect 3912 7731 4312 7848
rect 4367 7827 4405 7879
rect 3912 7685 3947 7731
rect 3993 7685 4312 7731
rect 3912 7568 4312 7685
rect 4358 7662 4405 7827
rect 4367 7610 4405 7662
rect 3912 7522 3947 7568
rect 3993 7522 4312 7568
rect 3912 7405 4312 7522
rect 4358 7444 4405 7610
rect 3912 7359 3947 7405
rect 3993 7359 4312 7405
rect 4367 7392 4405 7444
rect 3912 7242 4312 7359
rect 3912 7196 3947 7242
rect 3993 7196 4312 7242
rect 4358 7226 4405 7392
rect 3912 7078 4312 7196
rect 4367 7174 4405 7226
rect 3912 7032 3947 7078
rect 3993 7032 4312 7078
rect 3912 6915 4312 7032
rect 4358 7008 4405 7174
rect 4367 6956 4405 7008
rect 3912 6869 3947 6915
rect 3993 6869 4312 6915
rect 3912 6752 4312 6869
rect 4358 6791 4405 6956
rect 3912 6706 3947 6752
rect 3993 6706 4312 6752
rect 4367 6739 4405 6791
rect 3912 6588 4312 6706
rect 3912 6542 3947 6588
rect 3993 6542 4312 6588
rect 3912 6425 4312 6542
rect 3912 6379 3947 6425
rect 3993 6379 4312 6425
rect 3912 6262 4312 6379
rect 3912 6216 3947 6262
rect 3993 6216 4312 6262
rect 3912 6098 4312 6216
rect 3912 6052 3947 6098
rect 3993 6052 4312 6098
rect 3912 5935 4312 6052
rect 3912 5889 3947 5935
rect 3993 5889 4312 5935
rect 3912 5772 4312 5889
rect 3912 5726 3947 5772
rect 3993 5726 4312 5772
rect 3405 5574 3443 5614
rect 3319 5522 3355 5574
rect 3407 5522 3443 5574
rect 3319 5356 3359 5522
rect 3405 5356 3443 5522
rect 3912 5609 4312 5726
rect 3912 5563 3947 5609
rect 3993 5563 4312 5609
rect 3912 5446 4312 5563
rect 3912 5400 3947 5446
rect 3993 5400 4312 5446
rect 3912 5363 4312 5400
rect 3319 5304 3355 5356
rect 3407 5304 3443 5356
rect 3319 5268 3359 5304
rect 3405 5268 3443 5304
rect 3319 5264 3443 5268
rect 3987 5268 4312 5363
rect 4358 6699 4405 6739
rect 4358 6698 4399 6699
rect 4358 5268 4392 6698
rect 3359 5255 3405 5264
rect 3987 5263 4392 5268
rect 4496 5574 4536 5614
rect 4582 7902 4616 7964
rect 4826 7964 4872 7977
rect 4791 6699 4826 7920
rect 5015 7964 5130 8270
rect 5652 8316 6083 8375
rect 6227 9152 6273 9165
rect 6227 9048 6273 9106
rect 6227 8944 6273 9002
rect 6227 8840 6273 8898
rect 6227 8736 6273 8794
rect 6227 8631 6273 8690
rect 6475 9152 6603 9257
rect 6475 9146 6517 9152
rect 6563 9146 6603 9152
rect 6475 9094 6513 9146
rect 6565 9094 6603 9146
rect 6475 9048 6603 9094
rect 6475 9002 6517 9048
rect 6563 9002 6603 9048
rect 6475 8944 6603 9002
rect 6475 8928 6517 8944
rect 6563 8928 6603 8944
rect 6475 8876 6513 8928
rect 6565 8876 6603 8928
rect 6475 8840 6603 8876
rect 6475 8794 6517 8840
rect 6563 8794 6603 8840
rect 6475 8736 6603 8794
rect 6475 8710 6517 8736
rect 6563 8710 6603 8736
rect 6475 8658 6513 8710
rect 6565 8658 6603 8710
rect 6475 8631 6603 8658
rect 6475 8618 6517 8631
rect 6227 8526 6273 8585
rect 6227 8421 6273 8480
rect 6227 8326 6273 8375
rect 6563 8618 6603 8631
rect 6741 9152 6787 9165
rect 6741 9048 6787 9106
rect 7327 9106 13864 9257
rect 7327 9102 7671 9106
rect 7633 9054 7671 9102
rect 7723 9102 8119 9106
rect 7723 9054 7761 9102
rect 6741 8944 6787 9002
rect 6741 8840 6787 8898
rect 6741 8736 6787 8794
rect 6741 8631 6787 8690
rect 7450 9008 7496 9021
rect 7450 8880 7496 8962
rect 7450 8753 7496 8834
rect 7450 8650 7496 8707
rect 7633 9008 7761 9054
rect 8081 9054 8119 9102
rect 8171 9102 8567 9106
rect 8171 9054 8209 9102
rect 7898 9012 7944 9021
rect 7633 8962 7674 9008
rect 7720 8962 7761 9008
rect 7633 8888 7761 8962
rect 7633 8836 7671 8888
rect 7723 8836 7761 8888
rect 7633 8834 7674 8836
rect 7720 8834 7761 8836
rect 7633 8753 7761 8834
rect 7633 8707 7674 8753
rect 7720 8707 7761 8753
rect 7633 8670 7761 8707
rect 6517 8526 6563 8585
rect 6517 8421 6563 8480
rect 5652 8270 6003 8316
rect 6049 8270 6083 8316
rect 5652 8265 6083 8270
rect 6192 8316 6307 8326
rect 6192 8270 6227 8316
rect 6273 8270 6307 8316
rect 6003 8257 6049 8265
rect 5748 8176 6088 8183
rect 6192 8176 6307 8270
rect 6517 8316 6563 8375
rect 6741 8526 6787 8585
rect 6741 8421 6787 8480
rect 6741 8326 6787 8375
rect 7416 8626 7531 8650
rect 7416 8580 7450 8626
rect 7496 8580 7531 8626
rect 7416 8491 7531 8580
rect 7633 8618 7671 8670
rect 7723 8618 7761 8670
rect 7633 8580 7674 8618
rect 7720 8580 7761 8618
rect 7633 8578 7761 8580
rect 7859 9008 7987 9012
rect 7859 8973 7898 9008
rect 7944 8973 7987 9008
rect 7859 8921 7897 8973
rect 7949 8921 7987 8973
rect 7859 8880 7987 8921
rect 7859 8834 7898 8880
rect 7944 8834 7987 8880
rect 7859 8755 7987 8834
rect 7859 8703 7897 8755
rect 7949 8703 7987 8755
rect 7859 8626 7987 8703
rect 7859 8580 7898 8626
rect 7944 8580 7987 8626
rect 7674 8567 7720 8578
rect 7859 8537 7987 8580
rect 8081 9008 8209 9054
rect 8529 9054 8567 9102
rect 8619 9102 9304 9106
rect 8619 9054 8657 9102
rect 8346 9012 8392 9021
rect 8081 8962 8122 9008
rect 8168 8962 8209 9008
rect 8081 8888 8209 8962
rect 8081 8836 8119 8888
rect 8171 8836 8209 8888
rect 8081 8834 8122 8836
rect 8168 8834 8209 8836
rect 8081 8753 8209 8834
rect 8081 8707 8122 8753
rect 8168 8707 8209 8753
rect 8081 8670 8209 8707
rect 8081 8618 8119 8670
rect 8171 8618 8209 8670
rect 8081 8580 8122 8618
rect 8168 8580 8209 8618
rect 8081 8578 8209 8580
rect 8303 9008 8431 9012
rect 8303 8973 8346 9008
rect 8392 8973 8431 9008
rect 8303 8921 8341 8973
rect 8393 8921 8431 8973
rect 8303 8880 8431 8921
rect 8303 8834 8346 8880
rect 8392 8834 8431 8880
rect 8303 8755 8431 8834
rect 8303 8703 8341 8755
rect 8393 8703 8431 8755
rect 8303 8626 8431 8703
rect 8303 8580 8346 8626
rect 8392 8580 8431 8626
rect 8122 8567 8168 8578
rect 7859 8491 7897 8537
rect 7416 8485 7897 8491
rect 7949 8485 7987 8537
rect 7416 8445 7987 8485
rect 8303 8537 8431 8580
rect 8529 9008 8657 9054
rect 9266 9054 9304 9102
rect 9356 9102 9752 9106
rect 9356 9054 9394 9102
rect 8529 8962 8570 9008
rect 8616 8962 8657 9008
rect 8529 8888 8657 8962
rect 8529 8836 8567 8888
rect 8619 8836 8657 8888
rect 8529 8834 8570 8836
rect 8616 8834 8657 8836
rect 8529 8753 8657 8834
rect 8529 8707 8570 8753
rect 8616 8707 8657 8753
rect 8529 8670 8657 8707
rect 8529 8618 8567 8670
rect 8619 8618 8657 8670
rect 8794 9008 8840 9021
rect 8794 8880 8840 8962
rect 8794 8753 8840 8834
rect 8794 8650 8840 8707
rect 9083 9008 9129 9021
rect 9083 8880 9129 8962
rect 9083 8753 9129 8834
rect 9083 8650 9129 8707
rect 9266 9008 9394 9054
rect 9714 9054 9752 9102
rect 9804 9102 10200 9106
rect 9804 9054 9842 9102
rect 9531 9012 9577 9021
rect 9266 8962 9307 9008
rect 9353 8962 9394 9008
rect 9266 8888 9394 8962
rect 9266 8836 9304 8888
rect 9356 8836 9394 8888
rect 9266 8834 9307 8836
rect 9353 8834 9394 8836
rect 9266 8753 9394 8834
rect 9266 8707 9307 8753
rect 9353 8707 9394 8753
rect 9266 8670 9394 8707
rect 8529 8580 8570 8618
rect 8616 8580 8657 8618
rect 8529 8578 8657 8580
rect 8759 8626 8874 8650
rect 8759 8580 8794 8626
rect 8840 8580 8874 8626
rect 8570 8567 8616 8578
rect 8303 8485 8341 8537
rect 8393 8491 8431 8537
rect 8759 8491 8874 8580
rect 8393 8485 8874 8491
rect 8303 8445 8874 8485
rect 7416 8444 7979 8445
rect 8311 8444 8874 8445
rect 7416 8372 7978 8444
rect 6517 8257 6563 8270
rect 6706 8316 6821 8326
rect 6706 8270 6741 8316
rect 6787 8270 6821 8316
rect 5748 8142 6105 8176
rect 5748 8090 5786 8142
rect 5838 8139 5998 8142
rect 6050 8139 6105 8142
rect 5838 8093 5866 8139
rect 5912 8093 5998 8139
rect 6070 8093 6105 8139
rect 5838 8090 5998 8093
rect 6050 8090 6105 8093
rect 5748 8056 6105 8090
rect 6192 8139 6615 8176
rect 6192 8093 6376 8139
rect 6422 8093 6534 8139
rect 6580 8093 6615 8139
rect 6192 8056 6615 8093
rect 5748 8050 6088 8056
rect 6003 7967 6049 7977
rect 4872 7879 4919 7920
rect 5015 7902 5050 7964
rect 4881 7827 4919 7879
rect 4872 7662 4919 7827
rect 4881 7610 4919 7662
rect 4872 7444 4919 7610
rect 4881 7392 4919 7444
rect 4872 7226 4919 7392
rect 4881 7174 4919 7226
rect 4872 7008 4919 7174
rect 4881 6956 4919 7008
rect 4872 6791 4919 6956
rect 4881 6739 4919 6791
rect 4797 6698 4826 6699
rect 4582 5574 4620 5614
rect 4496 5522 4532 5574
rect 4584 5522 4620 5574
rect 4496 5356 4536 5522
rect 4582 5356 4620 5522
rect 4496 5304 4532 5356
rect 4584 5304 4620 5356
rect 4496 5268 4536 5304
rect 4582 5268 4620 5304
rect 4496 5264 4620 5268
rect 4872 6699 4919 6739
rect 4872 6698 4913 6699
rect 4312 5255 4358 5263
rect 4536 5255 4582 5264
rect 4826 5255 4872 5268
rect 5010 5574 5050 5614
rect 5096 7902 5130 7964
rect 5678 7964 6083 7967
rect 5678 7931 6003 7964
rect 5603 7894 6003 7931
rect 5603 7848 5638 7894
rect 5684 7848 6003 7894
rect 6049 7920 6083 7964
rect 6192 7964 6307 8056
rect 6049 7879 6096 7920
rect 6192 7902 6227 7964
rect 5603 7731 6003 7848
rect 6058 7827 6096 7879
rect 5603 7685 5638 7731
rect 5684 7685 6003 7731
rect 5603 7568 6003 7685
rect 6049 7662 6096 7827
rect 6058 7610 6096 7662
rect 5603 7522 5638 7568
rect 5684 7522 6003 7568
rect 5603 7405 6003 7522
rect 6049 7444 6096 7610
rect 5603 7359 5638 7405
rect 5684 7359 6003 7405
rect 6058 7392 6096 7444
rect 5603 7242 6003 7359
rect 5603 7196 5638 7242
rect 5684 7196 6003 7242
rect 6049 7226 6096 7392
rect 5603 7078 6003 7196
rect 6058 7174 6096 7226
rect 5603 7032 5638 7078
rect 5684 7032 6003 7078
rect 5603 6915 6003 7032
rect 6049 7008 6096 7174
rect 6058 6956 6096 7008
rect 5603 6869 5638 6915
rect 5684 6869 6003 6915
rect 5603 6752 6003 6869
rect 6049 6791 6096 6956
rect 5603 6706 5638 6752
rect 5684 6706 6003 6752
rect 6058 6739 6096 6791
rect 5603 6588 6003 6706
rect 5603 6542 5638 6588
rect 5684 6542 6003 6588
rect 5603 6425 6003 6542
rect 5603 6379 5638 6425
rect 5684 6379 6003 6425
rect 5603 6262 6003 6379
rect 5603 6216 5638 6262
rect 5684 6216 6003 6262
rect 5603 6098 6003 6216
rect 5603 6052 5638 6098
rect 5684 6052 6003 6098
rect 5603 5935 6003 6052
rect 5603 5889 5638 5935
rect 5684 5889 6003 5935
rect 5603 5772 6003 5889
rect 5603 5726 5638 5772
rect 5684 5726 6003 5772
rect 5096 5574 5134 5614
rect 5010 5522 5046 5574
rect 5098 5522 5134 5574
rect 5010 5356 5050 5522
rect 5096 5356 5134 5522
rect 5603 5609 6003 5726
rect 5603 5563 5638 5609
rect 5684 5563 6003 5609
rect 5603 5446 6003 5563
rect 5603 5400 5638 5446
rect 5684 5400 6003 5446
rect 5603 5363 6003 5400
rect 5010 5304 5046 5356
rect 5098 5304 5134 5356
rect 5010 5268 5050 5304
rect 5096 5268 5134 5304
rect 5010 5264 5134 5268
rect 5678 5268 6003 5363
rect 6049 6699 6096 6739
rect 6049 6698 6090 6699
rect 6049 5268 6083 6698
rect 5050 5255 5096 5264
rect 5678 5263 6083 5268
rect 6187 5574 6227 5614
rect 6273 7902 6307 7964
rect 6517 7964 6563 7977
rect 6482 6699 6517 7920
rect 6706 7964 6821 8270
rect 7416 8273 7531 8372
rect 7863 8371 7978 8372
rect 7416 8227 7450 8273
rect 7496 8227 7531 8273
rect 7674 8273 7720 8286
rect 7864 8273 7978 8371
rect 8312 8372 8874 8444
rect 8312 8371 8427 8372
rect 7864 8227 7898 8273
rect 7944 8227 7978 8273
rect 8122 8273 8168 8286
rect 8312 8273 8426 8371
rect 8312 8227 8346 8273
rect 8392 8227 8426 8273
rect 8570 8273 8616 8286
rect 8759 8273 8874 8372
rect 8759 8227 8794 8273
rect 8840 8227 8874 8273
rect 9049 8626 9164 8650
rect 9049 8580 9083 8626
rect 9129 8580 9164 8626
rect 9049 8491 9164 8580
rect 9266 8618 9304 8670
rect 9356 8618 9394 8670
rect 9266 8580 9307 8618
rect 9353 8580 9394 8618
rect 9266 8578 9394 8580
rect 9492 9008 9620 9012
rect 9492 8973 9531 9008
rect 9577 8973 9620 9008
rect 9492 8921 9530 8973
rect 9582 8921 9620 8973
rect 9492 8880 9620 8921
rect 9492 8834 9531 8880
rect 9577 8834 9620 8880
rect 9492 8755 9620 8834
rect 9492 8703 9530 8755
rect 9582 8703 9620 8755
rect 9492 8626 9620 8703
rect 9492 8580 9531 8626
rect 9577 8580 9620 8626
rect 9307 8567 9353 8578
rect 9492 8537 9620 8580
rect 9714 9008 9842 9054
rect 10162 9054 10200 9102
rect 10252 9102 10938 9106
rect 10252 9054 10290 9102
rect 9979 9012 10025 9021
rect 9714 8962 9755 9008
rect 9801 8962 9842 9008
rect 9714 8888 9842 8962
rect 9714 8836 9752 8888
rect 9804 8836 9842 8888
rect 9714 8834 9755 8836
rect 9801 8834 9842 8836
rect 9714 8753 9842 8834
rect 9714 8707 9755 8753
rect 9801 8707 9842 8753
rect 9714 8670 9842 8707
rect 9714 8618 9752 8670
rect 9804 8618 9842 8670
rect 9714 8580 9755 8618
rect 9801 8580 9842 8618
rect 9714 8578 9842 8580
rect 9936 9008 10064 9012
rect 9936 8973 9979 9008
rect 10025 8973 10064 9008
rect 9936 8921 9974 8973
rect 10026 8921 10064 8973
rect 9936 8880 10064 8921
rect 9936 8834 9979 8880
rect 10025 8834 10064 8880
rect 9936 8755 10064 8834
rect 9936 8703 9974 8755
rect 10026 8703 10064 8755
rect 9936 8626 10064 8703
rect 9936 8580 9979 8626
rect 10025 8580 10064 8626
rect 9755 8567 9801 8578
rect 9492 8491 9530 8537
rect 9049 8485 9530 8491
rect 9582 8485 9620 8537
rect 9049 8445 9620 8485
rect 9936 8537 10064 8580
rect 10162 9008 10290 9054
rect 10900 9054 10938 9102
rect 10990 9102 11386 9106
rect 10990 9054 11028 9102
rect 10162 8962 10203 9008
rect 10249 8962 10290 9008
rect 10162 8888 10290 8962
rect 10162 8836 10200 8888
rect 10252 8836 10290 8888
rect 10162 8834 10203 8836
rect 10249 8834 10290 8836
rect 10162 8753 10290 8834
rect 10162 8707 10203 8753
rect 10249 8707 10290 8753
rect 10162 8670 10290 8707
rect 10162 8618 10200 8670
rect 10252 8618 10290 8670
rect 10427 9008 10473 9021
rect 10427 8880 10473 8962
rect 10427 8753 10473 8834
rect 10427 8650 10473 8707
rect 10717 9008 10763 9021
rect 10717 8880 10763 8962
rect 10717 8753 10763 8834
rect 10717 8650 10763 8707
rect 10900 9008 11028 9054
rect 11348 9054 11386 9102
rect 11438 9102 11834 9106
rect 11438 9054 11476 9102
rect 11165 9012 11211 9021
rect 10900 8962 10941 9008
rect 10987 8962 11028 9008
rect 10900 8888 11028 8962
rect 10900 8836 10938 8888
rect 10990 8836 11028 8888
rect 10900 8834 10941 8836
rect 10987 8834 11028 8836
rect 10900 8753 11028 8834
rect 10900 8707 10941 8753
rect 10987 8707 11028 8753
rect 10900 8670 11028 8707
rect 10162 8580 10203 8618
rect 10249 8580 10290 8618
rect 10162 8578 10290 8580
rect 10392 8626 10507 8650
rect 10392 8580 10427 8626
rect 10473 8580 10507 8626
rect 10203 8567 10249 8578
rect 9936 8485 9974 8537
rect 10026 8491 10064 8537
rect 10392 8491 10507 8580
rect 10026 8485 10507 8491
rect 9936 8445 10507 8485
rect 9049 8444 9612 8445
rect 9944 8444 10507 8445
rect 9049 8372 9611 8444
rect 9049 8273 9164 8372
rect 9496 8371 9611 8372
rect 9049 8227 9083 8273
rect 9129 8227 9164 8273
rect 9307 8273 9353 8286
rect 9497 8273 9611 8371
rect 9945 8372 10507 8444
rect 9945 8371 10060 8372
rect 9497 8227 9531 8273
rect 9577 8227 9611 8273
rect 9755 8273 9801 8286
rect 9945 8273 10059 8371
rect 9945 8227 9979 8273
rect 10025 8227 10059 8273
rect 10203 8273 10249 8286
rect 10392 8273 10507 8372
rect 10392 8227 10427 8273
rect 10473 8227 10507 8273
rect 10683 8626 10798 8650
rect 10683 8580 10717 8626
rect 10763 8580 10798 8626
rect 10683 8491 10798 8580
rect 10900 8618 10938 8670
rect 10990 8618 11028 8670
rect 10900 8580 10941 8618
rect 10987 8580 11028 8618
rect 10900 8578 11028 8580
rect 11126 9008 11254 9012
rect 11126 8973 11165 9008
rect 11211 8973 11254 9008
rect 11126 8921 11164 8973
rect 11216 8921 11254 8973
rect 11126 8880 11254 8921
rect 11126 8834 11165 8880
rect 11211 8834 11254 8880
rect 11126 8755 11254 8834
rect 11126 8703 11164 8755
rect 11216 8703 11254 8755
rect 11126 8626 11254 8703
rect 11126 8580 11165 8626
rect 11211 8580 11254 8626
rect 10941 8567 10987 8578
rect 11126 8537 11254 8580
rect 11348 9008 11476 9054
rect 11796 9054 11834 9102
rect 11886 9102 12572 9106
rect 11886 9054 11924 9102
rect 11613 9012 11659 9021
rect 11348 8962 11389 9008
rect 11435 8962 11476 9008
rect 11348 8888 11476 8962
rect 11348 8836 11386 8888
rect 11438 8836 11476 8888
rect 11348 8834 11389 8836
rect 11435 8834 11476 8836
rect 11348 8753 11476 8834
rect 11348 8707 11389 8753
rect 11435 8707 11476 8753
rect 11348 8670 11476 8707
rect 11348 8618 11386 8670
rect 11438 8618 11476 8670
rect 11348 8580 11389 8618
rect 11435 8580 11476 8618
rect 11348 8578 11476 8580
rect 11570 9008 11698 9012
rect 11570 8973 11613 9008
rect 11659 8973 11698 9008
rect 11570 8921 11608 8973
rect 11660 8921 11698 8973
rect 11570 8880 11698 8921
rect 11570 8834 11613 8880
rect 11659 8834 11698 8880
rect 11570 8755 11698 8834
rect 11570 8703 11608 8755
rect 11660 8703 11698 8755
rect 11570 8626 11698 8703
rect 11570 8580 11613 8626
rect 11659 8580 11698 8626
rect 11389 8567 11435 8578
rect 11126 8491 11164 8537
rect 10683 8485 11164 8491
rect 11216 8485 11254 8537
rect 10683 8445 11254 8485
rect 11570 8537 11698 8580
rect 11796 9008 11924 9054
rect 12534 9054 12572 9102
rect 12624 9102 13020 9106
rect 12624 9054 12662 9102
rect 11796 8962 11837 9008
rect 11883 8962 11924 9008
rect 11796 8888 11924 8962
rect 11796 8836 11834 8888
rect 11886 8836 11924 8888
rect 11796 8834 11837 8836
rect 11883 8834 11924 8836
rect 11796 8753 11924 8834
rect 11796 8707 11837 8753
rect 11883 8707 11924 8753
rect 11796 8670 11924 8707
rect 11796 8618 11834 8670
rect 11886 8618 11924 8670
rect 12061 9008 12107 9021
rect 12061 8880 12107 8962
rect 12061 8753 12107 8834
rect 12061 8650 12107 8707
rect 12351 9008 12397 9021
rect 12351 8880 12397 8962
rect 12351 8753 12397 8834
rect 12351 8650 12397 8707
rect 12534 9008 12662 9054
rect 12982 9054 13020 9102
rect 13072 9102 13468 9106
rect 13072 9054 13110 9102
rect 12799 9012 12845 9021
rect 12534 8962 12575 9008
rect 12621 8962 12662 9008
rect 12534 8888 12662 8962
rect 12534 8836 12572 8888
rect 12624 8836 12662 8888
rect 12534 8834 12575 8836
rect 12621 8834 12662 8836
rect 12534 8753 12662 8834
rect 12534 8707 12575 8753
rect 12621 8707 12662 8753
rect 12534 8670 12662 8707
rect 11796 8580 11837 8618
rect 11883 8580 11924 8618
rect 11796 8578 11924 8580
rect 12026 8626 12141 8650
rect 12026 8580 12061 8626
rect 12107 8580 12141 8626
rect 11837 8567 11883 8578
rect 11570 8485 11608 8537
rect 11660 8491 11698 8537
rect 12026 8491 12141 8580
rect 11660 8485 12141 8491
rect 11570 8445 12141 8485
rect 10683 8444 11246 8445
rect 11578 8444 12141 8445
rect 10683 8372 11245 8444
rect 10683 8273 10798 8372
rect 11130 8371 11245 8372
rect 10683 8227 10717 8273
rect 10763 8227 10798 8273
rect 10941 8273 10987 8286
rect 11131 8273 11245 8371
rect 11579 8372 12141 8444
rect 11579 8371 11694 8372
rect 11131 8227 11165 8273
rect 11211 8227 11245 8273
rect 11389 8273 11435 8286
rect 11579 8273 11693 8371
rect 11579 8227 11613 8273
rect 11659 8227 11693 8273
rect 11837 8273 11883 8286
rect 12026 8273 12141 8372
rect 12026 8227 12061 8273
rect 12107 8227 12141 8273
rect 12317 8626 12432 8650
rect 12317 8580 12351 8626
rect 12397 8580 12432 8626
rect 12317 8491 12432 8580
rect 12534 8618 12572 8670
rect 12624 8618 12662 8670
rect 12534 8580 12575 8618
rect 12621 8580 12662 8618
rect 12534 8578 12662 8580
rect 12760 9008 12888 9012
rect 12760 8973 12799 9008
rect 12845 8973 12888 9008
rect 12760 8921 12798 8973
rect 12850 8921 12888 8973
rect 12760 8880 12888 8921
rect 12760 8834 12799 8880
rect 12845 8834 12888 8880
rect 12760 8755 12888 8834
rect 12760 8703 12798 8755
rect 12850 8703 12888 8755
rect 12760 8626 12888 8703
rect 12760 8580 12799 8626
rect 12845 8580 12888 8626
rect 12575 8567 12621 8578
rect 12760 8537 12888 8580
rect 12982 9008 13110 9054
rect 13430 9054 13468 9102
rect 13520 9102 13864 9106
rect 13520 9054 13558 9102
rect 13247 9012 13293 9021
rect 12982 8962 13023 9008
rect 13069 8962 13110 9008
rect 12982 8888 13110 8962
rect 12982 8836 13020 8888
rect 13072 8836 13110 8888
rect 12982 8834 13023 8836
rect 13069 8834 13110 8836
rect 12982 8753 13110 8834
rect 12982 8707 13023 8753
rect 13069 8707 13110 8753
rect 12982 8670 13110 8707
rect 12982 8618 13020 8670
rect 13072 8618 13110 8670
rect 12982 8580 13023 8618
rect 13069 8580 13110 8618
rect 12982 8578 13110 8580
rect 13204 9008 13332 9012
rect 13204 8973 13247 9008
rect 13293 8973 13332 9008
rect 13204 8921 13242 8973
rect 13294 8921 13332 8973
rect 13204 8880 13332 8921
rect 13204 8834 13247 8880
rect 13293 8834 13332 8880
rect 13204 8755 13332 8834
rect 13204 8703 13242 8755
rect 13294 8703 13332 8755
rect 13204 8626 13332 8703
rect 13204 8580 13247 8626
rect 13293 8580 13332 8626
rect 13023 8567 13069 8578
rect 12760 8491 12798 8537
rect 12317 8485 12798 8491
rect 12850 8485 12888 8537
rect 12317 8445 12888 8485
rect 13204 8537 13332 8580
rect 13430 9008 13558 9054
rect 13430 8962 13471 9008
rect 13517 8962 13558 9008
rect 13430 8888 13558 8962
rect 13430 8836 13468 8888
rect 13520 8836 13558 8888
rect 13430 8834 13471 8836
rect 13517 8834 13558 8836
rect 13430 8753 13558 8834
rect 13430 8707 13471 8753
rect 13517 8707 13558 8753
rect 13430 8670 13558 8707
rect 13430 8618 13468 8670
rect 13520 8618 13558 8670
rect 13695 9008 13741 9021
rect 13695 8880 13741 8962
rect 13695 8753 13741 8834
rect 13695 8650 13741 8707
rect 13430 8580 13471 8618
rect 13517 8580 13558 8618
rect 13430 8578 13558 8580
rect 13660 8626 13775 8650
rect 13660 8580 13695 8626
rect 13741 8580 13775 8626
rect 13471 8567 13517 8578
rect 13204 8485 13242 8537
rect 13294 8491 13332 8537
rect 13660 8491 13775 8580
rect 13294 8485 13775 8491
rect 13204 8445 13775 8485
rect 12317 8444 12880 8445
rect 13212 8444 13775 8445
rect 12317 8372 12879 8444
rect 12317 8273 12432 8372
rect 12764 8371 12879 8372
rect 12317 8227 12351 8273
rect 12397 8227 12432 8273
rect 12575 8273 12621 8286
rect 12765 8273 12879 8371
rect 13213 8372 13775 8444
rect 13213 8371 13328 8372
rect 12765 8227 12799 8273
rect 12845 8227 12879 8273
rect 13023 8273 13069 8286
rect 13213 8273 13327 8371
rect 13213 8227 13247 8273
rect 13293 8227 13327 8273
rect 13471 8273 13517 8286
rect 13660 8273 13775 8372
rect 13660 8227 13695 8273
rect 13741 8227 13775 8273
rect 6563 7879 6610 7920
rect 6706 7902 6741 7964
rect 6572 7827 6610 7879
rect 6563 7662 6610 7827
rect 6572 7610 6610 7662
rect 6563 7444 6610 7610
rect 6572 7392 6610 7444
rect 6563 7226 6610 7392
rect 6572 7174 6610 7226
rect 6563 7008 6610 7174
rect 6572 6956 6610 7008
rect 6563 6791 6610 6956
rect 6572 6739 6610 6791
rect 6488 6698 6517 6699
rect 6273 5574 6311 5614
rect 6187 5522 6223 5574
rect 6275 5522 6311 5574
rect 6187 5356 6227 5522
rect 6273 5356 6311 5522
rect 6187 5304 6223 5356
rect 6275 5304 6311 5356
rect 6187 5268 6227 5304
rect 6273 5268 6311 5304
rect 6187 5264 6311 5268
rect 6563 6699 6610 6739
rect 6563 6698 6604 6699
rect 6003 5255 6049 5263
rect 6227 5255 6273 5264
rect 6517 5255 6563 5268
rect 6701 5574 6741 5614
rect 6787 7902 6821 7964
rect 7450 8164 7496 8227
rect 7450 8055 7496 8118
rect 7450 7947 7496 8009
rect 7450 7839 7496 7901
rect 7674 8164 7720 8227
rect 7674 8055 7720 8118
rect 7674 7947 7720 8009
rect 7674 7858 7720 7901
rect 7898 8164 7944 8227
rect 7898 8055 7944 8118
rect 7898 7947 7944 8009
rect 7450 7731 7496 7793
rect 7450 7623 7496 7685
rect 7450 7515 7496 7577
rect 7450 7407 7496 7469
rect 7450 7299 7496 7361
rect 7633 7839 7761 7858
rect 7633 7819 7674 7839
rect 7720 7819 7761 7839
rect 7633 7767 7671 7819
rect 7723 7767 7761 7819
rect 7633 7731 7761 7767
rect 7633 7685 7674 7731
rect 7720 7685 7761 7731
rect 7633 7623 7761 7685
rect 7633 7601 7674 7623
rect 7720 7601 7761 7623
rect 7633 7549 7671 7601
rect 7723 7549 7761 7601
rect 7633 7515 7761 7549
rect 7633 7469 7674 7515
rect 7720 7469 7761 7515
rect 7633 7407 7761 7469
rect 7633 7383 7674 7407
rect 7720 7383 7761 7407
rect 7633 7331 7671 7383
rect 7723 7331 7761 7383
rect 7633 7299 7761 7331
rect 7633 7291 7674 7299
rect 7450 7191 7496 7253
rect 7450 7132 7496 7145
rect 7720 7291 7761 7299
rect 7898 7839 7944 7901
rect 8122 8164 8168 8227
rect 8122 8055 8168 8118
rect 8122 7947 8168 8009
rect 8122 7858 8168 7901
rect 8346 8164 8392 8227
rect 8346 8055 8392 8118
rect 8346 7947 8392 8009
rect 7898 7731 7944 7793
rect 7898 7623 7944 7685
rect 7898 7515 7944 7577
rect 7898 7407 7944 7469
rect 7898 7299 7944 7361
rect 7674 7191 7720 7253
rect 7674 7132 7720 7145
rect 8081 7839 8209 7858
rect 8081 7819 8122 7839
rect 8168 7819 8209 7839
rect 8081 7767 8119 7819
rect 8171 7767 8209 7819
rect 8081 7731 8209 7767
rect 8081 7685 8122 7731
rect 8168 7685 8209 7731
rect 8081 7623 8209 7685
rect 8081 7601 8122 7623
rect 8168 7601 8209 7623
rect 8081 7549 8119 7601
rect 8171 7549 8209 7601
rect 8081 7515 8209 7549
rect 8081 7469 8122 7515
rect 8168 7469 8209 7515
rect 8081 7407 8209 7469
rect 8081 7383 8122 7407
rect 8168 7383 8209 7407
rect 8081 7331 8119 7383
rect 8171 7331 8209 7383
rect 8081 7299 8209 7331
rect 8081 7291 8122 7299
rect 7898 7191 7944 7253
rect 7898 7132 7944 7145
rect 8168 7291 8209 7299
rect 8346 7839 8392 7901
rect 8570 8164 8616 8227
rect 8570 8055 8616 8118
rect 8570 7947 8616 8009
rect 8570 7858 8616 7901
rect 8794 8164 8840 8227
rect 8794 8055 8840 8118
rect 8794 7947 8840 8009
rect 8346 7731 8392 7793
rect 8346 7623 8392 7685
rect 8346 7515 8392 7577
rect 8346 7407 8392 7469
rect 8346 7299 8392 7361
rect 8122 7191 8168 7253
rect 8122 7132 8168 7145
rect 8529 7839 8657 7858
rect 8529 7819 8570 7839
rect 8616 7819 8657 7839
rect 8529 7767 8567 7819
rect 8619 7767 8657 7819
rect 8529 7731 8657 7767
rect 8529 7685 8570 7731
rect 8616 7685 8657 7731
rect 8529 7623 8657 7685
rect 8529 7601 8570 7623
rect 8616 7601 8657 7623
rect 8529 7549 8567 7601
rect 8619 7549 8657 7601
rect 8529 7515 8657 7549
rect 8529 7469 8570 7515
rect 8616 7469 8657 7515
rect 8529 7407 8657 7469
rect 8529 7383 8570 7407
rect 8616 7383 8657 7407
rect 8529 7331 8567 7383
rect 8619 7331 8657 7383
rect 8529 7299 8657 7331
rect 8529 7291 8570 7299
rect 8346 7191 8392 7253
rect 8346 7132 8392 7145
rect 8616 7291 8657 7299
rect 8794 7839 8840 7901
rect 8794 7731 8840 7793
rect 8794 7623 8840 7685
rect 8794 7515 8840 7577
rect 8794 7407 8840 7469
rect 8794 7299 8840 7361
rect 8570 7191 8616 7253
rect 8570 7132 8616 7145
rect 8794 7191 8840 7253
rect 8794 7132 8840 7145
rect 9083 8164 9129 8227
rect 9083 8055 9129 8118
rect 9083 7947 9129 8009
rect 9083 7839 9129 7901
rect 9307 8164 9353 8227
rect 9307 8055 9353 8118
rect 9307 7947 9353 8009
rect 9307 7858 9353 7901
rect 9531 8164 9577 8227
rect 9531 8055 9577 8118
rect 9531 7947 9577 8009
rect 9083 7731 9129 7793
rect 9083 7623 9129 7685
rect 9083 7515 9129 7577
rect 9083 7407 9129 7469
rect 9083 7299 9129 7361
rect 9266 7839 9394 7858
rect 9266 7819 9307 7839
rect 9353 7819 9394 7839
rect 9266 7767 9304 7819
rect 9356 7767 9394 7819
rect 9266 7731 9394 7767
rect 9266 7685 9307 7731
rect 9353 7685 9394 7731
rect 9266 7623 9394 7685
rect 9266 7601 9307 7623
rect 9353 7601 9394 7623
rect 9266 7549 9304 7601
rect 9356 7549 9394 7601
rect 9266 7515 9394 7549
rect 9266 7469 9307 7515
rect 9353 7469 9394 7515
rect 9266 7407 9394 7469
rect 9266 7383 9307 7407
rect 9353 7383 9394 7407
rect 9266 7331 9304 7383
rect 9356 7331 9394 7383
rect 9266 7299 9394 7331
rect 9266 7291 9307 7299
rect 9083 7191 9129 7253
rect 9083 7132 9129 7145
rect 9353 7291 9394 7299
rect 9531 7839 9577 7901
rect 9755 8164 9801 8227
rect 9755 8055 9801 8118
rect 9755 7947 9801 8009
rect 9755 7858 9801 7901
rect 9979 8164 10025 8227
rect 9979 8055 10025 8118
rect 9979 7947 10025 8009
rect 9531 7731 9577 7793
rect 9531 7623 9577 7685
rect 9531 7515 9577 7577
rect 9531 7407 9577 7469
rect 9531 7299 9577 7361
rect 9307 7191 9353 7253
rect 9307 7132 9353 7145
rect 9714 7839 9842 7858
rect 9714 7819 9755 7839
rect 9801 7819 9842 7839
rect 9714 7767 9752 7819
rect 9804 7767 9842 7819
rect 9714 7731 9842 7767
rect 9714 7685 9755 7731
rect 9801 7685 9842 7731
rect 9714 7623 9842 7685
rect 9714 7601 9755 7623
rect 9801 7601 9842 7623
rect 9714 7549 9752 7601
rect 9804 7549 9842 7601
rect 9714 7515 9842 7549
rect 9714 7469 9755 7515
rect 9801 7469 9842 7515
rect 9714 7407 9842 7469
rect 9714 7383 9755 7407
rect 9801 7383 9842 7407
rect 9714 7331 9752 7383
rect 9804 7331 9842 7383
rect 9714 7299 9842 7331
rect 9714 7291 9755 7299
rect 9531 7191 9577 7253
rect 9531 7132 9577 7145
rect 9801 7291 9842 7299
rect 9979 7839 10025 7901
rect 10203 8164 10249 8227
rect 10203 8055 10249 8118
rect 10203 7947 10249 8009
rect 10203 7858 10249 7901
rect 10427 8164 10473 8227
rect 10427 8055 10473 8118
rect 10427 7947 10473 8009
rect 9979 7731 10025 7793
rect 9979 7623 10025 7685
rect 9979 7515 10025 7577
rect 9979 7407 10025 7469
rect 9979 7299 10025 7361
rect 9755 7191 9801 7253
rect 9755 7132 9801 7145
rect 10162 7839 10290 7858
rect 10162 7819 10203 7839
rect 10249 7819 10290 7839
rect 10162 7767 10200 7819
rect 10252 7767 10290 7819
rect 10162 7731 10290 7767
rect 10162 7685 10203 7731
rect 10249 7685 10290 7731
rect 10162 7623 10290 7685
rect 10162 7601 10203 7623
rect 10249 7601 10290 7623
rect 10162 7549 10200 7601
rect 10252 7549 10290 7601
rect 10162 7515 10290 7549
rect 10162 7469 10203 7515
rect 10249 7469 10290 7515
rect 10162 7407 10290 7469
rect 10162 7383 10203 7407
rect 10249 7383 10290 7407
rect 10162 7331 10200 7383
rect 10252 7331 10290 7383
rect 10162 7299 10290 7331
rect 10162 7291 10203 7299
rect 9979 7191 10025 7253
rect 9979 7132 10025 7145
rect 10249 7291 10290 7299
rect 10427 7839 10473 7901
rect 10427 7731 10473 7793
rect 10427 7623 10473 7685
rect 10427 7515 10473 7577
rect 10427 7407 10473 7469
rect 10427 7299 10473 7361
rect 10203 7191 10249 7253
rect 10203 7132 10249 7145
rect 10427 7191 10473 7253
rect 10427 7132 10473 7145
rect 10717 8164 10763 8227
rect 10717 8055 10763 8118
rect 10717 7947 10763 8009
rect 10717 7839 10763 7901
rect 10941 8164 10987 8227
rect 10941 8055 10987 8118
rect 10941 7947 10987 8009
rect 10941 7858 10987 7901
rect 11165 8164 11211 8227
rect 11165 8055 11211 8118
rect 11165 7947 11211 8009
rect 10717 7731 10763 7793
rect 10717 7623 10763 7685
rect 10717 7515 10763 7577
rect 10717 7407 10763 7469
rect 10717 7299 10763 7361
rect 10900 7839 11028 7858
rect 10900 7819 10941 7839
rect 10987 7819 11028 7839
rect 10900 7767 10938 7819
rect 10990 7767 11028 7819
rect 10900 7731 11028 7767
rect 10900 7685 10941 7731
rect 10987 7685 11028 7731
rect 10900 7623 11028 7685
rect 10900 7601 10941 7623
rect 10987 7601 11028 7623
rect 10900 7549 10938 7601
rect 10990 7549 11028 7601
rect 10900 7515 11028 7549
rect 10900 7469 10941 7515
rect 10987 7469 11028 7515
rect 10900 7407 11028 7469
rect 10900 7383 10941 7407
rect 10987 7383 11028 7407
rect 10900 7331 10938 7383
rect 10990 7331 11028 7383
rect 10900 7299 11028 7331
rect 10900 7291 10941 7299
rect 10717 7191 10763 7253
rect 10717 7132 10763 7145
rect 10987 7291 11028 7299
rect 11165 7839 11211 7901
rect 11389 8164 11435 8227
rect 11389 8055 11435 8118
rect 11389 7947 11435 8009
rect 11389 7858 11435 7901
rect 11613 8164 11659 8227
rect 11613 8055 11659 8118
rect 11613 7947 11659 8009
rect 11165 7731 11211 7793
rect 11165 7623 11211 7685
rect 11165 7515 11211 7577
rect 11165 7407 11211 7469
rect 11165 7299 11211 7361
rect 10941 7191 10987 7253
rect 10941 7132 10987 7145
rect 11348 7839 11476 7858
rect 11348 7819 11389 7839
rect 11435 7819 11476 7839
rect 11348 7767 11386 7819
rect 11438 7767 11476 7819
rect 11348 7731 11476 7767
rect 11348 7685 11389 7731
rect 11435 7685 11476 7731
rect 11348 7623 11476 7685
rect 11348 7601 11389 7623
rect 11435 7601 11476 7623
rect 11348 7549 11386 7601
rect 11438 7549 11476 7601
rect 11348 7515 11476 7549
rect 11348 7469 11389 7515
rect 11435 7469 11476 7515
rect 11348 7407 11476 7469
rect 11348 7383 11389 7407
rect 11435 7383 11476 7407
rect 11348 7331 11386 7383
rect 11438 7331 11476 7383
rect 11348 7299 11476 7331
rect 11348 7291 11389 7299
rect 11165 7191 11211 7253
rect 11165 7132 11211 7145
rect 11435 7291 11476 7299
rect 11613 7839 11659 7901
rect 11837 8164 11883 8227
rect 11837 8055 11883 8118
rect 11837 7947 11883 8009
rect 11837 7858 11883 7901
rect 12061 8164 12107 8227
rect 12061 8055 12107 8118
rect 12061 7947 12107 8009
rect 11613 7731 11659 7793
rect 11613 7623 11659 7685
rect 11613 7515 11659 7577
rect 11613 7407 11659 7469
rect 11613 7299 11659 7361
rect 11389 7191 11435 7253
rect 11389 7132 11435 7145
rect 11796 7839 11924 7858
rect 11796 7819 11837 7839
rect 11883 7819 11924 7839
rect 11796 7767 11834 7819
rect 11886 7767 11924 7819
rect 11796 7731 11924 7767
rect 11796 7685 11837 7731
rect 11883 7685 11924 7731
rect 11796 7623 11924 7685
rect 11796 7601 11837 7623
rect 11883 7601 11924 7623
rect 11796 7549 11834 7601
rect 11886 7549 11924 7601
rect 11796 7515 11924 7549
rect 11796 7469 11837 7515
rect 11883 7469 11924 7515
rect 11796 7407 11924 7469
rect 11796 7383 11837 7407
rect 11883 7383 11924 7407
rect 11796 7331 11834 7383
rect 11886 7331 11924 7383
rect 11796 7299 11924 7331
rect 11796 7291 11837 7299
rect 11613 7191 11659 7253
rect 11613 7132 11659 7145
rect 11883 7291 11924 7299
rect 12061 7839 12107 7901
rect 12061 7731 12107 7793
rect 12061 7623 12107 7685
rect 12061 7515 12107 7577
rect 12061 7407 12107 7469
rect 12061 7299 12107 7361
rect 11837 7191 11883 7253
rect 11837 7132 11883 7145
rect 12061 7191 12107 7253
rect 12061 7132 12107 7145
rect 12351 8164 12397 8227
rect 12351 8055 12397 8118
rect 12351 7947 12397 8009
rect 12351 7839 12397 7901
rect 12575 8164 12621 8227
rect 12575 8055 12621 8118
rect 12575 7947 12621 8009
rect 12575 7858 12621 7901
rect 12799 8164 12845 8227
rect 12799 8055 12845 8118
rect 12799 7947 12845 8009
rect 12351 7731 12397 7793
rect 12351 7623 12397 7685
rect 12351 7515 12397 7577
rect 12351 7407 12397 7469
rect 12351 7299 12397 7361
rect 12534 7839 12662 7858
rect 12534 7819 12575 7839
rect 12621 7819 12662 7839
rect 12534 7767 12572 7819
rect 12624 7767 12662 7819
rect 12534 7731 12662 7767
rect 12534 7685 12575 7731
rect 12621 7685 12662 7731
rect 12534 7623 12662 7685
rect 12534 7601 12575 7623
rect 12621 7601 12662 7623
rect 12534 7549 12572 7601
rect 12624 7549 12662 7601
rect 12534 7515 12662 7549
rect 12534 7469 12575 7515
rect 12621 7469 12662 7515
rect 12534 7407 12662 7469
rect 12534 7383 12575 7407
rect 12621 7383 12662 7407
rect 12534 7331 12572 7383
rect 12624 7331 12662 7383
rect 12534 7299 12662 7331
rect 12534 7291 12575 7299
rect 12351 7191 12397 7253
rect 12351 7132 12397 7145
rect 12621 7291 12662 7299
rect 12799 7839 12845 7901
rect 13023 8164 13069 8227
rect 13023 8055 13069 8118
rect 13023 7947 13069 8009
rect 13023 7858 13069 7901
rect 13247 8164 13293 8227
rect 13247 8055 13293 8118
rect 13247 7947 13293 8009
rect 12799 7731 12845 7793
rect 12799 7623 12845 7685
rect 12799 7515 12845 7577
rect 12799 7407 12845 7469
rect 12799 7299 12845 7361
rect 12575 7191 12621 7253
rect 12575 7132 12621 7145
rect 12982 7839 13110 7858
rect 12982 7819 13023 7839
rect 13069 7819 13110 7839
rect 12982 7767 13020 7819
rect 13072 7767 13110 7819
rect 12982 7731 13110 7767
rect 12982 7685 13023 7731
rect 13069 7685 13110 7731
rect 12982 7623 13110 7685
rect 12982 7601 13023 7623
rect 13069 7601 13110 7623
rect 12982 7549 13020 7601
rect 13072 7549 13110 7601
rect 12982 7515 13110 7549
rect 12982 7469 13023 7515
rect 13069 7469 13110 7515
rect 12982 7407 13110 7469
rect 12982 7383 13023 7407
rect 13069 7383 13110 7407
rect 12982 7331 13020 7383
rect 13072 7331 13110 7383
rect 12982 7299 13110 7331
rect 12982 7291 13023 7299
rect 12799 7191 12845 7253
rect 12799 7132 12845 7145
rect 13069 7291 13110 7299
rect 13247 7839 13293 7901
rect 13471 8164 13517 8227
rect 13471 8055 13517 8118
rect 13471 7947 13517 8009
rect 13471 7858 13517 7901
rect 13695 8164 13741 8227
rect 13695 8055 13741 8118
rect 13695 7947 13741 8009
rect 13247 7731 13293 7793
rect 13247 7623 13293 7685
rect 13247 7515 13293 7577
rect 13247 7407 13293 7469
rect 13247 7299 13293 7361
rect 13023 7191 13069 7253
rect 13023 7132 13069 7145
rect 13430 7839 13558 7858
rect 13430 7819 13471 7839
rect 13517 7819 13558 7839
rect 13430 7767 13468 7819
rect 13520 7767 13558 7819
rect 13430 7731 13558 7767
rect 13430 7685 13471 7731
rect 13517 7685 13558 7731
rect 13430 7623 13558 7685
rect 13430 7601 13471 7623
rect 13517 7601 13558 7623
rect 13430 7549 13468 7601
rect 13520 7549 13558 7601
rect 13430 7515 13558 7549
rect 13430 7469 13471 7515
rect 13517 7469 13558 7515
rect 13430 7407 13558 7469
rect 13430 7383 13471 7407
rect 13517 7383 13558 7407
rect 13430 7331 13468 7383
rect 13520 7331 13558 7383
rect 13430 7299 13558 7331
rect 13430 7291 13471 7299
rect 13247 7191 13293 7253
rect 13247 7132 13293 7145
rect 13517 7291 13558 7299
rect 13695 7839 13741 7901
rect 13695 7731 13741 7793
rect 13695 7623 13741 7685
rect 13695 7515 13741 7577
rect 13695 7407 13741 7469
rect 13695 7299 13741 7361
rect 13471 7191 13517 7253
rect 13471 7132 13517 7145
rect 13695 7191 13741 7253
rect 13695 7132 13741 7145
rect 7416 7044 8090 7081
rect 7416 6998 7678 7044
rect 7912 6998 8090 7044
rect 7416 6962 8090 6998
rect 8200 7044 8874 7081
rect 8200 6998 8378 7044
rect 8612 6998 8874 7044
rect 8200 6962 8874 6998
rect 7416 6406 7531 6962
rect 7640 6808 8650 6845
rect 7640 6762 7727 6808
rect 7773 6762 7885 6808
rect 7931 6762 8043 6808
rect 8089 6762 8201 6808
rect 8247 6762 8359 6808
rect 8405 6762 8517 6808
rect 8563 6762 8650 6808
rect 7640 6750 8650 6762
rect 7416 6386 7450 6406
rect 7496 6386 7531 6406
rect 7638 6726 8652 6750
rect 7638 6709 7765 6726
rect 7638 6657 7675 6709
rect 7727 6657 7765 6709
rect 7638 6492 7765 6657
rect 7638 6440 7675 6492
rect 7727 6440 7765 6492
rect 7638 6406 7765 6440
rect 8081 6710 8209 6726
rect 8081 6658 8119 6710
rect 8171 6658 8209 6710
rect 8081 6492 8209 6658
rect 8081 6440 8119 6492
rect 8171 6440 8209 6492
rect 7450 6300 7496 6360
rect 7450 6194 7496 6254
rect 7450 6088 7496 6148
rect 7450 5982 7496 6042
rect 7450 5876 7496 5936
rect 7450 5770 7496 5830
rect 7638 6360 7674 6406
rect 7720 6360 7765 6406
rect 7638 6300 7765 6360
rect 7638 6254 7674 6300
rect 7720 6274 7765 6300
rect 7638 6222 7675 6254
rect 7727 6222 7765 6274
rect 7638 6194 7765 6222
rect 7638 6148 7674 6194
rect 7720 6148 7765 6194
rect 7638 6088 7765 6148
rect 7638 6042 7674 6088
rect 7720 6056 7765 6088
rect 7638 6004 7675 6042
rect 7727 6004 7765 6056
rect 7638 5982 7765 6004
rect 7638 5936 7674 5982
rect 7720 5936 7765 5982
rect 7638 5876 7765 5936
rect 7638 5830 7674 5876
rect 7720 5839 7765 5876
rect 7638 5787 7675 5830
rect 7727 5787 7765 5839
rect 7638 5770 7765 5787
rect 7638 5746 7674 5770
rect 7450 5664 7496 5724
rect 7411 5618 7450 5644
rect 7720 5746 7765 5770
rect 7898 6406 7944 6419
rect 7898 6300 7944 6360
rect 7898 6194 7944 6254
rect 7898 6088 7944 6148
rect 7898 5982 7944 6042
rect 7898 5876 7944 5936
rect 7898 5770 7944 5830
rect 7674 5664 7720 5724
rect 7496 5618 7535 5644
rect 6787 5574 6825 5614
rect 6701 5522 6737 5574
rect 6789 5522 6825 5574
rect 6701 5356 6741 5522
rect 6787 5356 6825 5522
rect 6701 5304 6737 5356
rect 6789 5304 6825 5356
rect 6701 5268 6741 5304
rect 6787 5268 6825 5304
rect 7411 5604 7535 5618
rect 7411 5552 7447 5604
rect 7499 5552 7535 5604
rect 7411 5512 7450 5552
rect 7496 5512 7535 5552
rect 7411 5451 7535 5512
rect 7411 5405 7450 5451
rect 7496 5405 7535 5451
rect 7411 5386 7535 5405
rect 7411 5334 7447 5386
rect 7499 5334 7535 5386
rect 7411 5298 7450 5334
rect 7496 5298 7535 5334
rect 7411 5294 7535 5298
rect 7898 5664 7944 5724
rect 7674 5558 7720 5618
rect 7674 5451 7720 5512
rect 7674 5344 7720 5405
rect 7450 5285 7496 5294
rect 7674 5285 7720 5298
rect 7859 5618 7898 5644
rect 8081 6406 8209 6440
rect 8525 6709 8652 6726
rect 8525 6657 8563 6709
rect 8615 6657 8652 6709
rect 8525 6492 8652 6657
rect 8525 6440 8563 6492
rect 8615 6440 8652 6492
rect 8081 6360 8122 6406
rect 8168 6360 8209 6406
rect 8081 6300 8209 6360
rect 8081 6275 8122 6300
rect 8168 6275 8209 6300
rect 8081 6223 8119 6275
rect 8171 6223 8209 6275
rect 8081 6194 8209 6223
rect 8081 6148 8122 6194
rect 8168 6148 8209 6194
rect 8081 6088 8209 6148
rect 8081 6057 8122 6088
rect 8168 6057 8209 6088
rect 8081 6005 8119 6057
rect 8171 6005 8209 6057
rect 8081 5982 8209 6005
rect 8081 5936 8122 5982
rect 8168 5936 8209 5982
rect 8081 5876 8209 5936
rect 8081 5839 8122 5876
rect 8168 5839 8209 5876
rect 8081 5787 8119 5839
rect 8171 5787 8209 5839
rect 8081 5770 8209 5787
rect 8081 5724 8122 5770
rect 8168 5724 8209 5770
rect 8081 5664 8209 5724
rect 7944 5618 7983 5644
rect 7859 5604 7983 5618
rect 7859 5552 7895 5604
rect 7947 5552 7983 5604
rect 7859 5512 7898 5552
rect 7944 5512 7983 5552
rect 7859 5451 7983 5512
rect 7859 5405 7898 5451
rect 7944 5405 7983 5451
rect 7859 5386 7983 5405
rect 7859 5334 7895 5386
rect 7947 5334 7983 5386
rect 7859 5298 7898 5334
rect 7944 5298 7983 5334
rect 8081 5622 8122 5664
rect 8168 5622 8209 5664
rect 8346 6406 8392 6419
rect 8346 6300 8392 6360
rect 8346 6194 8392 6254
rect 8346 6088 8392 6148
rect 8346 5982 8392 6042
rect 8346 5876 8392 5936
rect 8346 5770 8392 5830
rect 8525 6406 8652 6440
rect 8525 6360 8570 6406
rect 8616 6360 8652 6406
rect 8759 6406 8874 6962
rect 8759 6386 8794 6406
rect 8525 6300 8652 6360
rect 8525 6274 8570 6300
rect 8525 6222 8563 6274
rect 8616 6254 8652 6300
rect 8615 6222 8652 6254
rect 8525 6194 8652 6222
rect 8525 6148 8570 6194
rect 8616 6148 8652 6194
rect 8525 6088 8652 6148
rect 8525 6056 8570 6088
rect 8525 6004 8563 6056
rect 8616 6042 8652 6088
rect 8615 6004 8652 6042
rect 8525 5982 8652 6004
rect 8525 5936 8570 5982
rect 8616 5936 8652 5982
rect 8525 5876 8652 5936
rect 8525 5839 8570 5876
rect 8525 5787 8563 5839
rect 8616 5830 8652 5876
rect 8615 5787 8652 5830
rect 8525 5770 8652 5787
rect 8525 5746 8570 5770
rect 8346 5664 8392 5724
rect 8081 5570 8119 5622
rect 8171 5570 8209 5622
rect 8081 5558 8209 5570
rect 8081 5512 8122 5558
rect 8168 5512 8209 5558
rect 8081 5451 8209 5512
rect 8081 5405 8122 5451
rect 8168 5405 8209 5451
rect 8081 5404 8209 5405
rect 8081 5352 8119 5404
rect 8171 5352 8209 5404
rect 8081 5344 8209 5352
rect 8081 5311 8122 5344
rect 7859 5294 7983 5298
rect 8168 5311 8209 5344
rect 8307 5618 8346 5644
rect 8616 5746 8652 5770
rect 8840 6386 8874 6406
rect 9049 7044 9723 7081
rect 9049 6998 9311 7044
rect 9545 6998 9723 7044
rect 9049 6962 9723 6998
rect 9833 7044 10507 7081
rect 9833 6998 10011 7044
rect 10245 6998 10507 7044
rect 9833 6962 10507 6998
rect 9049 6406 9164 6962
rect 9273 6808 10283 6845
rect 9273 6762 9360 6808
rect 9406 6762 9518 6808
rect 9564 6762 9676 6808
rect 9722 6762 9834 6808
rect 9880 6762 9992 6808
rect 10038 6762 10150 6808
rect 10196 6762 10283 6808
rect 9273 6750 10283 6762
rect 9049 6386 9083 6406
rect 8794 6300 8840 6360
rect 8794 6194 8840 6254
rect 8794 6088 8840 6148
rect 8794 5982 8840 6042
rect 8794 5876 8840 5936
rect 8794 5770 8840 5830
rect 8570 5664 8616 5724
rect 8392 5618 8431 5644
rect 8307 5604 8431 5618
rect 8307 5552 8343 5604
rect 8395 5552 8431 5604
rect 8307 5512 8346 5552
rect 8392 5512 8431 5552
rect 8307 5451 8431 5512
rect 8307 5405 8346 5451
rect 8392 5405 8431 5451
rect 8307 5386 8431 5405
rect 8307 5334 8343 5386
rect 8395 5334 8431 5386
rect 7898 5285 7944 5294
rect 8122 5285 8168 5298
rect 8307 5298 8346 5334
rect 8392 5298 8431 5334
rect 8307 5294 8431 5298
rect 8794 5664 8840 5724
rect 8570 5558 8616 5618
rect 8570 5451 8616 5512
rect 8570 5344 8616 5405
rect 8346 5285 8392 5294
rect 8570 5285 8616 5298
rect 8755 5618 8794 5644
rect 9129 6386 9164 6406
rect 9271 6726 10285 6750
rect 9271 6709 9398 6726
rect 9271 6657 9308 6709
rect 9360 6657 9398 6709
rect 9271 6492 9398 6657
rect 9271 6440 9308 6492
rect 9360 6440 9398 6492
rect 9271 6406 9398 6440
rect 9714 6710 9842 6726
rect 9714 6658 9752 6710
rect 9804 6658 9842 6710
rect 9714 6492 9842 6658
rect 9714 6440 9752 6492
rect 9804 6440 9842 6492
rect 9083 6300 9129 6360
rect 9083 6194 9129 6254
rect 9083 6088 9129 6148
rect 9083 5982 9129 6042
rect 9083 5876 9129 5936
rect 9083 5770 9129 5830
rect 9271 6360 9307 6406
rect 9353 6360 9398 6406
rect 9271 6300 9398 6360
rect 9271 6254 9307 6300
rect 9353 6274 9398 6300
rect 9271 6222 9308 6254
rect 9360 6222 9398 6274
rect 9271 6194 9398 6222
rect 9271 6148 9307 6194
rect 9353 6148 9398 6194
rect 9271 6088 9398 6148
rect 9271 6042 9307 6088
rect 9353 6056 9398 6088
rect 9271 6004 9308 6042
rect 9360 6004 9398 6056
rect 9271 5982 9398 6004
rect 9271 5936 9307 5982
rect 9353 5936 9398 5982
rect 9271 5876 9398 5936
rect 9271 5830 9307 5876
rect 9353 5839 9398 5876
rect 9271 5787 9308 5830
rect 9360 5787 9398 5839
rect 9271 5770 9398 5787
rect 9271 5746 9307 5770
rect 9083 5664 9129 5724
rect 8840 5618 8879 5644
rect 8755 5604 8879 5618
rect 8755 5552 8791 5604
rect 8843 5552 8879 5604
rect 8755 5512 8794 5552
rect 8840 5512 8879 5552
rect 8755 5451 8879 5512
rect 8755 5405 8794 5451
rect 8840 5405 8879 5451
rect 8755 5386 8879 5405
rect 8755 5334 8791 5386
rect 8843 5334 8879 5386
rect 8755 5298 8794 5334
rect 8840 5298 8879 5334
rect 8755 5294 8879 5298
rect 9044 5618 9083 5644
rect 9353 5746 9398 5770
rect 9531 6406 9577 6419
rect 9531 6300 9577 6360
rect 9531 6194 9577 6254
rect 9531 6088 9577 6148
rect 9531 5982 9577 6042
rect 9531 5876 9577 5936
rect 9531 5770 9577 5830
rect 9307 5664 9353 5724
rect 9129 5618 9168 5644
rect 9044 5604 9168 5618
rect 9044 5552 9080 5604
rect 9132 5552 9168 5604
rect 9044 5512 9083 5552
rect 9129 5512 9168 5552
rect 9044 5451 9168 5512
rect 9044 5405 9083 5451
rect 9129 5405 9168 5451
rect 9044 5386 9168 5405
rect 9044 5334 9080 5386
rect 9132 5334 9168 5386
rect 9044 5298 9083 5334
rect 9129 5298 9168 5334
rect 9044 5294 9168 5298
rect 9531 5664 9577 5724
rect 9307 5558 9353 5618
rect 9307 5451 9353 5512
rect 9307 5344 9353 5405
rect 8794 5285 8840 5294
rect 9083 5285 9129 5294
rect 9307 5285 9353 5298
rect 9492 5618 9531 5644
rect 9714 6406 9842 6440
rect 10158 6709 10285 6726
rect 10158 6657 10196 6709
rect 10248 6657 10285 6709
rect 10158 6492 10285 6657
rect 10158 6440 10196 6492
rect 10248 6440 10285 6492
rect 9714 6360 9755 6406
rect 9801 6360 9842 6406
rect 9714 6300 9842 6360
rect 9714 6275 9755 6300
rect 9801 6275 9842 6300
rect 9714 6223 9752 6275
rect 9804 6223 9842 6275
rect 9714 6194 9842 6223
rect 9714 6148 9755 6194
rect 9801 6148 9842 6194
rect 9714 6088 9842 6148
rect 9714 6057 9755 6088
rect 9801 6057 9842 6088
rect 9714 6005 9752 6057
rect 9804 6005 9842 6057
rect 9714 5982 9842 6005
rect 9714 5936 9755 5982
rect 9801 5936 9842 5982
rect 9714 5876 9842 5936
rect 9714 5839 9755 5876
rect 9801 5839 9842 5876
rect 9714 5787 9752 5839
rect 9804 5787 9842 5839
rect 9714 5770 9842 5787
rect 9714 5724 9755 5770
rect 9801 5724 9842 5770
rect 9714 5664 9842 5724
rect 9577 5618 9616 5644
rect 9492 5604 9616 5618
rect 9492 5552 9528 5604
rect 9580 5552 9616 5604
rect 9492 5512 9531 5552
rect 9577 5512 9616 5552
rect 9492 5451 9616 5512
rect 9492 5405 9531 5451
rect 9577 5405 9616 5451
rect 9492 5386 9616 5405
rect 9492 5334 9528 5386
rect 9580 5334 9616 5386
rect 9492 5298 9531 5334
rect 9577 5298 9616 5334
rect 9714 5622 9755 5664
rect 9801 5622 9842 5664
rect 9979 6406 10025 6419
rect 9979 6300 10025 6360
rect 9979 6194 10025 6254
rect 9979 6088 10025 6148
rect 9979 5982 10025 6042
rect 9979 5876 10025 5936
rect 9979 5770 10025 5830
rect 10158 6406 10285 6440
rect 10158 6360 10203 6406
rect 10249 6360 10285 6406
rect 10392 6406 10507 6962
rect 10392 6386 10427 6406
rect 10158 6300 10285 6360
rect 10158 6274 10203 6300
rect 10158 6222 10196 6274
rect 10249 6254 10285 6300
rect 10248 6222 10285 6254
rect 10158 6194 10285 6222
rect 10158 6148 10203 6194
rect 10249 6148 10285 6194
rect 10158 6088 10285 6148
rect 10158 6056 10203 6088
rect 10158 6004 10196 6056
rect 10249 6042 10285 6088
rect 10248 6004 10285 6042
rect 10158 5982 10285 6004
rect 10158 5936 10203 5982
rect 10249 5936 10285 5982
rect 10158 5876 10285 5936
rect 10158 5839 10203 5876
rect 10158 5787 10196 5839
rect 10249 5830 10285 5876
rect 10248 5787 10285 5830
rect 10158 5770 10285 5787
rect 10158 5746 10203 5770
rect 9979 5664 10025 5724
rect 9714 5570 9752 5622
rect 9804 5570 9842 5622
rect 9714 5558 9842 5570
rect 9714 5512 9755 5558
rect 9801 5512 9842 5558
rect 9714 5451 9842 5512
rect 9714 5405 9755 5451
rect 9801 5405 9842 5451
rect 9714 5404 9842 5405
rect 9714 5352 9752 5404
rect 9804 5352 9842 5404
rect 9714 5344 9842 5352
rect 9714 5311 9755 5344
rect 9492 5294 9616 5298
rect 9801 5311 9842 5344
rect 9940 5618 9979 5644
rect 10249 5746 10285 5770
rect 10473 6386 10507 6406
rect 10683 7044 11357 7081
rect 10683 6998 10945 7044
rect 11179 6998 11357 7044
rect 10683 6962 11357 6998
rect 11467 7044 12141 7081
rect 11467 6998 11645 7044
rect 11879 6998 12141 7044
rect 11467 6962 12141 6998
rect 10683 6406 10798 6962
rect 10907 6808 11917 6845
rect 10907 6762 10994 6808
rect 11040 6762 11152 6808
rect 11198 6762 11310 6808
rect 11356 6762 11468 6808
rect 11514 6762 11626 6808
rect 11672 6762 11784 6808
rect 11830 6762 11917 6808
rect 10907 6750 11917 6762
rect 10683 6386 10717 6406
rect 10427 6300 10473 6360
rect 10427 6194 10473 6254
rect 10427 6088 10473 6148
rect 10427 5982 10473 6042
rect 10427 5876 10473 5936
rect 10427 5770 10473 5830
rect 10203 5664 10249 5724
rect 10025 5618 10064 5644
rect 9940 5604 10064 5618
rect 9940 5552 9976 5604
rect 10028 5552 10064 5604
rect 9940 5512 9979 5552
rect 10025 5512 10064 5552
rect 9940 5451 10064 5512
rect 9940 5405 9979 5451
rect 10025 5405 10064 5451
rect 9940 5386 10064 5405
rect 9940 5334 9976 5386
rect 10028 5334 10064 5386
rect 9531 5285 9577 5294
rect 9755 5285 9801 5298
rect 9940 5298 9979 5334
rect 10025 5298 10064 5334
rect 9940 5294 10064 5298
rect 10427 5664 10473 5724
rect 10203 5558 10249 5618
rect 10203 5451 10249 5512
rect 10203 5344 10249 5405
rect 9979 5285 10025 5294
rect 10203 5285 10249 5298
rect 10388 5618 10427 5644
rect 10763 6386 10798 6406
rect 10905 6726 11919 6750
rect 10905 6709 11032 6726
rect 10905 6657 10942 6709
rect 10994 6657 11032 6709
rect 10905 6492 11032 6657
rect 10905 6440 10942 6492
rect 10994 6440 11032 6492
rect 10905 6406 11032 6440
rect 11348 6710 11476 6726
rect 11348 6658 11386 6710
rect 11438 6658 11476 6710
rect 11348 6492 11476 6658
rect 11348 6440 11386 6492
rect 11438 6440 11476 6492
rect 10717 6300 10763 6360
rect 10717 6194 10763 6254
rect 10717 6088 10763 6148
rect 10717 5982 10763 6042
rect 10717 5876 10763 5936
rect 10717 5770 10763 5830
rect 10905 6360 10941 6406
rect 10987 6360 11032 6406
rect 10905 6300 11032 6360
rect 10905 6254 10941 6300
rect 10987 6274 11032 6300
rect 10905 6222 10942 6254
rect 10994 6222 11032 6274
rect 10905 6194 11032 6222
rect 10905 6148 10941 6194
rect 10987 6148 11032 6194
rect 10905 6088 11032 6148
rect 10905 6042 10941 6088
rect 10987 6056 11032 6088
rect 10905 6004 10942 6042
rect 10994 6004 11032 6056
rect 10905 5982 11032 6004
rect 10905 5936 10941 5982
rect 10987 5936 11032 5982
rect 10905 5876 11032 5936
rect 10905 5830 10941 5876
rect 10987 5839 11032 5876
rect 10905 5787 10942 5830
rect 10994 5787 11032 5839
rect 10905 5770 11032 5787
rect 10905 5746 10941 5770
rect 10717 5664 10763 5724
rect 10473 5618 10512 5644
rect 10388 5604 10512 5618
rect 10388 5552 10424 5604
rect 10476 5552 10512 5604
rect 10388 5512 10427 5552
rect 10473 5512 10512 5552
rect 10388 5451 10512 5512
rect 10388 5405 10427 5451
rect 10473 5405 10512 5451
rect 10388 5386 10512 5405
rect 10388 5334 10424 5386
rect 10476 5334 10512 5386
rect 10388 5298 10427 5334
rect 10473 5298 10512 5334
rect 10388 5294 10512 5298
rect 10678 5618 10717 5644
rect 10987 5746 11032 5770
rect 11165 6406 11211 6419
rect 11165 6300 11211 6360
rect 11165 6194 11211 6254
rect 11165 6088 11211 6148
rect 11165 5982 11211 6042
rect 11165 5876 11211 5936
rect 11165 5770 11211 5830
rect 10941 5664 10987 5724
rect 10763 5618 10802 5644
rect 10678 5604 10802 5618
rect 10678 5552 10714 5604
rect 10766 5552 10802 5604
rect 10678 5512 10717 5552
rect 10763 5512 10802 5552
rect 10678 5451 10802 5512
rect 10678 5405 10717 5451
rect 10763 5405 10802 5451
rect 10678 5386 10802 5405
rect 10678 5334 10714 5386
rect 10766 5334 10802 5386
rect 10678 5298 10717 5334
rect 10763 5298 10802 5334
rect 10678 5294 10802 5298
rect 11165 5664 11211 5724
rect 10941 5558 10987 5618
rect 10941 5451 10987 5512
rect 10941 5344 10987 5405
rect 10427 5285 10473 5294
rect 10717 5285 10763 5294
rect 10941 5285 10987 5298
rect 11126 5618 11165 5644
rect 11348 6406 11476 6440
rect 11792 6709 11919 6726
rect 11792 6657 11830 6709
rect 11882 6657 11919 6709
rect 11792 6492 11919 6657
rect 11792 6440 11830 6492
rect 11882 6440 11919 6492
rect 11348 6360 11389 6406
rect 11435 6360 11476 6406
rect 11348 6300 11476 6360
rect 11348 6275 11389 6300
rect 11435 6275 11476 6300
rect 11348 6223 11386 6275
rect 11438 6223 11476 6275
rect 11348 6194 11476 6223
rect 11348 6148 11389 6194
rect 11435 6148 11476 6194
rect 11348 6088 11476 6148
rect 11348 6057 11389 6088
rect 11435 6057 11476 6088
rect 11348 6005 11386 6057
rect 11438 6005 11476 6057
rect 11348 5982 11476 6005
rect 11348 5936 11389 5982
rect 11435 5936 11476 5982
rect 11348 5876 11476 5936
rect 11348 5839 11389 5876
rect 11435 5839 11476 5876
rect 11348 5787 11386 5839
rect 11438 5787 11476 5839
rect 11348 5770 11476 5787
rect 11348 5724 11389 5770
rect 11435 5724 11476 5770
rect 11348 5664 11476 5724
rect 11211 5618 11250 5644
rect 11126 5604 11250 5618
rect 11126 5552 11162 5604
rect 11214 5552 11250 5604
rect 11126 5512 11165 5552
rect 11211 5512 11250 5552
rect 11126 5451 11250 5512
rect 11126 5405 11165 5451
rect 11211 5405 11250 5451
rect 11126 5386 11250 5405
rect 11126 5334 11162 5386
rect 11214 5334 11250 5386
rect 11126 5298 11165 5334
rect 11211 5298 11250 5334
rect 11348 5622 11389 5664
rect 11435 5622 11476 5664
rect 11613 6406 11659 6419
rect 11613 6300 11659 6360
rect 11613 6194 11659 6254
rect 11613 6088 11659 6148
rect 11613 5982 11659 6042
rect 11613 5876 11659 5936
rect 11613 5770 11659 5830
rect 11792 6406 11919 6440
rect 11792 6360 11837 6406
rect 11883 6360 11919 6406
rect 12026 6406 12141 6962
rect 12026 6386 12061 6406
rect 11792 6300 11919 6360
rect 11792 6274 11837 6300
rect 11792 6222 11830 6274
rect 11883 6254 11919 6300
rect 11882 6222 11919 6254
rect 11792 6194 11919 6222
rect 11792 6148 11837 6194
rect 11883 6148 11919 6194
rect 11792 6088 11919 6148
rect 11792 6056 11837 6088
rect 11792 6004 11830 6056
rect 11883 6042 11919 6088
rect 11882 6004 11919 6042
rect 11792 5982 11919 6004
rect 11792 5936 11837 5982
rect 11883 5936 11919 5982
rect 11792 5876 11919 5936
rect 11792 5839 11837 5876
rect 11792 5787 11830 5839
rect 11883 5830 11919 5876
rect 11882 5787 11919 5830
rect 11792 5770 11919 5787
rect 11792 5746 11837 5770
rect 11613 5664 11659 5724
rect 11348 5570 11386 5622
rect 11438 5570 11476 5622
rect 11348 5558 11476 5570
rect 11348 5512 11389 5558
rect 11435 5512 11476 5558
rect 11348 5451 11476 5512
rect 11348 5405 11389 5451
rect 11435 5405 11476 5451
rect 11348 5404 11476 5405
rect 11348 5352 11386 5404
rect 11438 5352 11476 5404
rect 11348 5344 11476 5352
rect 11348 5311 11389 5344
rect 11126 5294 11250 5298
rect 11435 5311 11476 5344
rect 11574 5618 11613 5644
rect 11883 5746 11919 5770
rect 12107 6386 12141 6406
rect 12317 7044 12991 7081
rect 12317 6998 12579 7044
rect 12813 6998 12991 7044
rect 12317 6962 12991 6998
rect 13101 7044 13775 7081
rect 13101 6998 13279 7044
rect 13513 6998 13775 7044
rect 13101 6962 13775 6998
rect 12317 6406 12432 6962
rect 12541 6808 13551 6845
rect 12541 6762 12628 6808
rect 12674 6762 12786 6808
rect 12832 6762 12944 6808
rect 12990 6762 13102 6808
rect 13148 6762 13260 6808
rect 13306 6762 13418 6808
rect 13464 6762 13551 6808
rect 12541 6750 13551 6762
rect 12317 6386 12351 6406
rect 12061 6300 12107 6360
rect 12061 6194 12107 6254
rect 12061 6088 12107 6148
rect 12061 5982 12107 6042
rect 12061 5876 12107 5936
rect 12061 5770 12107 5830
rect 11837 5664 11883 5724
rect 11659 5618 11698 5644
rect 11574 5604 11698 5618
rect 11574 5552 11610 5604
rect 11662 5552 11698 5604
rect 11574 5512 11613 5552
rect 11659 5512 11698 5552
rect 11574 5451 11698 5512
rect 11574 5405 11613 5451
rect 11659 5405 11698 5451
rect 11574 5386 11698 5405
rect 11574 5334 11610 5386
rect 11662 5334 11698 5386
rect 11165 5285 11211 5294
rect 11389 5285 11435 5298
rect 11574 5298 11613 5334
rect 11659 5298 11698 5334
rect 11574 5294 11698 5298
rect 12061 5664 12107 5724
rect 11837 5558 11883 5618
rect 11837 5451 11883 5512
rect 11837 5344 11883 5405
rect 11613 5285 11659 5294
rect 11837 5285 11883 5298
rect 12022 5618 12061 5644
rect 12397 6386 12432 6406
rect 12539 6726 13553 6750
rect 12539 6709 12666 6726
rect 12539 6657 12576 6709
rect 12628 6657 12666 6709
rect 12539 6492 12666 6657
rect 12539 6440 12576 6492
rect 12628 6440 12666 6492
rect 12539 6406 12666 6440
rect 12982 6710 13110 6726
rect 12982 6658 13020 6710
rect 13072 6658 13110 6710
rect 12982 6492 13110 6658
rect 12982 6440 13020 6492
rect 13072 6440 13110 6492
rect 12351 6300 12397 6360
rect 12351 6194 12397 6254
rect 12351 6088 12397 6148
rect 12351 5982 12397 6042
rect 12351 5876 12397 5936
rect 12351 5770 12397 5830
rect 12539 6360 12575 6406
rect 12621 6360 12666 6406
rect 12539 6300 12666 6360
rect 12539 6254 12575 6300
rect 12621 6274 12666 6300
rect 12539 6222 12576 6254
rect 12628 6222 12666 6274
rect 12539 6194 12666 6222
rect 12539 6148 12575 6194
rect 12621 6148 12666 6194
rect 12539 6088 12666 6148
rect 12539 6042 12575 6088
rect 12621 6056 12666 6088
rect 12539 6004 12576 6042
rect 12628 6004 12666 6056
rect 12539 5982 12666 6004
rect 12539 5936 12575 5982
rect 12621 5936 12666 5982
rect 12539 5876 12666 5936
rect 12539 5830 12575 5876
rect 12621 5839 12666 5876
rect 12539 5787 12576 5830
rect 12628 5787 12666 5839
rect 12539 5770 12666 5787
rect 12539 5746 12575 5770
rect 12351 5664 12397 5724
rect 12107 5618 12146 5644
rect 12022 5604 12146 5618
rect 12022 5552 12058 5604
rect 12110 5552 12146 5604
rect 12022 5512 12061 5552
rect 12107 5512 12146 5552
rect 12022 5451 12146 5512
rect 12022 5405 12061 5451
rect 12107 5405 12146 5451
rect 12022 5386 12146 5405
rect 12022 5334 12058 5386
rect 12110 5334 12146 5386
rect 12022 5298 12061 5334
rect 12107 5298 12146 5334
rect 12022 5294 12146 5298
rect 12312 5618 12351 5644
rect 12621 5746 12666 5770
rect 12799 6406 12845 6419
rect 12799 6300 12845 6360
rect 12799 6194 12845 6254
rect 12799 6088 12845 6148
rect 12799 5982 12845 6042
rect 12799 5876 12845 5936
rect 12799 5770 12845 5830
rect 12575 5664 12621 5724
rect 12397 5618 12436 5644
rect 12312 5604 12436 5618
rect 12312 5552 12348 5604
rect 12400 5552 12436 5604
rect 12312 5512 12351 5552
rect 12397 5512 12436 5552
rect 12312 5451 12436 5512
rect 12312 5405 12351 5451
rect 12397 5405 12436 5451
rect 12312 5386 12436 5405
rect 12312 5334 12348 5386
rect 12400 5334 12436 5386
rect 12312 5298 12351 5334
rect 12397 5298 12436 5334
rect 12312 5294 12436 5298
rect 12799 5664 12845 5724
rect 12575 5558 12621 5618
rect 12575 5451 12621 5512
rect 12575 5344 12621 5405
rect 12061 5285 12107 5294
rect 12351 5285 12397 5294
rect 12575 5285 12621 5298
rect 12760 5618 12799 5644
rect 12982 6406 13110 6440
rect 13426 6709 13553 6726
rect 13426 6657 13464 6709
rect 13516 6657 13553 6709
rect 13426 6492 13553 6657
rect 13426 6440 13464 6492
rect 13516 6440 13553 6492
rect 12982 6360 13023 6406
rect 13069 6360 13110 6406
rect 12982 6300 13110 6360
rect 12982 6275 13023 6300
rect 13069 6275 13110 6300
rect 12982 6223 13020 6275
rect 13072 6223 13110 6275
rect 12982 6194 13110 6223
rect 12982 6148 13023 6194
rect 13069 6148 13110 6194
rect 12982 6088 13110 6148
rect 12982 6057 13023 6088
rect 13069 6057 13110 6088
rect 12982 6005 13020 6057
rect 13072 6005 13110 6057
rect 12982 5982 13110 6005
rect 12982 5936 13023 5982
rect 13069 5936 13110 5982
rect 12982 5876 13110 5936
rect 12982 5839 13023 5876
rect 13069 5839 13110 5876
rect 12982 5787 13020 5839
rect 13072 5787 13110 5839
rect 12982 5770 13110 5787
rect 12982 5724 13023 5770
rect 13069 5724 13110 5770
rect 12982 5664 13110 5724
rect 12845 5618 12884 5644
rect 12760 5604 12884 5618
rect 12760 5552 12796 5604
rect 12848 5552 12884 5604
rect 12760 5512 12799 5552
rect 12845 5512 12884 5552
rect 12760 5451 12884 5512
rect 12760 5405 12799 5451
rect 12845 5405 12884 5451
rect 12760 5386 12884 5405
rect 12760 5334 12796 5386
rect 12848 5334 12884 5386
rect 12760 5298 12799 5334
rect 12845 5298 12884 5334
rect 12982 5622 13023 5664
rect 13069 5622 13110 5664
rect 13247 6406 13293 6419
rect 13247 6300 13293 6360
rect 13247 6194 13293 6254
rect 13247 6088 13293 6148
rect 13247 5982 13293 6042
rect 13247 5876 13293 5936
rect 13247 5770 13293 5830
rect 13426 6406 13553 6440
rect 13426 6360 13471 6406
rect 13517 6360 13553 6406
rect 13660 6406 13775 6962
rect 13660 6386 13695 6406
rect 13426 6300 13553 6360
rect 13426 6274 13471 6300
rect 13426 6222 13464 6274
rect 13517 6254 13553 6300
rect 13516 6222 13553 6254
rect 13426 6194 13553 6222
rect 13426 6148 13471 6194
rect 13517 6148 13553 6194
rect 13426 6088 13553 6148
rect 13426 6056 13471 6088
rect 13426 6004 13464 6056
rect 13517 6042 13553 6088
rect 13516 6004 13553 6042
rect 13426 5982 13553 6004
rect 13426 5936 13471 5982
rect 13517 5936 13553 5982
rect 13426 5876 13553 5936
rect 13426 5839 13471 5876
rect 13426 5787 13464 5839
rect 13517 5830 13553 5876
rect 13516 5787 13553 5830
rect 13426 5770 13553 5787
rect 13426 5746 13471 5770
rect 13247 5664 13293 5724
rect 12982 5570 13020 5622
rect 13072 5570 13110 5622
rect 12982 5558 13110 5570
rect 12982 5512 13023 5558
rect 13069 5512 13110 5558
rect 12982 5451 13110 5512
rect 12982 5405 13023 5451
rect 13069 5405 13110 5451
rect 12982 5404 13110 5405
rect 12982 5352 13020 5404
rect 13072 5352 13110 5404
rect 12982 5344 13110 5352
rect 12982 5311 13023 5344
rect 12760 5294 12884 5298
rect 13069 5311 13110 5344
rect 13208 5618 13247 5644
rect 13517 5746 13553 5770
rect 13741 6386 13775 6406
rect 13695 6300 13741 6360
rect 13695 6194 13741 6254
rect 13695 6088 13741 6148
rect 13695 5982 13741 6042
rect 13695 5876 13741 5936
rect 13695 5770 13741 5830
rect 13471 5664 13517 5724
rect 13293 5618 13332 5644
rect 13208 5604 13332 5618
rect 13208 5552 13244 5604
rect 13296 5552 13332 5604
rect 13208 5512 13247 5552
rect 13293 5512 13332 5552
rect 13208 5451 13332 5512
rect 13208 5405 13247 5451
rect 13293 5405 13332 5451
rect 13208 5386 13332 5405
rect 13208 5334 13244 5386
rect 13296 5334 13332 5386
rect 12799 5285 12845 5294
rect 13023 5285 13069 5298
rect 13208 5298 13247 5334
rect 13293 5298 13332 5334
rect 13208 5294 13332 5298
rect 13695 5664 13741 5724
rect 13471 5558 13517 5618
rect 13471 5451 13517 5512
rect 13471 5344 13517 5405
rect 13247 5285 13293 5294
rect 13471 5285 13517 5298
rect 13656 5618 13695 5644
rect 13741 5618 13780 5644
rect 13656 5604 13780 5618
rect 13656 5552 13692 5604
rect 13744 5552 13780 5604
rect 13656 5512 13695 5552
rect 13741 5512 13780 5552
rect 13656 5451 13780 5512
rect 13656 5405 13695 5451
rect 13741 5405 13780 5451
rect 13656 5386 13780 5405
rect 13656 5334 13692 5386
rect 13744 5334 13780 5386
rect 13656 5298 13695 5334
rect 13741 5298 13780 5334
rect 13656 5294 13780 5298
rect 13695 5285 13741 5294
rect 6701 5264 6825 5268
rect 6741 5255 6787 5264
rect 7527 5161 7642 5173
rect 8647 5161 8762 5173
rect 9160 5161 9275 5173
rect 10280 5161 10395 5173
rect 1931 5137 13921 5161
rect 1931 5091 7562 5137
rect 7608 5091 8682 5137
rect 8728 5091 9195 5137
rect 9241 5091 10315 5137
rect 10361 5091 13921 5137
rect 1931 5069 13921 5091
rect 1931 5068 7280 5069
rect 7527 5054 7642 5069
rect 8647 5054 8762 5069
rect 9160 5054 9275 5069
rect 10280 5054 10395 5069
rect 4494 4959 4623 4980
rect 7751 4959 7866 4974
rect 8423 4959 8538 4974
rect 11018 4959 11133 4974
rect 11690 4959 11805 4974
rect 1931 4939 13921 4959
rect 1931 4887 4533 4939
rect 4585 4938 13921 4939
rect 4585 4892 7786 4938
rect 7832 4892 8458 4938
rect 8504 4892 11053 4938
rect 11099 4892 11725 4938
rect 11771 4892 13921 4938
rect 4585 4887 13921 4892
rect 1931 4867 13921 4887
rect 1931 4866 7280 4867
rect 4494 4846 4623 4866
rect 7751 4855 7866 4867
rect 8423 4855 8538 4867
rect 11018 4855 11133 4867
rect 11690 4855 11805 4867
rect 6184 4757 6313 4778
rect 7975 4757 8090 4770
rect 9608 4757 9723 4770
rect 11242 4757 11357 4770
rect 12876 4757 12991 4770
rect 1931 4737 13921 4757
rect 1931 4685 6223 4737
rect 6275 4734 13921 4737
rect 6275 4688 8010 4734
rect 8056 4688 9643 4734
rect 9689 4688 11277 4734
rect 11323 4688 12911 4734
rect 12957 4688 13921 4734
rect 6275 4685 13921 4688
rect 1931 4665 13921 4685
rect 6184 4644 6313 4665
rect 7975 4651 8090 4665
rect 9608 4651 9723 4665
rect 11242 4651 11357 4665
rect 12876 4651 12991 4665
rect 3316 4555 3445 4576
rect 10794 4555 10909 4568
rect 11914 4555 12029 4568
rect 12428 4555 12543 4568
rect 13548 4555 13663 4568
rect 1931 4535 13921 4555
rect 1931 4483 3355 4535
rect 3407 4532 13921 4535
rect 3407 4486 10829 4532
rect 10875 4486 11949 4532
rect 11995 4486 12463 4532
rect 12509 4486 13583 4532
rect 13629 4486 13921 4532
rect 3407 4483 13921 4486
rect 1931 4463 13921 4483
rect 3316 4442 3445 4463
rect 10794 4449 10909 4463
rect 11914 4449 12029 4463
rect 12428 4449 12543 4463
rect 13548 4449 13663 4463
rect 5007 4354 5136 4374
rect 9384 4354 9499 4366
rect 10056 4354 10171 4366
rect 12652 4354 12767 4366
rect 13324 4354 13439 4366
rect 1931 4333 13921 4354
rect 1931 4281 5046 4333
rect 5098 4330 13921 4333
rect 5098 4284 9419 4330
rect 9465 4284 10091 4330
rect 10137 4284 12687 4330
rect 12733 4284 13359 4330
rect 13405 4284 13921 4330
rect 5098 4281 13921 4284
rect 1931 4262 13921 4281
rect 1931 4261 7280 4262
rect 5007 4240 5136 4261
rect 9384 4247 9499 4262
rect 10056 4247 10171 4262
rect 12652 4247 12767 4262
rect 13324 4247 13439 4262
rect 6698 4152 6827 4173
rect 8199 4152 8314 4165
rect 9832 4152 9947 4165
rect 11466 4152 11581 4165
rect 13100 4152 13215 4165
rect 1931 4132 13921 4152
rect 1931 4080 6737 4132
rect 6789 4129 13921 4132
rect 6789 4083 8234 4129
rect 8280 4083 9867 4129
rect 9913 4083 11501 4129
rect 11547 4083 13135 4129
rect 13181 4083 13921 4129
rect 6789 4080 13921 4083
rect 1931 4060 13921 4080
rect 1931 4059 7280 4060
rect 6698 4039 6827 4059
rect 8199 4046 8314 4060
rect 9832 4046 9947 4060
rect 11466 4046 11581 4060
rect 13100 4046 13215 4060
rect 7416 3866 7531 3903
rect 7416 3820 7450 3866
rect 7496 3820 7531 3866
rect 7416 3753 7531 3820
rect 8088 3866 8202 3903
rect 8088 3820 8122 3866
rect 8168 3820 8202 3866
rect 8088 3807 8202 3820
rect 8759 3866 8874 3903
rect 8759 3820 8794 3866
rect 8840 3820 8874 3866
rect 7410 3712 7537 3753
rect 7410 3660 7447 3712
rect 7499 3660 7537 3712
rect 7410 3652 7450 3660
rect 7496 3652 7537 3660
rect 7410 3530 7537 3652
rect 7410 3495 7450 3530
rect 7496 3495 7537 3530
rect 7410 3443 7447 3495
rect 7499 3443 7537 3495
rect 7410 3363 7537 3443
rect 7410 3317 7450 3363
rect 7496 3317 7537 3363
rect 7410 3277 7537 3317
rect 2368 3211 2492 3251
rect 2368 3159 2404 3211
rect 2456 3159 2492 3211
rect 2368 2993 2492 3159
rect 2368 2941 2404 2993
rect 2456 2941 2492 2993
rect 2368 2901 2492 2941
rect 4059 3211 4183 3251
rect 4059 3159 4095 3211
rect 4147 3159 4183 3211
rect 4059 2993 4183 3159
rect 4059 2941 4095 2993
rect 4147 2941 4183 2993
rect 4059 2901 4183 2941
rect 5750 3211 5874 3251
rect 5750 3159 5786 3211
rect 5838 3159 5874 3211
rect 5750 2993 5874 3159
rect 5750 2941 5786 2993
rect 5838 2941 5874 2993
rect 5750 2901 5874 2941
rect 7410 3225 7447 3277
rect 7499 3225 7537 3277
rect 7410 3195 7537 3225
rect 7410 3149 7450 3195
rect 7496 3149 7537 3195
rect 7410 3059 7537 3149
rect 7410 3007 7447 3059
rect 7499 3007 7537 3059
rect 7410 2981 7450 3007
rect 7496 2981 7537 3007
rect 7410 2859 7537 2981
rect 7410 2842 7450 2859
rect 7496 2842 7537 2859
rect 7410 2790 7447 2842
rect 7499 2790 7537 2842
rect 7410 2749 7537 2790
rect 8087 3698 8203 3807
rect 8759 3753 8874 3820
rect 9049 3866 9164 3903
rect 9049 3820 9083 3866
rect 9129 3820 9164 3866
rect 9049 3753 9164 3820
rect 9721 3866 9835 3903
rect 9721 3820 9755 3866
rect 9801 3820 9835 3866
rect 9721 3807 9835 3820
rect 10392 3866 10507 3903
rect 10392 3820 10427 3866
rect 10473 3820 10507 3866
rect 8087 3652 8122 3698
rect 8168 3652 8203 3698
rect 8087 3584 8203 3652
rect 7416 2692 7531 2749
rect 1714 1117 1844 1158
rect 1714 1065 1753 1117
rect 1805 1065 1844 1117
rect 1714 899 1844 1065
rect 1714 847 1753 899
rect 1805 847 1844 899
rect 1714 807 1844 847
rect 1714 806 1843 807
rect 6960 756 7089 2678
rect 7416 2646 7450 2692
rect 7496 2646 7531 2692
rect 7416 2559 7531 2646
rect 8087 2596 8119 3584
rect 8171 2596 8203 3584
rect 8753 3712 8880 3753
rect 8753 3660 8791 3712
rect 8843 3660 8880 3712
rect 8753 3652 8794 3660
rect 8840 3652 8880 3660
rect 8753 3530 8880 3652
rect 8753 3495 8794 3530
rect 8840 3495 8880 3530
rect 8753 3443 8791 3495
rect 8843 3443 8880 3495
rect 8753 3363 8880 3443
rect 8753 3317 8794 3363
rect 8840 3317 8880 3363
rect 8753 3277 8880 3317
rect 8753 3225 8791 3277
rect 8843 3225 8880 3277
rect 8753 3195 8880 3225
rect 8753 3149 8794 3195
rect 8840 3149 8880 3195
rect 8753 3059 8880 3149
rect 8753 3007 8791 3059
rect 8843 3007 8880 3059
rect 8753 2981 8794 3007
rect 8840 2981 8880 3007
rect 8753 2859 8880 2981
rect 8753 2842 8794 2859
rect 8840 2842 8880 2859
rect 8753 2790 8791 2842
rect 8843 2790 8880 2842
rect 8753 2749 8880 2790
rect 9043 3712 9170 3753
rect 9043 3660 9080 3712
rect 9132 3660 9170 3712
rect 9043 3652 9083 3660
rect 9129 3652 9170 3660
rect 9043 3530 9170 3652
rect 9043 3495 9083 3530
rect 9129 3495 9170 3530
rect 9043 3443 9080 3495
rect 9132 3443 9170 3495
rect 9043 3363 9170 3443
rect 9043 3317 9083 3363
rect 9129 3317 9170 3363
rect 9043 3277 9170 3317
rect 9043 3225 9080 3277
rect 9132 3225 9170 3277
rect 9043 3195 9170 3225
rect 9043 3149 9083 3195
rect 9129 3149 9170 3195
rect 9043 3059 9170 3149
rect 9043 3007 9080 3059
rect 9132 3007 9170 3059
rect 9043 2981 9083 3007
rect 9129 2981 9170 3007
rect 9043 2859 9170 2981
rect 9043 2842 9083 2859
rect 9129 2842 9170 2859
rect 9043 2790 9080 2842
rect 9132 2790 9170 2842
rect 9043 2749 9170 2790
rect 9720 3698 9836 3807
rect 10392 3753 10507 3820
rect 10683 3866 10798 3903
rect 10683 3820 10717 3866
rect 10763 3820 10798 3866
rect 10683 3753 10798 3820
rect 11355 3866 11469 3903
rect 11355 3820 11389 3866
rect 11435 3820 11469 3866
rect 11355 3807 11469 3820
rect 12026 3866 12141 3903
rect 12026 3820 12061 3866
rect 12107 3820 12141 3866
rect 9720 3652 9755 3698
rect 9801 3652 9836 3698
rect 9720 3584 9836 3652
rect 8087 2470 8203 2596
rect 8759 2692 8874 2749
rect 8759 2646 8794 2692
rect 8840 2646 8874 2692
rect 8759 2559 8874 2646
rect 9049 2692 9164 2749
rect 9049 2646 9083 2692
rect 9129 2646 9164 2692
rect 9049 2559 9164 2646
rect 9720 2596 9753 3584
rect 9805 2596 9836 3584
rect 10386 3712 10513 3753
rect 10386 3660 10424 3712
rect 10476 3660 10513 3712
rect 10386 3652 10427 3660
rect 10473 3652 10513 3660
rect 10386 3530 10513 3652
rect 10386 3495 10427 3530
rect 10473 3495 10513 3530
rect 10386 3443 10424 3495
rect 10476 3443 10513 3495
rect 10386 3363 10513 3443
rect 10386 3317 10427 3363
rect 10473 3317 10513 3363
rect 10386 3277 10513 3317
rect 10386 3225 10424 3277
rect 10476 3225 10513 3277
rect 10386 3195 10513 3225
rect 10386 3149 10427 3195
rect 10473 3149 10513 3195
rect 10386 3059 10513 3149
rect 10386 3007 10424 3059
rect 10476 3007 10513 3059
rect 10386 2981 10427 3007
rect 10473 2981 10513 3007
rect 10386 2859 10513 2981
rect 10386 2842 10427 2859
rect 10473 2842 10513 2859
rect 10386 2790 10424 2842
rect 10476 2790 10513 2842
rect 10386 2749 10513 2790
rect 10677 3712 10804 3753
rect 10677 3660 10714 3712
rect 10766 3660 10804 3712
rect 10677 3652 10717 3660
rect 10763 3652 10804 3660
rect 10677 3530 10804 3652
rect 10677 3495 10717 3530
rect 10763 3495 10804 3530
rect 10677 3443 10714 3495
rect 10766 3443 10804 3495
rect 10677 3363 10804 3443
rect 10677 3317 10717 3363
rect 10763 3317 10804 3363
rect 10677 3277 10804 3317
rect 10677 3225 10714 3277
rect 10766 3225 10804 3277
rect 10677 3195 10804 3225
rect 10677 3149 10717 3195
rect 10763 3149 10804 3195
rect 10677 3059 10804 3149
rect 10677 3007 10714 3059
rect 10766 3007 10804 3059
rect 10677 2981 10717 3007
rect 10763 2981 10804 3007
rect 10677 2859 10804 2981
rect 10677 2842 10717 2859
rect 10763 2842 10804 2859
rect 10677 2790 10714 2842
rect 10766 2790 10804 2842
rect 10677 2749 10804 2790
rect 11354 3698 11470 3807
rect 12026 3753 12141 3820
rect 12317 3866 12432 3903
rect 12317 3820 12351 3866
rect 12397 3820 12432 3866
rect 12317 3753 12432 3820
rect 12989 3866 13103 3903
rect 12989 3820 13023 3866
rect 13069 3820 13103 3866
rect 12989 3807 13103 3820
rect 13660 3866 13775 3903
rect 13660 3820 13695 3866
rect 13741 3820 13775 3866
rect 11354 3652 11389 3698
rect 11435 3652 11470 3698
rect 11354 3584 11470 3652
rect 9720 2470 9836 2596
rect 10392 2692 10507 2749
rect 10392 2646 10427 2692
rect 10473 2646 10507 2692
rect 10392 2559 10507 2646
rect 10683 2692 10798 2749
rect 10683 2646 10717 2692
rect 10763 2646 10798 2692
rect 10683 2559 10798 2646
rect 11354 2596 11386 3584
rect 11438 2596 11470 3584
rect 12020 3712 12147 3753
rect 12020 3660 12058 3712
rect 12110 3660 12147 3712
rect 12020 3652 12061 3660
rect 12107 3652 12147 3660
rect 12020 3530 12147 3652
rect 12020 3495 12061 3530
rect 12107 3495 12147 3530
rect 12020 3443 12058 3495
rect 12110 3443 12147 3495
rect 12020 3363 12147 3443
rect 12020 3317 12061 3363
rect 12107 3317 12147 3363
rect 12020 3277 12147 3317
rect 12020 3225 12058 3277
rect 12110 3225 12147 3277
rect 12020 3195 12147 3225
rect 12020 3149 12061 3195
rect 12107 3149 12147 3195
rect 12020 3059 12147 3149
rect 12020 3007 12058 3059
rect 12110 3007 12147 3059
rect 12020 2981 12061 3007
rect 12107 2981 12147 3007
rect 12020 2859 12147 2981
rect 12020 2842 12061 2859
rect 12107 2842 12147 2859
rect 12020 2790 12058 2842
rect 12110 2790 12147 2842
rect 12020 2749 12147 2790
rect 12311 3712 12438 3753
rect 12311 3660 12348 3712
rect 12400 3660 12438 3712
rect 12311 3652 12351 3660
rect 12397 3652 12438 3660
rect 12311 3530 12438 3652
rect 12311 3495 12351 3530
rect 12397 3495 12438 3530
rect 12311 3443 12348 3495
rect 12400 3443 12438 3495
rect 12311 3363 12438 3443
rect 12311 3317 12351 3363
rect 12397 3317 12438 3363
rect 12311 3277 12438 3317
rect 12311 3225 12348 3277
rect 12400 3225 12438 3277
rect 12311 3195 12438 3225
rect 12311 3149 12351 3195
rect 12397 3149 12438 3195
rect 12311 3059 12438 3149
rect 12311 3007 12348 3059
rect 12400 3007 12438 3059
rect 12311 2981 12351 3007
rect 12397 2981 12438 3007
rect 12311 2859 12438 2981
rect 12311 2842 12351 2859
rect 12397 2842 12438 2859
rect 12311 2790 12348 2842
rect 12400 2790 12438 2842
rect 12311 2749 12438 2790
rect 12988 3698 13104 3807
rect 13660 3753 13775 3820
rect 12988 3652 13023 3698
rect 13069 3652 13104 3698
rect 12988 3584 13104 3652
rect 11354 2470 11470 2596
rect 12026 2692 12141 2749
rect 12026 2646 12061 2692
rect 12107 2646 12141 2692
rect 12026 2559 12141 2646
rect 12317 2692 12432 2749
rect 12317 2646 12351 2692
rect 12397 2646 12432 2692
rect 12317 2559 12432 2646
rect 12988 2596 13020 3584
rect 13072 2596 13104 3584
rect 13654 3712 13781 3753
rect 13654 3660 13692 3712
rect 13744 3660 13781 3712
rect 13654 3652 13695 3660
rect 13741 3652 13781 3660
rect 13654 3530 13781 3652
rect 13654 3495 13695 3530
rect 13741 3495 13781 3530
rect 13654 3443 13692 3495
rect 13744 3443 13781 3495
rect 13654 3363 13781 3443
rect 13654 3317 13695 3363
rect 13741 3317 13781 3363
rect 13654 3277 13781 3317
rect 13654 3225 13692 3277
rect 13744 3225 13781 3277
rect 13654 3195 13781 3225
rect 13654 3149 13695 3195
rect 13741 3149 13781 3195
rect 13654 3059 13781 3149
rect 13654 3007 13692 3059
rect 13744 3007 13781 3059
rect 13654 2981 13695 3007
rect 13741 2981 13781 3007
rect 13654 2859 13781 2981
rect 13654 2842 13695 2859
rect 13741 2842 13781 2859
rect 13654 2790 13692 2842
rect 13744 2790 13781 2842
rect 13654 2749 13781 2790
rect 12988 2470 13104 2596
rect 13660 2692 13775 2749
rect 13660 2646 13695 2692
rect 13741 2646 13775 2692
rect 13660 2559 13775 2646
rect 7327 2274 13864 2470
rect 7327 2228 7558 2274
rect 7604 2228 7716 2274
rect 7762 2228 7874 2274
rect 7920 2228 8032 2274
rect 8078 2228 8212 2274
rect 8258 2228 8370 2274
rect 8416 2228 8528 2274
rect 8574 2228 8686 2274
rect 8732 2228 9191 2274
rect 9237 2228 9349 2274
rect 9395 2228 9507 2274
rect 9553 2228 9665 2274
rect 9711 2228 9845 2274
rect 9891 2228 10003 2274
rect 10049 2228 10161 2274
rect 10207 2228 10319 2274
rect 10365 2228 10825 2274
rect 10871 2228 10983 2274
rect 11029 2228 11141 2274
rect 11187 2228 11299 2274
rect 11345 2228 11479 2274
rect 11525 2228 11637 2274
rect 11683 2228 11795 2274
rect 11841 2228 11953 2274
rect 11999 2228 12459 2274
rect 12505 2228 12617 2274
rect 12663 2228 12775 2274
rect 12821 2228 12933 2274
rect 12979 2228 13113 2274
rect 13159 2228 13271 2274
rect 13317 2228 13429 2274
rect 13475 2228 13587 2274
rect 13633 2228 13864 2274
rect 7327 2178 13864 2228
rect 7804 1917 7919 2178
rect 7803 1916 7919 1917
rect 8965 1926 9089 1966
rect 7802 1876 7926 1916
rect 7802 1824 7838 1876
rect 7890 1824 7926 1876
rect 8965 1874 9001 1926
rect 9053 1874 9089 1926
rect 7802 1816 7926 1824
rect 7802 1570 7838 1816
rect 7884 1658 7926 1816
rect 8062 1816 8108 1829
rect 7890 1606 7926 1658
rect 7884 1570 7926 1606
rect 7802 1566 7926 1570
rect 8028 1570 8062 1740
rect 8965 1771 9089 1874
rect 8108 1570 8143 1740
rect 8965 1708 9009 1771
rect 8965 1656 9001 1708
rect 8965 1631 9009 1656
rect 9055 1631 9089 1771
rect 8965 1616 9089 1631
rect 9208 1931 9254 2178
rect 9656 2008 13864 2178
rect 9656 1956 9900 2008
rect 9952 1956 10111 2008
rect 10163 1956 10321 2008
rect 10373 1956 10532 2008
rect 10584 1956 10743 2008
rect 10795 1956 10954 2008
rect 11006 1956 11165 2008
rect 11217 1956 11375 2008
rect 11427 1956 11586 2008
rect 11638 1956 11798 2008
rect 11850 1956 12009 2008
rect 12061 1956 12219 2008
rect 12271 1956 12430 2008
rect 12482 1956 12641 2008
rect 12693 1956 12852 2008
rect 12904 1956 13063 2008
rect 13115 1956 13273 2008
rect 13325 1956 13484 2008
rect 13536 1956 13864 2008
rect 9656 1948 13864 1956
rect 9208 1828 9254 1885
rect 9208 1725 9254 1782
rect 9208 1621 9254 1679
rect 7838 1557 7884 1566
rect 7182 1434 7306 1467
rect 8028 1434 8143 1570
rect 9208 1562 9254 1575
rect 9432 1931 9478 1944
rect 9432 1828 9478 1885
rect 9432 1725 9478 1782
rect 9432 1621 9478 1679
rect 9432 1475 9478 1575
rect 9656 1931 9960 1948
rect 9702 1902 9960 1931
rect 10006 1902 10118 1948
rect 10164 1902 10276 1948
rect 10322 1902 10434 1948
rect 10480 1902 10592 1948
rect 10638 1902 10750 1948
rect 10796 1902 10908 1948
rect 10954 1902 11066 1948
rect 11112 1902 11224 1948
rect 11270 1902 11383 1948
rect 11429 1902 11541 1948
rect 11587 1902 11699 1948
rect 11745 1902 11857 1948
rect 11903 1902 12015 1948
rect 12061 1902 12173 1948
rect 12219 1902 12332 1948
rect 12378 1902 12490 1948
rect 12536 1902 12648 1948
rect 12694 1902 12806 1948
rect 12852 1902 12964 1948
rect 13010 1902 13122 1948
rect 13168 1902 13280 1948
rect 13326 1902 13438 1948
rect 13484 1902 13596 1948
rect 13642 1902 13864 1948
rect 9702 1885 13864 1902
rect 9656 1828 13864 1885
rect 9702 1790 13864 1828
rect 9702 1782 9900 1790
rect 9656 1738 9900 1782
rect 9952 1784 10111 1790
rect 10163 1784 10321 1790
rect 10373 1784 10532 1790
rect 9952 1738 9960 1784
rect 10006 1738 10111 1784
rect 10164 1738 10276 1784
rect 10373 1738 10434 1784
rect 10480 1738 10532 1784
rect 10584 1784 10743 1790
rect 10795 1784 10954 1790
rect 10584 1738 10592 1784
rect 10638 1738 10743 1784
rect 10796 1738 10908 1784
rect 11006 1784 11165 1790
rect 11006 1738 11066 1784
rect 11112 1738 11165 1784
rect 11217 1784 11375 1790
rect 11427 1784 11586 1790
rect 11638 1784 11798 1790
rect 11217 1738 11224 1784
rect 11270 1738 11375 1784
rect 11429 1738 11541 1784
rect 11638 1738 11699 1784
rect 11745 1738 11798 1784
rect 11850 1784 12009 1790
rect 12061 1784 12219 1790
rect 11850 1738 11857 1784
rect 11903 1738 12009 1784
rect 12061 1738 12173 1784
rect 12271 1784 12430 1790
rect 12271 1738 12332 1784
rect 12378 1738 12430 1784
rect 12482 1784 12641 1790
rect 12693 1784 12852 1790
rect 12482 1738 12490 1784
rect 12536 1738 12641 1784
rect 12694 1738 12806 1784
rect 12904 1784 13063 1790
rect 12904 1738 12964 1784
rect 13010 1738 13063 1784
rect 13115 1784 13273 1790
rect 13325 1784 13484 1790
rect 13115 1738 13122 1784
rect 13168 1738 13273 1784
rect 13326 1738 13438 1784
rect 13536 1784 13864 1790
rect 13536 1738 13596 1784
rect 13642 1738 13864 1784
rect 9656 1725 13864 1738
rect 9702 1688 13864 1725
rect 9656 1621 9702 1679
rect 20764 1590 22476 1636
rect 9656 1562 9702 1575
rect 7180 1427 8143 1434
rect 7180 1375 7218 1427
rect 7270 1375 8143 1427
rect 8630 1451 8914 1463
rect 8630 1399 8642 1451
rect 8902 1399 8914 1451
rect 8630 1387 8754 1399
rect 8743 1386 8754 1387
rect 8800 1387 8914 1399
rect 8800 1386 8811 1387
rect 8743 1375 8811 1386
rect 7180 1300 8143 1375
rect 9192 1355 9478 1475
rect 9601 1451 9885 1463
rect 9601 1399 9613 1451
rect 9873 1399 9885 1451
rect 9601 1387 9885 1399
rect 7182 1209 7306 1300
rect 7182 1157 7218 1209
rect 7270 1157 7306 1209
rect 7182 1117 7306 1157
rect 7411 1183 7535 1200
rect 7411 1170 7778 1183
rect 7411 1160 7732 1170
rect 7411 1108 7447 1160
rect 7499 1124 7732 1160
rect 7499 1108 7778 1124
rect 7411 1035 7778 1108
rect 7411 989 7732 1035
rect 7411 942 7778 989
rect 7411 890 7447 942
rect 7499 900 7778 942
rect 7499 890 7732 900
rect 7411 854 7732 890
rect 7411 841 7778 854
rect 7956 1170 8002 1300
rect 8438 1183 8562 1218
rect 7956 1035 8002 1124
rect 7956 900 8002 989
rect 7956 841 8002 854
rect 8180 1178 8842 1183
rect 8180 1170 8474 1178
rect 8226 1126 8474 1170
rect 8526 1126 8842 1178
rect 8226 1124 8842 1126
rect 8180 1123 8842 1124
rect 8180 1077 8761 1123
rect 8807 1077 8842 1123
rect 8180 1035 8842 1077
rect 8226 989 8842 1035
rect 8180 960 8842 989
rect 8180 908 8474 960
rect 8526 919 8842 960
rect 8526 908 8761 919
rect 8180 900 8761 908
rect 8226 873 8761 900
rect 8807 873 8842 919
rect 8226 854 8842 873
rect 8180 841 8842 854
rect 8726 836 8842 841
rect 9192 1123 9271 1355
rect 9192 1077 9209 1123
rect 9255 1077 9271 1123
rect 9192 919 9271 1077
rect 9192 873 9209 919
rect 9255 873 9271 919
rect 7857 762 8113 773
rect 7857 756 7868 762
rect 6960 716 7868 756
rect 8102 756 8113 762
rect 9192 756 9271 873
rect 9622 1173 13649 1241
rect 9622 1123 9660 1173
rect 9622 1077 9657 1123
rect 9712 1121 9871 1173
rect 9923 1121 10082 1173
rect 10134 1121 10293 1173
rect 10345 1121 10504 1173
rect 10556 1121 10714 1173
rect 10766 1121 10925 1173
rect 10977 1121 11136 1173
rect 11188 1121 11347 1173
rect 11399 1121 11558 1173
rect 11610 1121 11769 1173
rect 11821 1121 11980 1173
rect 12032 1121 12191 1173
rect 12243 1121 12402 1173
rect 12454 1121 12612 1173
rect 12664 1121 12823 1173
rect 12875 1121 13034 1173
rect 13086 1121 13245 1173
rect 13297 1121 13456 1173
rect 13508 1121 13649 1173
rect 9703 1107 13649 1121
rect 9703 1077 9931 1107
rect 9622 1061 9931 1077
rect 9977 1061 10089 1107
rect 10135 1061 10247 1107
rect 10293 1061 10405 1107
rect 10451 1061 10563 1107
rect 10609 1061 10721 1107
rect 10767 1061 10879 1107
rect 10925 1061 11037 1107
rect 11083 1061 11195 1107
rect 11241 1061 11354 1107
rect 11400 1061 11512 1107
rect 11558 1061 11670 1107
rect 11716 1061 11828 1107
rect 11874 1061 11986 1107
rect 12032 1061 12144 1107
rect 12190 1061 12303 1107
rect 12349 1061 12461 1107
rect 12507 1061 12619 1107
rect 12665 1061 12777 1107
rect 12823 1061 12935 1107
rect 12981 1061 13093 1107
rect 13139 1061 13251 1107
rect 13297 1061 13409 1107
rect 13455 1061 13567 1107
rect 13613 1061 13649 1107
rect 9622 955 13649 1061
rect 9622 919 9660 955
rect 9622 873 9657 919
rect 9712 903 9871 955
rect 9923 943 10082 955
rect 10134 943 10293 955
rect 9923 903 9931 943
rect 9703 897 9931 903
rect 9977 903 10082 943
rect 9977 897 10089 903
rect 10135 897 10247 943
rect 10345 943 10504 955
rect 10345 903 10405 943
rect 10293 897 10405 903
rect 10451 903 10504 943
rect 10556 943 10714 955
rect 10766 943 10925 955
rect 10556 903 10563 943
rect 10451 897 10563 903
rect 10609 903 10714 943
rect 10609 897 10721 903
rect 10767 897 10879 943
rect 10977 943 11136 955
rect 10977 903 11037 943
rect 10925 897 11037 903
rect 11083 903 11136 943
rect 11188 943 11347 955
rect 11399 943 11558 955
rect 11188 903 11195 943
rect 11083 897 11195 903
rect 11241 903 11347 943
rect 11241 897 11354 903
rect 11400 897 11512 943
rect 11610 943 11769 955
rect 11610 903 11670 943
rect 11558 897 11670 903
rect 11716 903 11769 943
rect 11821 943 11980 955
rect 12032 943 12191 955
rect 11821 903 11828 943
rect 11716 897 11828 903
rect 11874 903 11980 943
rect 11874 897 11986 903
rect 12032 897 12144 943
rect 12190 903 12191 943
rect 12243 943 12402 955
rect 12243 903 12303 943
rect 12190 897 12303 903
rect 12349 903 12402 943
rect 12454 943 12612 955
rect 12664 943 12823 955
rect 12454 903 12461 943
rect 12349 897 12461 903
rect 12507 903 12612 943
rect 12507 897 12619 903
rect 12665 897 12777 943
rect 12875 943 13034 955
rect 12875 903 12935 943
rect 12823 897 12935 903
rect 12981 903 13034 943
rect 13086 943 13245 955
rect 13297 943 13456 955
rect 13086 903 13093 943
rect 12981 897 13093 903
rect 13139 903 13245 943
rect 13139 897 13251 903
rect 13297 897 13409 943
rect 13455 903 13456 943
rect 13508 943 13649 955
rect 13508 903 13567 943
rect 13455 897 13567 903
rect 13613 897 13649 943
rect 9703 873 13649 897
rect 9622 836 13649 873
rect 8102 716 9271 756
rect 6960 636 9271 716
rect 22430 439 22476 1590
rect 28007 1130 28136 17115
rect 28007 1078 28045 1130
rect 28097 1078 28136 1130
rect 28007 912 28136 1078
rect 28007 860 28045 912
rect 28097 860 28136 912
rect 28007 694 28136 860
rect 28007 642 28045 694
rect 28097 642 28136 694
rect 28007 602 28136 642
rect 28248 1130 28378 17342
rect 28248 1078 28287 1130
rect 28339 1078 28378 1130
rect 28248 912 28378 1078
rect 28248 860 28287 912
rect 28339 860 28378 912
rect 28248 694 28378 860
rect 28248 642 28287 694
rect 28339 642 28378 694
rect 28248 602 28378 642
rect 28490 1130 28619 17568
rect 28490 1078 28529 1130
rect 28581 1078 28619 1130
rect 28490 912 28619 1078
rect 28490 860 28529 912
rect 28581 860 28619 912
rect 28490 694 28619 860
rect 28490 642 28529 694
rect 28581 642 28619 694
rect 28490 602 28619 642
rect 28731 1130 28861 17795
rect 29520 1155 29654 28726
rect 28731 1078 28770 1130
rect 28822 1078 28861 1130
rect 28731 912 28861 1078
rect 28731 860 28770 912
rect 28822 860 28861 912
rect 28731 694 28861 860
rect 29525 1117 29649 1155
rect 29525 1065 29561 1117
rect 29613 1065 29649 1117
rect 29525 899 29649 1065
rect 29525 847 29561 899
rect 29613 847 29649 899
rect 29525 807 29649 847
rect 28731 642 28770 694
rect 28822 642 28861 694
rect 28731 602 28861 642
rect 403 289 9220 330
rect 403 237 8918 289
rect 8970 237 9130 289
rect 9182 237 9220 289
rect 403 185 733 237
rect 785 185 945 237
rect 997 185 9220 237
rect 27841 237 29415 330
rect 403 71 9220 185
rect 13144 144 14721 190
rect 27841 185 29059 237
rect 29111 185 29271 237
rect 29323 185 29415 237
rect 403 19 8918 71
rect 8970 19 9130 71
rect 9182 19 9220 71
rect 403 -33 733 19
rect 785 -33 945 19
rect 997 -33 9220 19
rect 403 -126 9220 -33
rect 27841 19 29415 185
rect 27841 -33 29059 19
rect 29111 -33 29271 19
rect 29323 -33 29415 19
rect 27841 -126 29415 -33
<< via1 >>
rect 444 28944 496 28996
rect 444 28726 496 28778
rect 1656 28489 1659 28500
rect 1659 28489 1705 28500
rect 1705 28489 1708 28500
rect 1656 28448 1708 28489
rect 1656 28279 1659 28282
rect 1659 28279 1705 28282
rect 1705 28279 1708 28282
rect 1656 28230 1708 28279
rect 1656 28012 1708 28064
rect 1656 27804 1708 27846
rect 1656 27794 1659 27804
rect 1659 27794 1705 27804
rect 1705 27794 1708 27804
rect 2096 28489 2107 28500
rect 2107 28489 2148 28500
rect 2096 28448 2148 28489
rect 2096 28279 2107 28282
rect 2107 28279 2148 28282
rect 2096 28230 2148 28279
rect 2096 28012 2148 28064
rect 2096 27804 2148 27846
rect 2096 27794 2107 27804
rect 2107 27794 2148 27804
rect 2328 28489 2331 28500
rect 2331 28489 2377 28500
rect 2377 28489 2380 28500
rect 2328 28448 2380 28489
rect 2328 28279 2331 28282
rect 2331 28279 2377 28282
rect 2377 28279 2380 28282
rect 2328 28230 2380 28279
rect 2328 28012 2380 28064
rect 2328 27804 2380 27846
rect 2328 27794 2331 27804
rect 2331 27794 2377 27804
rect 2377 27794 2380 27804
rect 2776 28489 2779 28500
rect 2779 28489 2825 28500
rect 2825 28489 2828 28500
rect 2776 28448 2828 28489
rect 2776 28279 2779 28282
rect 2779 28279 2825 28282
rect 2825 28279 2828 28282
rect 2776 28230 2828 28279
rect 2776 28012 2828 28064
rect 2776 27804 2828 27846
rect 2776 27794 2779 27804
rect 2779 27794 2825 27804
rect 2825 27794 2828 27804
rect 3008 28489 3049 28500
rect 3049 28489 3060 28500
rect 3008 28448 3060 28489
rect 3008 28279 3049 28282
rect 3049 28279 3060 28282
rect 3008 28230 3060 28279
rect 3008 28012 3060 28064
rect 3008 27804 3060 27846
rect 3008 27794 3049 27804
rect 3049 27794 3060 27804
rect 3448 28489 3451 28500
rect 3451 28489 3497 28500
rect 3497 28489 3500 28500
rect 3448 28448 3500 28489
rect 3448 28279 3451 28282
rect 3451 28279 3497 28282
rect 3497 28279 3500 28282
rect 3448 28230 3500 28279
rect 3448 28012 3500 28064
rect 1656 27347 1708 27353
rect 1656 27301 1659 27347
rect 1659 27301 1705 27347
rect 1705 27301 1708 27347
rect 1656 27091 1659 27135
rect 1659 27091 1705 27135
rect 1705 27091 1708 27135
rect 1656 27083 1708 27091
rect 1656 26881 1659 26917
rect 1659 26881 1705 26917
rect 1705 26881 1708 26917
rect 1656 26865 1708 26881
rect 3448 27804 3500 27846
rect 3448 27794 3451 27804
rect 3451 27794 3497 27804
rect 3497 27794 3500 27804
rect 3888 28489 3899 28500
rect 3899 28489 3940 28500
rect 3888 28448 3940 28489
rect 3888 28279 3899 28282
rect 3899 28279 3940 28282
rect 3888 28230 3940 28279
rect 3888 28012 3940 28064
rect 2104 27347 2156 27353
rect 2104 27301 2107 27347
rect 2107 27301 2153 27347
rect 2153 27301 2156 27347
rect 2104 27091 2107 27135
rect 2107 27091 2153 27135
rect 2153 27091 2156 27135
rect 2104 27083 2156 27091
rect 2104 26881 2107 26917
rect 2107 26881 2153 26917
rect 2153 26881 2156 26917
rect 2104 26865 2156 26881
rect 2552 27347 2604 27353
rect 2552 27301 2555 27347
rect 2555 27301 2601 27347
rect 2601 27301 2604 27347
rect 2552 27091 2555 27135
rect 2555 27091 2601 27135
rect 2601 27091 2604 27135
rect 2552 27083 2604 27091
rect 2552 26881 2555 26917
rect 2555 26881 2601 26917
rect 2601 26881 2604 26917
rect 2552 26865 2604 26881
rect 3888 27804 3940 27846
rect 3888 27794 3899 27804
rect 3899 27794 3940 27804
rect 4120 28489 4123 28500
rect 4123 28489 4169 28500
rect 4169 28489 4172 28500
rect 4120 28448 4172 28489
rect 4120 28279 4123 28282
rect 4123 28279 4169 28282
rect 4169 28279 4172 28282
rect 4120 28230 4172 28279
rect 4120 28012 4172 28064
rect 4120 27804 4172 27846
rect 4120 27794 4123 27804
rect 4123 27794 4169 27804
rect 4169 27794 4172 27804
rect 4568 28489 4571 28500
rect 4571 28489 4617 28500
rect 4617 28489 4620 28500
rect 4568 28448 4620 28489
rect 4568 28279 4571 28282
rect 4571 28279 4617 28282
rect 4617 28279 4620 28282
rect 4568 28230 4620 28279
rect 4568 28012 4620 28064
rect 4568 27804 4620 27846
rect 4568 27794 4571 27804
rect 4571 27794 4617 27804
rect 4617 27794 4620 27804
rect 4800 28489 4841 28500
rect 4841 28489 4852 28500
rect 4800 28448 4852 28489
rect 4800 28279 4841 28282
rect 4841 28279 4852 28282
rect 4800 28230 4852 28279
rect 4800 28012 4852 28064
rect 4800 27804 4852 27846
rect 4800 27794 4841 27804
rect 4841 27794 4852 27804
rect 5240 28489 5243 28500
rect 5243 28489 5289 28500
rect 5289 28489 5292 28500
rect 5240 28448 5292 28489
rect 5240 28279 5243 28282
rect 5243 28279 5289 28282
rect 5289 28279 5292 28282
rect 5240 28230 5292 28279
rect 5240 28012 5292 28064
rect 5923 28349 5975 28401
rect 5923 28131 5975 28183
rect 6362 28349 6414 28401
rect 9035 28489 9038 28500
rect 9038 28489 9084 28500
rect 9084 28489 9087 28500
rect 9035 28448 9087 28489
rect 7746 28292 7798 28344
rect 5923 27913 5933 27965
rect 5933 27913 5975 27965
rect 3000 27347 3052 27353
rect 3000 27301 3003 27347
rect 3003 27301 3049 27347
rect 3049 27301 3052 27347
rect 3000 27091 3003 27135
rect 3003 27091 3049 27135
rect 3049 27091 3052 27135
rect 3000 27083 3052 27091
rect 3000 26881 3003 26917
rect 3003 26881 3049 26917
rect 3049 26881 3052 26917
rect 3000 26865 3052 26881
rect 3448 27347 3500 27353
rect 3448 27301 3451 27347
rect 3451 27301 3497 27347
rect 3497 27301 3500 27347
rect 3448 27091 3451 27135
rect 3451 27091 3497 27135
rect 3497 27091 3500 27135
rect 3448 27083 3500 27091
rect 3448 26881 3451 26917
rect 3451 26881 3497 26917
rect 3497 26881 3500 26917
rect 3448 26865 3500 26881
rect 5240 27804 5292 27846
rect 5240 27794 5243 27804
rect 5243 27794 5289 27804
rect 5289 27794 5292 27804
rect 6362 28131 6414 28183
rect 6362 27913 6381 27965
rect 6381 27913 6414 27965
rect 6582 28133 6634 28185
rect 7746 28074 7798 28126
rect 6582 27915 6587 27967
rect 6587 27915 6633 27967
rect 6633 27915 6634 27967
rect 5837 27637 5854 27683
rect 5854 27637 5993 27683
rect 5837 27631 5993 27637
rect 7746 27876 7798 27908
rect 7746 27856 7751 27876
rect 7751 27856 7797 27876
rect 7797 27856 7798 27876
rect 9035 28279 9038 28282
rect 9038 28279 9084 28282
rect 9084 28279 9087 28282
rect 9035 28230 9087 28279
rect 9035 28012 9087 28064
rect 9035 27804 9087 27846
rect 9035 27794 9038 27804
rect 9038 27794 9084 27804
rect 9084 27794 9087 27804
rect 9475 28489 9486 28500
rect 9486 28489 9527 28500
rect 9475 28448 9527 28489
rect 9475 28279 9486 28282
rect 9486 28279 9527 28282
rect 9475 28230 9527 28279
rect 9475 28012 9527 28064
rect 6765 27631 6921 27683
rect 3896 27347 3948 27353
rect 3896 27301 3899 27347
rect 3899 27301 3945 27347
rect 3945 27301 3948 27347
rect 3896 27091 3899 27135
rect 3899 27091 3945 27135
rect 3945 27091 3948 27135
rect 3896 27083 3948 27091
rect 3896 26881 3899 26917
rect 3899 26881 3945 26917
rect 3945 26881 3948 26917
rect 3896 26865 3948 26881
rect 4344 27347 4396 27353
rect 4344 27301 4347 27347
rect 4347 27301 4393 27347
rect 4393 27301 4396 27347
rect 4344 27091 4347 27135
rect 4347 27091 4393 27135
rect 4393 27091 4396 27135
rect 4344 27083 4396 27091
rect 4344 26881 4347 26917
rect 4347 26881 4393 26917
rect 4393 26881 4396 26917
rect 4344 26865 4396 26881
rect 4792 27347 4844 27353
rect 4792 27301 4795 27347
rect 4795 27301 4841 27347
rect 4841 27301 4844 27347
rect 4792 27091 4795 27135
rect 4795 27091 4841 27135
rect 4841 27091 4844 27135
rect 4792 27083 4844 27091
rect 4792 26881 4795 26917
rect 4795 26881 4841 26917
rect 4841 26881 4844 26917
rect 4792 26865 4844 26881
rect 5240 27347 5292 27353
rect 5240 27301 5243 27347
rect 5243 27301 5289 27347
rect 5289 27301 5292 27347
rect 5240 27091 5243 27135
rect 5243 27091 5289 27135
rect 5289 27091 5292 27135
rect 5240 27083 5292 27091
rect 5647 27326 5649 27378
rect 5649 27326 5695 27378
rect 5695 27326 5699 27378
rect 5647 27144 5649 27160
rect 5649 27144 5695 27160
rect 5695 27144 5699 27160
rect 5647 27108 5699 27144
rect 5923 27336 5933 27378
rect 5933 27336 5975 27378
rect 5923 27326 5975 27336
rect 5923 27132 5933 27160
rect 5933 27132 5975 27160
rect 5923 27108 5975 27132
rect 8778 27643 8830 27695
rect 9475 27804 9527 27846
rect 9475 27794 9486 27804
rect 9486 27794 9527 27804
rect 9707 28489 9710 28500
rect 9710 28489 9756 28500
rect 9756 28489 9759 28500
rect 9707 28448 9759 28489
rect 9707 28279 9710 28282
rect 9710 28279 9756 28282
rect 9756 28279 9759 28282
rect 9707 28230 9759 28279
rect 9707 28012 9759 28064
rect 9707 27804 9759 27846
rect 9707 27794 9710 27804
rect 9710 27794 9756 27804
rect 9756 27794 9759 27804
rect 10155 28489 10158 28500
rect 10158 28489 10204 28500
rect 10204 28489 10207 28500
rect 10155 28448 10207 28489
rect 10155 28279 10158 28282
rect 10158 28279 10204 28282
rect 10204 28279 10207 28282
rect 10155 28230 10207 28279
rect 10155 28012 10207 28064
rect 10155 27804 10207 27846
rect 10155 27794 10158 27804
rect 10158 27794 10204 27804
rect 10204 27794 10207 27804
rect 10387 28489 10428 28500
rect 10428 28489 10439 28500
rect 10387 28448 10439 28489
rect 10387 28279 10428 28282
rect 10428 28279 10439 28282
rect 10387 28230 10439 28279
rect 10387 28012 10439 28064
rect 10387 27804 10439 27846
rect 10387 27794 10428 27804
rect 10428 27794 10439 27804
rect 10827 28489 10830 28500
rect 10830 28489 10876 28500
rect 10876 28489 10879 28500
rect 10827 28448 10879 28489
rect 10827 28279 10830 28282
rect 10830 28279 10876 28282
rect 10876 28279 10879 28282
rect 10827 28230 10879 28279
rect 10827 28012 10879 28064
rect 5240 26881 5243 26917
rect 5243 26881 5289 26917
rect 5289 26881 5292 26917
rect 5240 26865 5292 26881
rect 7007 27158 7059 27210
rect 7219 27158 7271 27210
rect 8136 27378 8188 27392
rect 8136 27340 8141 27378
rect 8141 27340 8187 27378
rect 8187 27340 8188 27378
rect 8778 27425 8830 27477
rect 8136 27144 8141 27174
rect 8141 27144 8187 27174
rect 8187 27144 8188 27174
rect 8136 27122 8188 27144
rect 9035 27347 9087 27353
rect 9035 27301 9038 27347
rect 9038 27301 9084 27347
rect 9084 27301 9087 27347
rect 9035 27091 9038 27135
rect 9038 27091 9084 27135
rect 9084 27091 9087 27135
rect 9035 27083 9087 27091
rect 7005 26922 7057 26974
rect 7217 26922 7269 26974
rect 9035 26881 9038 26917
rect 9038 26881 9084 26917
rect 9084 26881 9087 26917
rect 9035 26865 9087 26881
rect 10827 27804 10879 27846
rect 10827 27794 10830 27804
rect 10830 27794 10876 27804
rect 10876 27794 10879 27804
rect 11267 28489 11278 28500
rect 11278 28489 11319 28500
rect 11267 28448 11319 28489
rect 11267 28279 11278 28282
rect 11278 28279 11319 28282
rect 11267 28230 11319 28279
rect 11267 28012 11319 28064
rect 5874 26462 5926 26514
rect 6081 26462 6091 26514
rect 6091 26462 6133 26514
rect 5874 26244 5926 26296
rect 6081 26276 6091 26296
rect 6091 26276 6133 26296
rect 6081 26244 6133 26276
rect 5874 26026 5926 26078
rect 6081 26070 6091 26078
rect 6091 26070 6133 26078
rect 6081 26026 6133 26070
rect 5874 25808 5926 25860
rect 6081 25808 6133 25860
rect 6601 26446 6653 26491
rect 6601 26439 6605 26446
rect 6605 26439 6651 26446
rect 6651 26439 6653 26446
rect 7565 26462 7617 26514
rect 7772 26462 7782 26514
rect 7782 26462 7824 26514
rect 6601 26230 6653 26273
rect 6601 26221 6605 26230
rect 6605 26221 6651 26230
rect 6651 26221 6653 26230
rect 6601 26014 6653 26055
rect 6601 26003 6605 26014
rect 6605 26003 6651 26014
rect 6651 26003 6653 26014
rect 6601 25798 6653 25837
rect 6601 25785 6605 25798
rect 6605 25785 6651 25798
rect 6651 25785 6653 25798
rect 5874 25169 5926 25221
rect 6086 25218 6138 25221
rect 6086 25172 6112 25218
rect 6112 25172 6138 25218
rect 6086 25169 6138 25172
rect 1817 24721 1869 24773
rect 1817 24550 1869 24556
rect 1817 24504 1863 24550
rect 1863 24504 1869 24550
rect 1817 24286 1863 24338
rect 1863 24286 1869 24338
rect 1817 24069 1863 24121
rect 1863 24069 1869 24121
rect 1817 23851 1863 23903
rect 1863 23851 1869 23903
rect 1817 23633 1863 23685
rect 1863 23633 1869 23685
rect 1817 23415 1863 23467
rect 1863 23415 1869 23467
rect 1817 23198 1863 23250
rect 1863 23198 1869 23250
rect 1817 22980 1863 23032
rect 1863 22980 1869 23032
rect 1817 22763 1863 22815
rect 1863 22763 1869 22815
rect 2269 24721 2321 24773
rect 2552 24721 2604 24773
rect 2835 24721 2887 24773
rect 2269 24550 2321 24556
rect 2269 24504 2311 24550
rect 2311 24504 2321 24550
rect 2552 24504 2604 24556
rect 2835 24550 2887 24556
rect 2835 24504 2845 24550
rect 2845 24504 2887 24550
rect 2269 24286 2311 24338
rect 2311 24286 2321 24338
rect 2552 24286 2604 24338
rect 2835 24286 2845 24338
rect 2845 24286 2887 24338
rect 2269 24069 2311 24121
rect 2311 24069 2321 24121
rect 2552 24069 2604 24121
rect 2835 24069 2845 24121
rect 2845 24069 2887 24121
rect 2269 23851 2311 23903
rect 2311 23851 2321 23903
rect 2552 23851 2604 23903
rect 2835 23851 2845 23903
rect 2845 23851 2887 23903
rect 2269 23633 2311 23685
rect 2311 23633 2321 23685
rect 2552 23633 2604 23685
rect 2835 23633 2845 23685
rect 2845 23633 2887 23685
rect 2269 23415 2311 23467
rect 2311 23415 2321 23467
rect 2552 23415 2604 23467
rect 2835 23415 2845 23467
rect 2845 23415 2887 23467
rect 2269 23198 2311 23250
rect 2311 23198 2321 23250
rect 2552 23198 2604 23250
rect 2835 23198 2845 23250
rect 2845 23198 2887 23250
rect 2269 22980 2311 23032
rect 2311 22980 2321 23032
rect 2552 22980 2604 23032
rect 2835 22980 2845 23032
rect 2845 22980 2887 23032
rect 2269 22763 2311 22815
rect 2311 22763 2321 22815
rect 2552 22763 2604 22815
rect 2835 22763 2845 22815
rect 2845 22763 2887 22815
rect 2039 21790 2091 21842
rect 2039 21582 2091 21624
rect 2039 21572 2041 21582
rect 2041 21572 2087 21582
rect 2087 21572 2091 21582
rect 3287 24721 3339 24773
rect 3287 24550 3339 24556
rect 3287 24504 3293 24550
rect 3293 24504 3339 24550
rect 3287 24286 3293 24338
rect 3293 24286 3339 24338
rect 3287 24069 3293 24121
rect 3293 24069 3339 24121
rect 3287 23851 3293 23903
rect 3293 23851 3339 23903
rect 3287 23633 3293 23685
rect 3293 23633 3339 23685
rect 3287 23415 3293 23467
rect 3293 23415 3339 23467
rect 3287 23198 3293 23250
rect 3293 23198 3339 23250
rect 3287 22980 3293 23032
rect 3293 22980 3339 23032
rect 3287 22763 3293 22815
rect 3293 22763 3339 22815
rect 3609 24721 3661 24773
rect 3609 24550 3661 24556
rect 3609 24504 3655 24550
rect 3655 24504 3661 24550
rect 3609 24286 3655 24338
rect 3655 24286 3661 24338
rect 3609 24069 3655 24121
rect 3655 24069 3661 24121
rect 3609 23851 3655 23903
rect 3655 23851 3661 23903
rect 3609 23633 3655 23685
rect 3655 23633 3661 23685
rect 3609 23415 3655 23467
rect 3655 23415 3661 23467
rect 3609 23198 3655 23250
rect 3655 23198 3661 23250
rect 3609 22980 3655 23032
rect 3655 22980 3661 23032
rect 3609 22763 3655 22815
rect 3655 22763 3661 22815
rect 3065 21790 3117 21842
rect 3065 21582 3117 21624
rect 3065 21572 3069 21582
rect 3069 21572 3115 21582
rect 3115 21572 3117 21582
rect 4061 24721 4113 24773
rect 4344 24721 4396 24773
rect 4627 24721 4679 24773
rect 4061 24550 4113 24556
rect 4061 24504 4103 24550
rect 4103 24504 4113 24550
rect 4344 24504 4396 24556
rect 4627 24550 4679 24556
rect 4627 24504 4637 24550
rect 4637 24504 4679 24550
rect 4061 24286 4103 24338
rect 4103 24286 4113 24338
rect 4344 24286 4396 24338
rect 4627 24286 4637 24338
rect 4637 24286 4679 24338
rect 4061 24069 4103 24121
rect 4103 24069 4113 24121
rect 4344 24069 4396 24121
rect 4627 24069 4637 24121
rect 4637 24069 4679 24121
rect 4061 23851 4103 23903
rect 4103 23851 4113 23903
rect 4344 23851 4396 23903
rect 4627 23851 4637 23903
rect 4637 23851 4679 23903
rect 4061 23633 4103 23685
rect 4103 23633 4113 23685
rect 4344 23633 4396 23685
rect 4627 23633 4637 23685
rect 4637 23633 4679 23685
rect 4061 23415 4103 23467
rect 4103 23415 4113 23467
rect 4344 23415 4396 23467
rect 4627 23415 4637 23467
rect 4637 23415 4679 23467
rect 4061 23198 4103 23250
rect 4103 23198 4113 23250
rect 4344 23198 4396 23250
rect 4627 23198 4637 23250
rect 4637 23198 4679 23250
rect 4061 22980 4103 23032
rect 4103 22980 4113 23032
rect 4344 22980 4396 23032
rect 4627 22980 4637 23032
rect 4637 22980 4679 23032
rect 4061 22763 4103 22815
rect 4103 22763 4113 22815
rect 4344 22763 4396 22815
rect 4627 22763 4637 22815
rect 4637 22763 4679 22815
rect 3831 21790 3883 21842
rect 3831 21582 3883 21624
rect 3831 21572 3833 21582
rect 3833 21572 3879 21582
rect 3879 21572 3883 21582
rect 5079 24721 5131 24773
rect 5079 24550 5131 24556
rect 5079 24504 5085 24550
rect 5085 24504 5131 24550
rect 5079 24286 5085 24338
rect 5085 24286 5131 24338
rect 5079 24069 5085 24121
rect 5085 24069 5131 24121
rect 5079 23851 5085 23903
rect 5085 23851 5131 23903
rect 5079 23633 5085 23685
rect 5085 23633 5131 23685
rect 5079 23415 5085 23467
rect 5085 23415 5131 23467
rect 5079 23198 5085 23250
rect 5085 23198 5131 23250
rect 5079 22980 5085 23032
rect 5085 22980 5131 23032
rect 5079 22763 5085 22815
rect 5085 22763 5131 22815
rect 6094 24750 6137 24802
rect 6137 24750 6146 24802
rect 6094 24533 6137 24585
rect 6137 24533 6146 24585
rect 6094 24315 6137 24367
rect 6137 24315 6146 24367
rect 6094 24098 6137 24150
rect 6137 24098 6146 24150
rect 6094 23880 6137 23932
rect 6137 23880 6146 23932
rect 6094 23662 6137 23714
rect 6137 23662 6146 23714
rect 6094 23444 6137 23496
rect 6137 23444 6146 23496
rect 6094 23227 6137 23279
rect 6137 23227 6146 23279
rect 6094 23009 6137 23061
rect 6137 23009 6146 23061
rect 6094 22792 6137 22844
rect 6137 22792 6146 22844
rect 4857 21790 4909 21842
rect 4857 21582 4909 21624
rect 4857 21572 4861 21582
rect 4861 21572 4907 21582
rect 4907 21572 4909 21582
rect 7565 26244 7617 26296
rect 7772 26276 7782 26296
rect 7782 26276 7824 26296
rect 7772 26244 7824 26276
rect 7565 26026 7617 26078
rect 7772 26070 7782 26078
rect 7782 26070 7824 26078
rect 7772 26026 7824 26070
rect 7565 25808 7617 25860
rect 7772 25808 7824 25860
rect 8292 26446 8344 26491
rect 8292 26439 8296 26446
rect 8296 26439 8342 26446
rect 8342 26439 8344 26446
rect 8292 26230 8344 26273
rect 8292 26221 8296 26230
rect 8296 26221 8342 26230
rect 8342 26221 8344 26230
rect 8292 26014 8344 26055
rect 8292 26003 8296 26014
rect 8296 26003 8342 26014
rect 8342 26003 8344 26014
rect 8292 25798 8344 25837
rect 8292 25785 8296 25798
rect 8296 25785 8342 25798
rect 8342 25785 8344 25798
rect 7565 25169 7617 25221
rect 7777 25218 7829 25221
rect 7777 25172 7803 25218
rect 7803 25172 7829 25218
rect 7777 25169 7829 25172
rect 6608 24759 6651 24811
rect 6651 24759 6660 24811
rect 6608 24541 6651 24593
rect 6651 24541 6660 24593
rect 6608 24324 6651 24376
rect 6651 24324 6660 24376
rect 6608 24106 6651 24158
rect 6651 24106 6660 24158
rect 6608 23888 6651 23940
rect 6651 23888 6660 23940
rect 6608 23670 6651 23722
rect 6651 23670 6660 23722
rect 6608 23453 6651 23505
rect 6651 23453 6660 23505
rect 6608 23267 6660 23287
rect 6608 23235 6651 23267
rect 6651 23235 6660 23267
rect 7785 24750 7828 24802
rect 7828 24750 7837 24802
rect 7785 24533 7828 24585
rect 7828 24533 7837 24585
rect 7785 24315 7828 24367
rect 7828 24315 7837 24367
rect 7785 24098 7828 24150
rect 7828 24098 7837 24150
rect 7785 23880 7828 23932
rect 7828 23880 7837 23932
rect 7785 23662 7828 23714
rect 7828 23662 7837 23714
rect 7785 23444 7828 23496
rect 7828 23444 7837 23496
rect 7785 23227 7828 23279
rect 7828 23227 7837 23279
rect 7785 23009 7828 23061
rect 7828 23009 7837 23061
rect 6825 22651 6877 22703
rect 6825 22443 6877 22485
rect 6825 22433 6829 22443
rect 6829 22433 6875 22443
rect 6875 22433 6877 22443
rect 7785 22792 7828 22844
rect 7828 22792 7837 22844
rect 6311 21744 6315 21796
rect 6315 21744 6361 21796
rect 6361 21744 6363 21796
rect 6311 21526 6315 21578
rect 6315 21526 6361 21578
rect 6361 21526 6363 21578
rect 9483 27347 9535 27353
rect 9483 27301 9486 27347
rect 9486 27301 9532 27347
rect 9532 27301 9535 27347
rect 9483 27091 9486 27135
rect 9486 27091 9532 27135
rect 9532 27091 9535 27135
rect 9483 27083 9535 27091
rect 9483 26881 9486 26917
rect 9486 26881 9532 26917
rect 9532 26881 9535 26917
rect 9483 26865 9535 26881
rect 9931 27347 9983 27353
rect 9931 27301 9934 27347
rect 9934 27301 9980 27347
rect 9980 27301 9983 27347
rect 9931 27091 9934 27135
rect 9934 27091 9980 27135
rect 9980 27091 9983 27135
rect 9931 27083 9983 27091
rect 9931 26881 9934 26917
rect 9934 26881 9980 26917
rect 9980 26881 9983 26917
rect 9931 26865 9983 26881
rect 11267 27804 11319 27846
rect 11267 27794 11278 27804
rect 11278 27794 11319 27804
rect 29561 28944 29613 28996
rect 11499 28489 11502 28500
rect 11502 28489 11548 28500
rect 11548 28489 11551 28500
rect 11499 28448 11551 28489
rect 11499 28279 11502 28282
rect 11502 28279 11548 28282
rect 11548 28279 11551 28282
rect 11499 28230 11551 28279
rect 11499 28012 11551 28064
rect 11499 27804 11551 27846
rect 11499 27794 11502 27804
rect 11502 27794 11548 27804
rect 11548 27794 11551 27804
rect 11947 28489 11950 28500
rect 11950 28489 11996 28500
rect 11996 28489 11999 28500
rect 11947 28448 11999 28489
rect 11947 28279 11950 28282
rect 11950 28279 11996 28282
rect 11996 28279 11999 28282
rect 11947 28230 11999 28279
rect 11947 28012 11999 28064
rect 11947 27804 11999 27846
rect 11947 27794 11950 27804
rect 11950 27794 11996 27804
rect 11996 27794 11999 27804
rect 12179 28489 12220 28500
rect 12220 28489 12231 28500
rect 12179 28448 12231 28489
rect 12179 28279 12220 28282
rect 12220 28279 12231 28282
rect 12179 28230 12231 28279
rect 12179 28012 12231 28064
rect 12179 27804 12231 27846
rect 12179 27794 12220 27804
rect 12220 27794 12231 27804
rect 12619 28489 12622 28500
rect 12622 28489 12668 28500
rect 12668 28489 12671 28500
rect 12619 28448 12671 28489
rect 12619 28279 12622 28282
rect 12622 28279 12668 28282
rect 12668 28279 12671 28282
rect 12619 28230 12671 28279
rect 12619 28012 12671 28064
rect 13302 28349 13354 28401
rect 13302 28131 13354 28183
rect 13741 28349 13793 28401
rect 29561 28726 29613 28778
rect 15125 28292 15177 28344
rect 13302 27913 13312 27965
rect 13312 27913 13354 27965
rect 10379 27347 10431 27353
rect 10379 27301 10382 27347
rect 10382 27301 10428 27347
rect 10428 27301 10431 27347
rect 10379 27091 10382 27135
rect 10382 27091 10428 27135
rect 10428 27091 10431 27135
rect 10379 27083 10431 27091
rect 10379 26881 10382 26917
rect 10382 26881 10428 26917
rect 10428 26881 10431 26917
rect 10379 26865 10431 26881
rect 10827 27347 10879 27353
rect 10827 27301 10830 27347
rect 10830 27301 10876 27347
rect 10876 27301 10879 27347
rect 10827 27091 10830 27135
rect 10830 27091 10876 27135
rect 10876 27091 10879 27135
rect 10827 27083 10879 27091
rect 10827 26881 10830 26917
rect 10830 26881 10876 26917
rect 10876 26881 10879 26917
rect 10827 26865 10879 26881
rect 12619 27804 12671 27846
rect 12619 27794 12622 27804
rect 12622 27794 12668 27804
rect 12668 27794 12671 27804
rect 13741 28131 13793 28183
rect 13741 27913 13760 27965
rect 13760 27913 13793 27965
rect 13961 28133 14013 28185
rect 16918 28340 16970 28392
rect 17828 28340 17880 28392
rect 18552 28340 18604 28392
rect 19462 28340 19514 28392
rect 20185 28340 20237 28392
rect 21095 28340 21147 28392
rect 21819 28340 21871 28392
rect 22729 28340 22781 28392
rect 23787 28361 23839 28401
rect 24226 28361 24278 28401
rect 23787 28349 23839 28361
rect 24226 28349 24278 28361
rect 15125 28074 15177 28126
rect 16918 28122 16970 28174
rect 13961 27915 13966 27967
rect 13966 27915 14012 27967
rect 14012 27915 14013 27967
rect 13216 27637 13233 27683
rect 13233 27637 13372 27683
rect 13216 27631 13372 27637
rect 15125 27876 15177 27908
rect 15125 27856 15130 27876
rect 15130 27856 15176 27876
rect 15176 27856 15177 27876
rect 14144 27631 14300 27683
rect 11275 27347 11327 27353
rect 11275 27301 11278 27347
rect 11278 27301 11324 27347
rect 11324 27301 11327 27347
rect 11275 27091 11278 27135
rect 11278 27091 11324 27135
rect 11324 27091 11327 27135
rect 11275 27083 11327 27091
rect 11275 26881 11278 26917
rect 11278 26881 11324 26917
rect 11324 26881 11327 26917
rect 11275 26865 11327 26881
rect 11723 27347 11775 27353
rect 11723 27301 11726 27347
rect 11726 27301 11772 27347
rect 11772 27301 11775 27347
rect 11723 27091 11726 27135
rect 11726 27091 11772 27135
rect 11772 27091 11775 27135
rect 11723 27083 11775 27091
rect 11723 26881 11726 26917
rect 11726 26881 11772 26917
rect 11772 26881 11775 26917
rect 11723 26865 11775 26881
rect 12171 27347 12223 27353
rect 12171 27301 12174 27347
rect 12174 27301 12220 27347
rect 12220 27301 12223 27347
rect 12171 27091 12174 27135
rect 12174 27091 12220 27135
rect 12220 27091 12223 27135
rect 12171 27083 12223 27091
rect 12171 26881 12174 26917
rect 12174 26881 12220 26917
rect 12220 26881 12223 26917
rect 12171 26865 12223 26881
rect 12619 27347 12671 27353
rect 12619 27301 12622 27347
rect 12622 27301 12668 27347
rect 12668 27301 12671 27347
rect 12619 27091 12622 27135
rect 12622 27091 12668 27135
rect 12668 27091 12671 27135
rect 12619 27083 12671 27091
rect 13026 27326 13028 27378
rect 13028 27326 13074 27378
rect 13074 27326 13078 27378
rect 13026 27144 13028 27160
rect 13028 27144 13074 27160
rect 13074 27144 13078 27160
rect 13026 27108 13078 27144
rect 13302 27336 13312 27378
rect 13312 27336 13354 27378
rect 13302 27326 13354 27336
rect 13302 27132 13312 27160
rect 13312 27132 13354 27160
rect 13302 27108 13354 27132
rect 16157 27643 16209 27695
rect 17151 28030 17152 28041
rect 17152 28030 17198 28041
rect 17198 28030 17203 28041
rect 17151 27989 17203 28030
rect 16918 27925 16928 27956
rect 16928 27925 16970 27956
rect 16918 27904 16970 27925
rect 16918 27715 16928 27738
rect 16928 27715 16970 27738
rect 16918 27686 16970 27715
rect 12619 26881 12622 26917
rect 12622 26881 12668 26917
rect 12668 26881 12671 26917
rect 12619 26865 12671 26881
rect 14386 27158 14438 27210
rect 14598 27158 14650 27210
rect 15515 27378 15567 27392
rect 15515 27340 15520 27378
rect 15520 27340 15566 27378
rect 15566 27340 15567 27378
rect 16157 27425 16209 27477
rect 17828 28122 17880 28174
rect 17595 28030 17600 28041
rect 17600 28030 17646 28041
rect 17646 28030 17647 28041
rect 17595 27989 17647 28030
rect 17151 27820 17152 27823
rect 17152 27820 17198 27823
rect 17198 27820 17203 27823
rect 17151 27771 17203 27820
rect 17151 27553 17203 27605
rect 15515 27144 15520 27174
rect 15520 27144 15566 27174
rect 15566 27144 15567 27174
rect 15515 27122 15567 27144
rect 18552 28122 18604 28174
rect 17595 27820 17600 27823
rect 17600 27820 17646 27823
rect 17646 27820 17647 27823
rect 17595 27771 17647 27820
rect 17828 27925 17870 27956
rect 17870 27925 17880 27956
rect 17828 27904 17880 27925
rect 17828 27715 17870 27738
rect 17870 27715 17880 27738
rect 17828 27686 17880 27715
rect 17595 27553 17647 27605
rect 14384 26922 14436 26974
rect 14596 26922 14648 26974
rect 13253 26462 13305 26514
rect 13460 26462 13470 26514
rect 13470 26462 13512 26514
rect 13253 26244 13305 26296
rect 13460 26276 13470 26296
rect 13470 26276 13512 26296
rect 13460 26244 13512 26276
rect 13253 26026 13305 26078
rect 13460 26070 13470 26078
rect 13470 26070 13512 26078
rect 13460 26026 13512 26070
rect 13253 25808 13305 25860
rect 13460 25808 13512 25860
rect 13980 26446 14032 26491
rect 13980 26439 13984 26446
rect 13984 26439 14030 26446
rect 14030 26439 14032 26446
rect 14944 26462 14996 26514
rect 15151 26462 15161 26514
rect 15161 26462 15203 26514
rect 13980 26230 14032 26273
rect 13980 26221 13984 26230
rect 13984 26221 14030 26230
rect 14030 26221 14032 26230
rect 13980 26014 14032 26055
rect 13980 26003 13984 26014
rect 13984 26003 14030 26014
rect 14030 26003 14032 26014
rect 13980 25798 14032 25837
rect 13980 25785 13984 25798
rect 13984 25785 14030 25798
rect 14030 25785 14032 25798
rect 13253 25169 13305 25221
rect 13465 25218 13517 25221
rect 13465 25172 13491 25218
rect 13491 25172 13517 25218
rect 13465 25169 13517 25172
rect 8299 24759 8342 24811
rect 8342 24759 8351 24811
rect 8299 24541 8342 24593
rect 8342 24541 8351 24593
rect 8299 24324 8342 24376
rect 8342 24324 8351 24376
rect 8299 24106 8342 24158
rect 8342 24106 8351 24158
rect 8299 23888 8342 23940
rect 8342 23888 8351 23940
rect 8299 23670 8342 23722
rect 8342 23670 8351 23722
rect 8299 23453 8342 23505
rect 8342 23453 8351 23505
rect 8299 23267 8351 23287
rect 8299 23235 8342 23267
rect 8342 23235 8351 23267
rect 9196 24721 9248 24773
rect 9196 24550 9248 24556
rect 9196 24504 9242 24550
rect 9242 24504 9248 24550
rect 9196 24286 9242 24338
rect 9242 24286 9248 24338
rect 9196 24069 9242 24121
rect 9242 24069 9248 24121
rect 9196 23851 9242 23903
rect 9242 23851 9248 23903
rect 9196 23633 9242 23685
rect 9242 23633 9248 23685
rect 9196 23415 9242 23467
rect 9242 23415 9248 23467
rect 9196 23198 9242 23250
rect 9242 23198 9248 23250
rect 9196 22980 9242 23032
rect 9242 22980 9248 23032
rect 9196 22763 9242 22815
rect 9242 22763 9248 22815
rect 8516 22651 8568 22703
rect 8516 22443 8568 22485
rect 8516 22433 8520 22443
rect 8520 22433 8566 22443
rect 8566 22433 8568 22443
rect 9648 24721 9700 24773
rect 9931 24721 9983 24773
rect 10214 24721 10266 24773
rect 9648 24550 9700 24556
rect 8002 21744 8006 21796
rect 8006 21744 8052 21796
rect 8052 21744 8054 21796
rect 8002 21526 8006 21578
rect 8006 21526 8052 21578
rect 8052 21526 8054 21578
rect 9648 24504 9690 24550
rect 9690 24504 9700 24550
rect 9931 24504 9983 24556
rect 10214 24550 10266 24556
rect 10214 24504 10224 24550
rect 10224 24504 10266 24550
rect 9648 24286 9690 24338
rect 9690 24286 9700 24338
rect 9931 24286 9983 24338
rect 10214 24286 10224 24338
rect 10224 24286 10266 24338
rect 9648 24069 9690 24121
rect 9690 24069 9700 24121
rect 9931 24069 9983 24121
rect 10214 24069 10224 24121
rect 10224 24069 10266 24121
rect 9648 23851 9690 23903
rect 9690 23851 9700 23903
rect 9931 23851 9983 23903
rect 10214 23851 10224 23903
rect 10224 23851 10266 23903
rect 9648 23633 9690 23685
rect 9690 23633 9700 23685
rect 9931 23633 9983 23685
rect 10214 23633 10224 23685
rect 10224 23633 10266 23685
rect 9648 23415 9690 23467
rect 9690 23415 9700 23467
rect 9931 23415 9983 23467
rect 10214 23415 10224 23467
rect 10224 23415 10266 23467
rect 9648 23198 9690 23250
rect 9690 23198 9700 23250
rect 9931 23198 9983 23250
rect 10214 23198 10224 23250
rect 10224 23198 10266 23250
rect 9648 22980 9690 23032
rect 9690 22980 9700 23032
rect 9931 22980 9983 23032
rect 10214 22980 10224 23032
rect 10224 22980 10266 23032
rect 9648 22763 9690 22815
rect 9690 22763 9700 22815
rect 9931 22763 9983 22815
rect 10214 22763 10224 22815
rect 10224 22763 10266 22815
rect 9418 21790 9470 21842
rect 9418 21582 9470 21624
rect 9418 21572 9420 21582
rect 9420 21572 9466 21582
rect 9466 21572 9470 21582
rect 10666 24721 10718 24773
rect 10666 24550 10718 24556
rect 10666 24504 10672 24550
rect 10672 24504 10718 24550
rect 10666 24286 10672 24338
rect 10672 24286 10718 24338
rect 10666 24069 10672 24121
rect 10672 24069 10718 24121
rect 10666 23851 10672 23903
rect 10672 23851 10718 23903
rect 10666 23633 10672 23685
rect 10672 23633 10718 23685
rect 10666 23415 10672 23467
rect 10672 23415 10718 23467
rect 10666 23198 10672 23250
rect 10672 23198 10718 23250
rect 10666 22980 10672 23032
rect 10672 22980 10718 23032
rect 10666 22763 10672 22815
rect 10672 22763 10718 22815
rect 10988 24721 11040 24773
rect 10988 24550 11040 24556
rect 10988 24504 11034 24550
rect 11034 24504 11040 24550
rect 10988 24286 11034 24338
rect 11034 24286 11040 24338
rect 10988 24069 11034 24121
rect 11034 24069 11040 24121
rect 10988 23851 11034 23903
rect 11034 23851 11040 23903
rect 10988 23633 11034 23685
rect 11034 23633 11040 23685
rect 10988 23415 11034 23467
rect 11034 23415 11040 23467
rect 10988 23198 11034 23250
rect 11034 23198 11040 23250
rect 10988 22980 11034 23032
rect 11034 22980 11040 23032
rect 10988 22763 11034 22815
rect 11034 22763 11040 22815
rect 10444 21790 10496 21842
rect 10444 21582 10496 21624
rect 10444 21572 10448 21582
rect 10448 21572 10494 21582
rect 10494 21572 10496 21582
rect 11440 24721 11492 24773
rect 11723 24721 11775 24773
rect 12006 24721 12058 24773
rect 11440 24550 11492 24556
rect 11440 24504 11482 24550
rect 11482 24504 11492 24550
rect 11723 24504 11775 24556
rect 12006 24550 12058 24556
rect 12006 24504 12016 24550
rect 12016 24504 12058 24550
rect 11440 24286 11482 24338
rect 11482 24286 11492 24338
rect 11723 24286 11775 24338
rect 12006 24286 12016 24338
rect 12016 24286 12058 24338
rect 11440 24069 11482 24121
rect 11482 24069 11492 24121
rect 11723 24069 11775 24121
rect 12006 24069 12016 24121
rect 12016 24069 12058 24121
rect 11440 23851 11482 23903
rect 11482 23851 11492 23903
rect 11723 23851 11775 23903
rect 12006 23851 12016 23903
rect 12016 23851 12058 23903
rect 11440 23633 11482 23685
rect 11482 23633 11492 23685
rect 11723 23633 11775 23685
rect 12006 23633 12016 23685
rect 12016 23633 12058 23685
rect 11440 23415 11482 23467
rect 11482 23415 11492 23467
rect 11723 23415 11775 23467
rect 12006 23415 12016 23467
rect 12016 23415 12058 23467
rect 11440 23198 11482 23250
rect 11482 23198 11492 23250
rect 11723 23198 11775 23250
rect 12006 23198 12016 23250
rect 12016 23198 12058 23250
rect 11440 22980 11482 23032
rect 11482 22980 11492 23032
rect 11723 22980 11775 23032
rect 12006 22980 12016 23032
rect 12016 22980 12058 23032
rect 11440 22763 11482 22815
rect 11482 22763 11492 22815
rect 11723 22763 11775 22815
rect 12006 22763 12016 22815
rect 12016 22763 12058 22815
rect 11210 21790 11262 21842
rect 11210 21582 11262 21624
rect 11210 21572 11212 21582
rect 11212 21572 11258 21582
rect 11258 21572 11262 21582
rect 12458 24721 12510 24773
rect 12458 24550 12510 24556
rect 12458 24504 12464 24550
rect 12464 24504 12510 24550
rect 12458 24286 12464 24338
rect 12464 24286 12510 24338
rect 12458 24069 12464 24121
rect 12464 24069 12510 24121
rect 12458 23851 12464 23903
rect 12464 23851 12510 23903
rect 12458 23633 12464 23685
rect 12464 23633 12510 23685
rect 12458 23415 12464 23467
rect 12464 23415 12510 23467
rect 12458 23198 12464 23250
rect 12464 23198 12510 23250
rect 12458 22980 12464 23032
rect 12464 22980 12510 23032
rect 12458 22763 12464 22815
rect 12464 22763 12510 22815
rect 13473 24750 13516 24802
rect 13516 24750 13525 24802
rect 13473 24533 13516 24585
rect 13516 24533 13525 24585
rect 13473 24315 13516 24367
rect 13516 24315 13525 24367
rect 13473 24098 13516 24150
rect 13516 24098 13525 24150
rect 13473 23880 13516 23932
rect 13516 23880 13525 23932
rect 13473 23662 13516 23714
rect 13516 23662 13525 23714
rect 13473 23444 13516 23496
rect 13516 23444 13525 23496
rect 13473 23227 13516 23279
rect 13516 23227 13525 23279
rect 13473 23009 13516 23061
rect 13516 23009 13525 23061
rect 13473 22792 13516 22844
rect 13516 22792 13525 22844
rect 12236 21790 12288 21842
rect 12236 21582 12288 21624
rect 12236 21572 12240 21582
rect 12240 21572 12286 21582
rect 12286 21572 12288 21582
rect 14944 26244 14996 26296
rect 15151 26276 15161 26296
rect 15161 26276 15203 26296
rect 15151 26244 15203 26276
rect 14944 26026 14996 26078
rect 15151 26070 15161 26078
rect 15161 26070 15203 26078
rect 15151 26026 15203 26070
rect 14944 25808 14996 25860
rect 15151 25808 15203 25860
rect 15671 26446 15723 26491
rect 15671 26439 15675 26446
rect 15675 26439 15721 26446
rect 15721 26439 15723 26446
rect 15671 26230 15723 26273
rect 15671 26221 15675 26230
rect 15675 26221 15721 26230
rect 15721 26221 15723 26230
rect 15671 26014 15723 26055
rect 15671 26003 15675 26014
rect 15675 26003 15721 26014
rect 15721 26003 15723 26014
rect 15671 25798 15723 25837
rect 15671 25785 15675 25798
rect 15675 25785 15721 25798
rect 15721 25785 15723 25798
rect 14944 25169 14996 25221
rect 15156 25218 15208 25221
rect 15156 25172 15182 25218
rect 15182 25172 15208 25218
rect 15156 25169 15208 25172
rect 13987 24759 14030 24811
rect 14030 24759 14039 24811
rect 13987 24541 14030 24593
rect 14030 24541 14039 24593
rect 13987 24324 14030 24376
rect 14030 24324 14039 24376
rect 13987 24106 14030 24158
rect 14030 24106 14039 24158
rect 13987 23888 14030 23940
rect 14030 23888 14039 23940
rect 13987 23670 14030 23722
rect 14030 23670 14039 23722
rect 13987 23453 14030 23505
rect 14030 23453 14039 23505
rect 13987 23267 14039 23287
rect 13987 23235 14030 23267
rect 14030 23235 14039 23267
rect 15164 24750 15207 24802
rect 15207 24750 15216 24802
rect 15164 24533 15207 24585
rect 15207 24533 15216 24585
rect 15164 24315 15207 24367
rect 15207 24315 15216 24367
rect 15164 24098 15207 24150
rect 15207 24098 15216 24150
rect 15164 23880 15207 23932
rect 15207 23880 15216 23932
rect 15164 23662 15207 23714
rect 15207 23662 15216 23714
rect 15164 23444 15207 23496
rect 15207 23444 15216 23496
rect 15164 23227 15207 23279
rect 15207 23227 15216 23279
rect 15164 23009 15207 23061
rect 15207 23009 15216 23061
rect 14204 22651 14256 22703
rect 14204 22443 14256 22485
rect 14204 22433 14208 22443
rect 14208 22433 14254 22443
rect 14254 22433 14256 22443
rect 15164 22792 15207 22844
rect 15207 22792 15216 22844
rect 13690 21744 13694 21796
rect 13694 21744 13740 21796
rect 13740 21744 13742 21796
rect 13690 21526 13694 21578
rect 13694 21526 13740 21578
rect 13740 21526 13742 21578
rect 15678 24759 15721 24811
rect 15721 24759 15730 24811
rect 15678 24541 15721 24593
rect 15721 24541 15730 24593
rect 15678 24324 15721 24376
rect 15721 24324 15730 24376
rect 15678 24106 15721 24158
rect 15721 24106 15730 24158
rect 15678 23888 15721 23940
rect 15721 23888 15730 23940
rect 15678 23670 15721 23722
rect 15721 23670 15730 23722
rect 15678 23453 15721 23505
rect 15721 23453 15730 23505
rect 15678 23267 15730 23287
rect 15678 23235 15721 23267
rect 15721 23235 15730 23267
rect 18785 28030 18786 28041
rect 18786 28030 18832 28041
rect 18832 28030 18837 28041
rect 18785 27989 18837 28030
rect 18552 27925 18562 27956
rect 18562 27925 18604 27956
rect 18552 27904 18604 27925
rect 18552 27715 18562 27738
rect 18562 27715 18604 27738
rect 18552 27686 18604 27715
rect 19462 28122 19514 28174
rect 19229 28030 19234 28041
rect 19234 28030 19280 28041
rect 19280 28030 19281 28041
rect 19229 27989 19281 28030
rect 18785 27820 18786 27823
rect 18786 27820 18832 27823
rect 18832 27820 18837 27823
rect 18785 27771 18837 27820
rect 18785 27553 18837 27605
rect 16925 25270 16928 25300
rect 16928 25270 16974 25300
rect 16974 25270 16977 25300
rect 16925 25248 16977 25270
rect 16925 25062 16928 25082
rect 16928 25062 16974 25082
rect 16974 25062 16977 25082
rect 16925 25030 16977 25062
rect 16925 24854 16928 24864
rect 16928 24854 16974 24864
rect 16974 24854 16977 24864
rect 16925 24812 16977 24854
rect 17373 25270 17376 25300
rect 17376 25270 17422 25300
rect 17422 25270 17425 25300
rect 17373 25248 17425 25270
rect 17373 25062 17376 25082
rect 17376 25062 17422 25082
rect 17422 25062 17425 25082
rect 17373 25030 17425 25062
rect 17373 24854 17376 24864
rect 17376 24854 17422 24864
rect 17422 24854 17425 24864
rect 17373 24812 17425 24854
rect 20185 28122 20237 28174
rect 19229 27820 19234 27823
rect 19234 27820 19280 27823
rect 19280 27820 19281 27823
rect 19229 27771 19281 27820
rect 19462 27925 19504 27956
rect 19504 27925 19514 27956
rect 19462 27904 19514 27925
rect 19462 27715 19504 27738
rect 19504 27715 19514 27738
rect 19462 27686 19514 27715
rect 19229 27553 19281 27605
rect 17821 25270 17824 25300
rect 17824 25270 17870 25300
rect 17870 25270 17873 25300
rect 17821 25248 17873 25270
rect 17821 25062 17824 25082
rect 17824 25062 17870 25082
rect 17870 25062 17873 25082
rect 17821 25030 17873 25062
rect 17821 24854 17824 24864
rect 17824 24854 17870 24864
rect 17870 24854 17873 24864
rect 17821 24812 17873 24854
rect 20418 28030 20419 28041
rect 20419 28030 20465 28041
rect 20465 28030 20470 28041
rect 20418 27989 20470 28030
rect 20185 27925 20195 27956
rect 20195 27925 20237 27956
rect 20185 27904 20237 27925
rect 20185 27715 20195 27738
rect 20195 27715 20237 27738
rect 20185 27686 20237 27715
rect 21095 28122 21147 28174
rect 20862 28030 20867 28041
rect 20867 28030 20913 28041
rect 20913 28030 20914 28041
rect 20862 27989 20914 28030
rect 20418 27820 20419 27823
rect 20419 27820 20465 27823
rect 20465 27820 20470 27823
rect 20418 27771 20470 27820
rect 20418 27553 20470 27605
rect 18559 25270 18562 25300
rect 18562 25270 18608 25300
rect 18608 25270 18611 25300
rect 18559 25248 18611 25270
rect 18559 25062 18562 25082
rect 18562 25062 18608 25082
rect 18608 25062 18611 25082
rect 18559 25030 18611 25062
rect 18559 24854 18562 24864
rect 18562 24854 18608 24864
rect 18608 24854 18611 24864
rect 18559 24812 18611 24854
rect 19007 25270 19010 25300
rect 19010 25270 19056 25300
rect 19056 25270 19059 25300
rect 19007 25248 19059 25270
rect 19007 25062 19010 25082
rect 19010 25062 19056 25082
rect 19056 25062 19059 25082
rect 19007 25030 19059 25062
rect 19007 24854 19010 24864
rect 19010 24854 19056 24864
rect 19056 24854 19059 24864
rect 19007 24812 19059 24854
rect 21819 28122 21871 28174
rect 20862 27820 20867 27823
rect 20867 27820 20913 27823
rect 20913 27820 20914 27823
rect 20862 27771 20914 27820
rect 21095 27925 21137 27956
rect 21137 27925 21147 27956
rect 21095 27904 21147 27925
rect 21095 27715 21137 27738
rect 21137 27715 21147 27738
rect 21095 27686 21147 27715
rect 20862 27553 20914 27605
rect 19455 25270 19458 25300
rect 19458 25270 19504 25300
rect 19504 25270 19507 25300
rect 19455 25248 19507 25270
rect 19455 25062 19458 25082
rect 19458 25062 19504 25082
rect 19504 25062 19507 25082
rect 19455 25030 19507 25062
rect 19455 24854 19458 24864
rect 19458 24854 19504 24864
rect 19504 24854 19507 24864
rect 19455 24812 19507 24854
rect 22052 28030 22053 28041
rect 22053 28030 22099 28041
rect 22099 28030 22104 28041
rect 22052 27989 22104 28030
rect 21819 27925 21829 27956
rect 21829 27925 21871 27956
rect 21819 27904 21871 27925
rect 21819 27715 21829 27738
rect 21829 27715 21871 27738
rect 21819 27686 21871 27715
rect 22729 28122 22781 28174
rect 22496 28030 22501 28041
rect 22501 28030 22547 28041
rect 22547 28030 22548 28041
rect 22496 27989 22548 28030
rect 22052 27820 22053 27823
rect 22053 27820 22099 27823
rect 22099 27820 22104 27823
rect 22052 27771 22104 27820
rect 22052 27553 22104 27605
rect 20192 25270 20195 25300
rect 20195 25270 20241 25300
rect 20241 25270 20244 25300
rect 20192 25248 20244 25270
rect 20192 25062 20195 25082
rect 20195 25062 20241 25082
rect 20241 25062 20244 25082
rect 20192 25030 20244 25062
rect 20192 24854 20195 24864
rect 20195 24854 20241 24864
rect 20241 24854 20244 24864
rect 20192 24812 20244 24854
rect 20640 25270 20643 25300
rect 20643 25270 20689 25300
rect 20689 25270 20692 25300
rect 20640 25248 20692 25270
rect 20640 25062 20643 25082
rect 20643 25062 20689 25082
rect 20689 25062 20692 25082
rect 20640 25030 20692 25062
rect 20640 24854 20643 24864
rect 20643 24854 20689 24864
rect 20689 24854 20692 24864
rect 20640 24812 20692 24854
rect 23787 28144 23797 28183
rect 23797 28144 23839 28183
rect 23787 28131 23839 28144
rect 25610 28292 25662 28344
rect 22496 27820 22501 27823
rect 22501 27820 22547 27823
rect 22547 27820 22548 27823
rect 22496 27771 22548 27820
rect 22729 27925 22771 27956
rect 22771 27925 22781 27956
rect 22729 27904 22781 27925
rect 22729 27715 22771 27738
rect 22771 27715 22781 27738
rect 22729 27686 22781 27715
rect 22496 27553 22548 27605
rect 23787 27938 23797 27965
rect 23797 27938 23839 27965
rect 23787 27913 23839 27938
rect 24226 28144 24245 28183
rect 24245 28144 24278 28183
rect 24226 28131 24278 28144
rect 24226 27938 24245 27965
rect 24245 27938 24278 27965
rect 24226 27913 24278 27938
rect 21088 25270 21091 25300
rect 21091 25270 21137 25300
rect 21137 25270 21140 25300
rect 21088 25248 21140 25270
rect 21088 25062 21091 25082
rect 21091 25062 21137 25082
rect 21137 25062 21140 25082
rect 21088 25030 21140 25062
rect 21088 24854 21091 24864
rect 21091 24854 21137 24864
rect 21137 24854 21140 24864
rect 21088 24812 21140 24854
rect 23598 27643 23650 27695
rect 23810 27694 23862 27695
rect 23810 27648 23819 27694
rect 23819 27648 23862 27694
rect 23810 27643 23862 27648
rect 24446 28133 24498 28185
rect 24446 27915 24469 27967
rect 24469 27915 24498 27967
rect 25610 28076 25662 28126
rect 25610 28074 25616 28076
rect 25616 28074 25662 28076
rect 25610 27856 25616 27908
rect 25616 27856 25662 27908
rect 23787 27336 23797 27378
rect 23797 27336 23839 27378
rect 23787 27326 23839 27336
rect 23787 27132 23797 27160
rect 23797 27132 23839 27160
rect 23787 27108 23839 27132
rect 24572 27666 24728 27673
rect 24572 27621 24683 27666
rect 24683 27621 24728 27666
rect 26642 27634 26694 27686
rect 21826 25270 21829 25300
rect 21829 25270 21875 25300
rect 21875 25270 21878 25300
rect 21826 25248 21878 25270
rect 21826 25062 21829 25082
rect 21829 25062 21875 25082
rect 21875 25062 21878 25082
rect 21826 25030 21878 25062
rect 21826 24854 21829 24864
rect 21829 24854 21875 24864
rect 21875 24854 21878 24864
rect 21826 24812 21878 24854
rect 22274 25270 22277 25300
rect 22277 25270 22323 25300
rect 22323 25270 22326 25300
rect 22274 25248 22326 25270
rect 22274 25062 22277 25082
rect 22277 25062 22323 25082
rect 22323 25062 22326 25082
rect 22274 25030 22326 25062
rect 22274 24854 22277 24864
rect 22277 24854 22323 24864
rect 22323 24854 22326 24864
rect 22274 24812 22326 24854
rect 24973 27385 25025 27437
rect 24973 27167 25025 27219
rect 26001 27340 26053 27392
rect 26642 27416 26694 27468
rect 26001 27122 26053 27174
rect 24869 26922 24921 26974
rect 25081 26922 25133 26974
rect 23739 26483 23791 26535
rect 23946 26524 23998 26535
rect 23946 26483 23956 26524
rect 23956 26483 23998 26524
rect 23739 26265 23791 26317
rect 23946 26272 23956 26317
rect 23956 26272 23998 26317
rect 23946 26265 23998 26272
rect 23739 26047 23791 26099
rect 23946 26064 23956 26099
rect 23956 26064 23998 26099
rect 23946 26047 23998 26064
rect 23739 25829 23791 25881
rect 23946 25856 23956 25881
rect 23956 25856 23998 25881
rect 23946 25829 23998 25856
rect 24466 26524 24518 26535
rect 24466 26483 24470 26524
rect 24470 26483 24516 26524
rect 24516 26483 24518 26524
rect 24466 26272 24470 26317
rect 24470 26272 24516 26317
rect 24516 26272 24518 26317
rect 24466 26265 24518 26272
rect 24466 26064 24470 26099
rect 24470 26064 24516 26099
rect 24516 26064 24518 26099
rect 24466 26047 24518 26064
rect 24466 25856 24470 25881
rect 24470 25856 24516 25881
rect 24516 25856 24518 25881
rect 24466 25829 24518 25856
rect 22722 25270 22725 25300
rect 22725 25270 22771 25300
rect 22771 25270 22774 25300
rect 22722 25248 22774 25270
rect 22722 25062 22725 25082
rect 22725 25062 22771 25082
rect 22771 25062 22774 25082
rect 22722 25030 22774 25062
rect 22722 24854 22725 24864
rect 22725 24854 22771 24864
rect 22771 24854 22774 24864
rect 22722 24812 22774 24854
rect 25429 26483 25481 26535
rect 25636 26524 25688 26535
rect 25636 26483 25646 26524
rect 25646 26483 25688 26524
rect 25429 26265 25481 26317
rect 25636 26272 25646 26317
rect 25646 26272 25688 26317
rect 25636 26265 25688 26272
rect 25429 26047 25481 26099
rect 25636 26064 25646 26099
rect 25646 26064 25688 26099
rect 25636 26047 25688 26064
rect 25429 25829 25481 25881
rect 25636 25856 25646 25881
rect 25646 25856 25688 25881
rect 25636 25829 25688 25856
rect 23739 25260 23791 25312
rect 23951 25309 24003 25312
rect 23951 25263 23977 25309
rect 23977 25263 24003 25309
rect 23951 25260 24003 25263
rect 23959 24985 24002 24997
rect 24002 24985 24011 24997
rect 23959 24945 24011 24985
rect 23959 24779 24002 24780
rect 24002 24779 24011 24780
rect 23959 24728 24011 24779
rect 15895 22651 15947 22703
rect 15895 22443 15947 22485
rect 15895 22433 15899 22443
rect 15899 22433 15945 22443
rect 15945 22433 15947 22443
rect 16929 24128 16981 24180
rect 17373 24128 17425 24180
rect 16929 23910 16974 23962
rect 16974 23910 16981 23962
rect 16929 23693 16974 23745
rect 16974 23693 16981 23745
rect 16929 23475 16974 23527
rect 16974 23475 16981 23527
rect 16929 23257 16974 23309
rect 16974 23257 16981 23309
rect 16929 23040 16974 23092
rect 16974 23040 16981 23092
rect 16929 22822 16974 22874
rect 16974 22822 16981 22874
rect 16701 22178 16704 22230
rect 16704 22178 16750 22230
rect 16750 22178 16753 22230
rect 16701 21960 16704 22012
rect 16704 21960 16750 22012
rect 16750 21960 16753 22012
rect 17817 24128 17869 24180
rect 17373 23910 17376 23962
rect 17376 23910 17422 23962
rect 17422 23910 17425 23962
rect 17373 23693 17376 23745
rect 17376 23693 17422 23745
rect 17422 23693 17425 23745
rect 17373 23475 17376 23527
rect 17376 23475 17422 23527
rect 17422 23475 17425 23527
rect 17373 23257 17376 23309
rect 17376 23257 17422 23309
rect 17422 23257 17425 23309
rect 17373 23040 17376 23092
rect 17376 23040 17422 23092
rect 17422 23040 17425 23092
rect 17373 22822 17376 22874
rect 17376 22822 17422 22874
rect 17422 22822 17425 22874
rect 17149 22178 17152 22230
rect 17152 22178 17198 22230
rect 17198 22178 17201 22230
rect 17149 21960 17152 22012
rect 17152 21960 17198 22012
rect 17198 21960 17201 22012
rect 17817 23910 17824 23962
rect 17824 23910 17869 23962
rect 17817 23693 17824 23745
rect 17824 23693 17869 23745
rect 17817 23475 17824 23527
rect 17824 23475 17869 23527
rect 17817 23257 17824 23309
rect 17824 23257 17869 23309
rect 17817 23040 17824 23092
rect 17824 23040 17869 23092
rect 17817 22822 17824 22874
rect 17824 22822 17869 22874
rect 17597 22178 17600 22230
rect 17600 22178 17646 22230
rect 17646 22178 17649 22230
rect 17597 21960 17600 22012
rect 17600 21960 17646 22012
rect 17646 21960 17649 22012
rect 18045 22178 18048 22230
rect 18048 22178 18094 22230
rect 18094 22178 18097 22230
rect 18045 21960 18048 22012
rect 18048 21960 18094 22012
rect 18094 21960 18097 22012
rect 18563 24128 18615 24180
rect 19007 24128 19059 24180
rect 18563 23910 18608 23962
rect 18608 23910 18615 23962
rect 18563 23693 18608 23745
rect 18608 23693 18615 23745
rect 18563 23475 18608 23527
rect 18608 23475 18615 23527
rect 18563 23257 18608 23309
rect 18608 23257 18615 23309
rect 18563 23040 18608 23092
rect 18608 23040 18615 23092
rect 18563 22822 18608 22874
rect 18608 22822 18615 22874
rect 18335 22178 18338 22230
rect 18338 22178 18384 22230
rect 18384 22178 18387 22230
rect 18335 21960 18338 22012
rect 18338 21960 18384 22012
rect 18384 21960 18387 22012
rect 19451 24128 19503 24180
rect 19007 23910 19010 23962
rect 19010 23910 19056 23962
rect 19056 23910 19059 23962
rect 19007 23693 19010 23745
rect 19010 23693 19056 23745
rect 19056 23693 19059 23745
rect 19007 23475 19010 23527
rect 19010 23475 19056 23527
rect 19056 23475 19059 23527
rect 19007 23257 19010 23309
rect 19010 23257 19056 23309
rect 19056 23257 19059 23309
rect 19007 23040 19010 23092
rect 19010 23040 19056 23092
rect 19056 23040 19059 23092
rect 19007 22822 19010 22874
rect 19010 22822 19056 22874
rect 19056 22822 19059 22874
rect 18783 22178 18786 22230
rect 18786 22178 18832 22230
rect 18832 22178 18835 22230
rect 18783 21960 18786 22012
rect 18786 21960 18832 22012
rect 18832 21960 18835 22012
rect 19451 23910 19458 23962
rect 19458 23910 19503 23962
rect 19451 23693 19458 23745
rect 19458 23693 19503 23745
rect 19451 23475 19458 23527
rect 19458 23475 19503 23527
rect 19451 23257 19458 23309
rect 19458 23257 19503 23309
rect 19451 23040 19458 23092
rect 19458 23040 19503 23092
rect 19451 22822 19458 22874
rect 19458 22822 19503 22874
rect 19231 22178 19234 22230
rect 19234 22178 19280 22230
rect 19280 22178 19283 22230
rect 19231 21960 19234 22012
rect 19234 21960 19280 22012
rect 19280 21960 19283 22012
rect 19679 22178 19682 22230
rect 19682 22178 19728 22230
rect 19728 22178 19731 22230
rect 19679 21960 19682 22012
rect 19682 21960 19728 22012
rect 19728 21960 19731 22012
rect 20196 24128 20248 24180
rect 20640 24128 20692 24180
rect 20196 23910 20241 23962
rect 20241 23910 20248 23962
rect 20196 23693 20241 23745
rect 20241 23693 20248 23745
rect 20196 23475 20241 23527
rect 20241 23475 20248 23527
rect 20196 23257 20241 23309
rect 20241 23257 20248 23309
rect 20196 23040 20241 23092
rect 20241 23040 20248 23092
rect 20196 22822 20241 22874
rect 20241 22822 20248 22874
rect 19968 22178 19971 22230
rect 19971 22178 20017 22230
rect 20017 22178 20020 22230
rect 19968 21960 19971 22012
rect 19971 21960 20017 22012
rect 20017 21960 20020 22012
rect 21084 24128 21136 24180
rect 20640 23910 20643 23962
rect 20643 23910 20689 23962
rect 20689 23910 20692 23962
rect 20640 23693 20643 23745
rect 20643 23693 20689 23745
rect 20689 23693 20692 23745
rect 20640 23475 20643 23527
rect 20643 23475 20689 23527
rect 20689 23475 20692 23527
rect 20640 23257 20643 23309
rect 20643 23257 20689 23309
rect 20689 23257 20692 23309
rect 20640 23040 20643 23092
rect 20643 23040 20689 23092
rect 20689 23040 20692 23092
rect 20640 22822 20643 22874
rect 20643 22822 20689 22874
rect 20689 22822 20692 22874
rect 20416 22178 20419 22230
rect 20419 22178 20465 22230
rect 20465 22178 20468 22230
rect 20416 21960 20419 22012
rect 20419 21960 20465 22012
rect 20465 21960 20468 22012
rect 21084 23910 21091 23962
rect 21091 23910 21136 23962
rect 21084 23693 21091 23745
rect 21091 23693 21136 23745
rect 21084 23475 21091 23527
rect 21091 23475 21136 23527
rect 21084 23257 21091 23309
rect 21091 23257 21136 23309
rect 21084 23040 21091 23092
rect 21091 23040 21136 23092
rect 21084 22822 21091 22874
rect 21091 22822 21136 22874
rect 20864 22178 20867 22230
rect 20867 22178 20913 22230
rect 20913 22178 20916 22230
rect 20864 21960 20867 22012
rect 20867 21960 20913 22012
rect 20913 21960 20916 22012
rect 21312 22178 21315 22230
rect 21315 22178 21361 22230
rect 21361 22178 21364 22230
rect 21312 21960 21315 22012
rect 21315 21960 21361 22012
rect 21361 21960 21364 22012
rect 21830 24128 21882 24180
rect 22274 24128 22326 24180
rect 21830 23910 21875 23962
rect 21875 23910 21882 23962
rect 21830 23693 21875 23745
rect 21875 23693 21882 23745
rect 21830 23475 21875 23527
rect 21875 23475 21882 23527
rect 21830 23257 21875 23309
rect 21875 23257 21882 23309
rect 21830 23040 21875 23092
rect 21875 23040 21882 23092
rect 21830 22822 21875 22874
rect 21875 22822 21882 22874
rect 21602 22178 21605 22230
rect 21605 22178 21651 22230
rect 21651 22178 21654 22230
rect 21602 21960 21605 22012
rect 21605 21960 21651 22012
rect 21651 21960 21654 22012
rect 22718 24128 22770 24180
rect 22274 23910 22277 23962
rect 22277 23910 22323 23962
rect 22323 23910 22326 23962
rect 22274 23693 22277 23745
rect 22277 23693 22323 23745
rect 22323 23693 22326 23745
rect 22274 23475 22277 23527
rect 22277 23475 22323 23527
rect 22323 23475 22326 23527
rect 22274 23257 22277 23309
rect 22277 23257 22323 23309
rect 22323 23257 22326 23309
rect 22274 23040 22277 23092
rect 22277 23040 22323 23092
rect 22323 23040 22326 23092
rect 22274 22822 22277 22874
rect 22277 22822 22323 22874
rect 22323 22822 22326 22874
rect 22050 22178 22053 22230
rect 22053 22178 22099 22230
rect 22099 22178 22102 22230
rect 22050 21960 22053 22012
rect 22053 21960 22099 22012
rect 22099 21960 22102 22012
rect 22718 23910 22725 23962
rect 22725 23910 22770 23962
rect 22718 23693 22725 23745
rect 22725 23693 22770 23745
rect 22718 23475 22725 23527
rect 22725 23475 22770 23527
rect 22718 23257 22725 23309
rect 22725 23257 22770 23309
rect 22718 23040 22725 23092
rect 22725 23040 22770 23092
rect 22718 22822 22725 22874
rect 22725 22822 22770 22874
rect 22498 22178 22501 22230
rect 22501 22178 22547 22230
rect 22547 22178 22550 22230
rect 22498 21960 22501 22012
rect 22501 21960 22547 22012
rect 22547 21960 22550 22012
rect 23959 24516 24011 24562
rect 23959 24510 24002 24516
rect 24002 24510 24011 24516
rect 23959 24310 24011 24344
rect 23959 24292 24002 24310
rect 24002 24292 24011 24310
rect 23959 24104 24011 24126
rect 23959 24074 24002 24104
rect 24002 24074 24011 24104
rect 23959 23898 24011 23909
rect 23959 23857 24002 23898
rect 24002 23857 24011 23898
rect 26156 26524 26208 26535
rect 26156 26483 26160 26524
rect 26160 26483 26206 26524
rect 26206 26483 26208 26524
rect 26156 26272 26160 26317
rect 26160 26272 26206 26317
rect 26206 26272 26208 26317
rect 26156 26265 26208 26272
rect 26156 26064 26160 26099
rect 26160 26064 26206 26099
rect 26206 26064 26208 26099
rect 26156 26047 26208 26064
rect 26156 25856 26160 25881
rect 26160 25856 26206 25881
rect 26206 25856 26208 25881
rect 26156 25829 26208 25856
rect 27120 26483 27172 26535
rect 27327 26524 27379 26535
rect 27327 26483 27337 26524
rect 27337 26483 27379 26524
rect 27120 26265 27172 26317
rect 27327 26272 27337 26317
rect 27337 26272 27379 26317
rect 27327 26265 27379 26272
rect 27120 26047 27172 26099
rect 27327 26064 27337 26099
rect 27337 26064 27379 26099
rect 27327 26047 27379 26064
rect 27120 25829 27172 25881
rect 27327 25856 27337 25881
rect 27337 25856 27379 25881
rect 27327 25829 27379 25856
rect 25429 25260 25481 25312
rect 25641 25309 25693 25312
rect 25641 25263 25667 25309
rect 25667 25263 25693 25309
rect 25641 25260 25693 25263
rect 22946 22178 22949 22230
rect 22949 22178 22995 22230
rect 22995 22178 22998 22230
rect 22946 21960 22949 22012
rect 22949 21960 22995 22012
rect 22995 21960 22998 22012
rect 24473 24985 24516 24997
rect 24516 24985 24525 24997
rect 24473 24945 24525 24985
rect 24473 24779 24516 24780
rect 24516 24779 24525 24780
rect 24473 24728 24525 24779
rect 24473 24516 24525 24562
rect 24473 24510 24516 24516
rect 24516 24510 24525 24516
rect 24473 24310 24525 24344
rect 24473 24292 24516 24310
rect 24516 24292 24525 24310
rect 24473 24104 24525 24126
rect 24473 24074 24516 24104
rect 24516 24074 24525 24104
rect 24473 23898 24525 23909
rect 24473 23857 24516 23898
rect 24516 23857 24525 23898
rect 25649 24985 25692 24997
rect 25692 24985 25701 24997
rect 25649 24945 25701 24985
rect 24176 22148 24228 22200
rect 24176 21940 24228 21982
rect 24176 21930 24180 21940
rect 24180 21930 24226 21940
rect 24226 21930 24228 21940
rect 15381 21744 15385 21796
rect 15385 21744 15431 21796
rect 15431 21744 15433 21796
rect 25649 24779 25692 24780
rect 25692 24779 25701 24780
rect 25649 24728 25701 24779
rect 25649 24516 25701 24562
rect 25649 24510 25692 24516
rect 25692 24510 25701 24516
rect 25649 24310 25701 24344
rect 25649 24292 25692 24310
rect 25692 24292 25701 24310
rect 25649 24104 25701 24126
rect 25649 24074 25692 24104
rect 25692 24074 25701 24104
rect 25649 23898 25701 23909
rect 25649 23857 25692 23898
rect 25692 23857 25701 23898
rect 27847 26524 27899 26535
rect 27847 26483 27851 26524
rect 27851 26483 27897 26524
rect 27897 26483 27899 26524
rect 27847 26272 27851 26317
rect 27851 26272 27897 26317
rect 27897 26272 27899 26317
rect 27847 26265 27899 26272
rect 27847 26064 27851 26099
rect 27851 26064 27897 26099
rect 27897 26064 27899 26099
rect 27847 26047 27899 26064
rect 27847 25856 27851 25881
rect 27851 25856 27897 25881
rect 27897 25856 27899 25881
rect 27847 25829 27899 25856
rect 27120 25260 27172 25312
rect 27332 25309 27384 25312
rect 27332 25263 27358 25309
rect 27358 25263 27384 25309
rect 27332 25260 27384 25263
rect 24690 22148 24742 22200
rect 24690 21940 24742 21982
rect 24690 21930 24694 21940
rect 24694 21930 24740 21940
rect 24740 21930 24742 21940
rect 26163 24985 26206 24997
rect 26206 24985 26215 24997
rect 26163 24945 26215 24985
rect 26163 24779 26206 24780
rect 26206 24779 26215 24780
rect 26163 24728 26215 24779
rect 26163 24516 26215 24562
rect 26163 24510 26206 24516
rect 26206 24510 26215 24516
rect 26163 24310 26215 24344
rect 26163 24292 26206 24310
rect 26206 24292 26215 24310
rect 26163 24104 26215 24126
rect 26163 24074 26206 24104
rect 26206 24074 26215 24104
rect 26163 23898 26215 23909
rect 26163 23857 26206 23898
rect 26206 23857 26215 23898
rect 27340 24985 27383 24997
rect 27383 24985 27392 24997
rect 27340 24945 27392 24985
rect 25866 22148 25918 22200
rect 25866 21940 25918 21982
rect 25866 21930 25870 21940
rect 25870 21930 25916 21940
rect 25916 21930 25918 21940
rect 27340 24779 27383 24780
rect 27383 24779 27392 24780
rect 27340 24728 27392 24779
rect 27340 24516 27392 24562
rect 27340 24510 27383 24516
rect 27383 24510 27392 24516
rect 27340 24310 27392 24344
rect 27340 24292 27383 24310
rect 27383 24292 27392 24310
rect 27340 24104 27392 24126
rect 27340 24074 27383 24104
rect 27383 24074 27392 24104
rect 27340 23898 27392 23909
rect 27340 23857 27383 23898
rect 27383 23857 27392 23898
rect 26380 22148 26432 22200
rect 26380 21940 26432 21982
rect 26380 21930 26384 21940
rect 26384 21930 26430 21940
rect 26430 21930 26432 21940
rect 27854 24985 27897 24997
rect 27897 24985 27906 24997
rect 27854 24945 27906 24985
rect 27854 24779 27897 24780
rect 27897 24779 27906 24780
rect 27854 24728 27906 24779
rect 27854 24516 27906 24562
rect 27854 24510 27897 24516
rect 27897 24510 27906 24516
rect 27854 24310 27906 24344
rect 27854 24292 27897 24310
rect 27897 24292 27906 24310
rect 27854 24104 27906 24126
rect 27854 24074 27897 24104
rect 27897 24074 27906 24104
rect 27854 23898 27906 23909
rect 27854 23857 27897 23898
rect 27897 23857 27906 23898
rect 27557 22148 27609 22200
rect 27557 21940 27609 21982
rect 27557 21930 27561 21940
rect 27561 21930 27607 21940
rect 27607 21930 27609 21940
rect 28071 22148 28123 22200
rect 28071 21940 28123 21982
rect 28071 21930 28075 21940
rect 28075 21930 28121 21940
rect 28121 21930 28123 21940
rect 15381 21526 15385 21578
rect 15385 21526 15431 21578
rect 15431 21526 15433 21578
rect 25867 21513 25919 21565
rect 27558 21311 27610 21363
rect 6825 21110 6877 21162
rect 14204 21110 14256 21162
rect 24690 21110 24742 21162
rect 8002 20908 8054 20960
rect 15381 20908 15433 20960
rect 26381 20908 26433 20960
rect 8516 20706 8568 20758
rect 15895 20706 15947 20758
rect 28072 20706 28124 20758
rect 1814 20460 1817 20502
rect 1817 20460 1863 20502
rect 1863 20460 1866 20502
rect 1814 20450 1866 20460
rect 1814 20232 1866 20284
rect 1814 20015 1866 20067
rect 1814 19835 1866 19849
rect 1814 19797 1817 19835
rect 1817 19797 1863 19835
rect 1863 19797 1866 19835
rect 1814 19621 1817 19631
rect 1817 19621 1863 19631
rect 1863 19621 1866 19631
rect 1814 19579 1866 19621
rect 1814 19361 1866 19413
rect 1814 19164 1866 19196
rect 1814 19144 1817 19164
rect 1817 19144 1863 19164
rect 1863 19144 1866 19164
rect 1814 18950 1817 18978
rect 1817 18950 1863 18978
rect 1863 18950 1866 18978
rect 1814 18926 1866 18950
rect 2269 20338 2321 20364
rect 2269 20312 2312 20338
rect 2312 20312 2321 20338
rect 2552 20329 2604 20364
rect 2552 20312 2555 20329
rect 2555 20312 2601 20329
rect 2601 20312 2604 20329
rect 2835 20338 2887 20364
rect 2835 20312 2844 20338
rect 2844 20312 2887 20338
rect 2269 20125 2312 20146
rect 2312 20125 2321 20146
rect 2269 20094 2321 20125
rect 2552 20120 2555 20146
rect 2555 20120 2601 20146
rect 2601 20120 2604 20146
rect 2552 20094 2604 20120
rect 2835 20125 2844 20146
rect 2844 20125 2887 20146
rect 2835 20094 2887 20125
rect 2269 19877 2321 19929
rect 2552 19877 2604 19929
rect 2835 19877 2887 19929
rect 2269 19667 2321 19711
rect 2269 19659 2312 19667
rect 2312 19659 2321 19667
rect 2552 19676 2604 19711
rect 2552 19659 2555 19676
rect 2555 19659 2601 19676
rect 2601 19659 2604 19676
rect 2835 19667 2887 19711
rect 2835 19659 2844 19667
rect 2844 19659 2887 19667
rect 2269 19453 2312 19494
rect 2312 19453 2321 19494
rect 2269 19442 2321 19453
rect 2552 19467 2555 19494
rect 2555 19467 2601 19494
rect 2601 19467 2604 19494
rect 2552 19442 2604 19467
rect 2835 19453 2844 19494
rect 2844 19453 2887 19494
rect 2835 19442 2887 19453
rect 2269 19224 2321 19276
rect 2552 19224 2604 19276
rect 2835 19224 2887 19276
rect 2269 19006 2321 19058
rect 2552 19023 2604 19058
rect 2552 19006 2555 19023
rect 2555 19006 2601 19023
rect 2601 19006 2604 19023
rect 2835 19006 2887 19058
rect 3290 20460 3293 20502
rect 3293 20460 3339 20502
rect 3339 20460 3342 20502
rect 3290 20450 3342 20460
rect 3290 20232 3342 20284
rect 3290 20015 3342 20067
rect 3290 19835 3342 19849
rect 3290 19797 3293 19835
rect 3293 19797 3339 19835
rect 3339 19797 3342 19835
rect 3290 19621 3293 19631
rect 3293 19621 3339 19631
rect 3339 19621 3342 19631
rect 3290 19579 3342 19621
rect 3290 19361 3342 19413
rect 3290 19164 3342 19196
rect 3290 19144 3293 19164
rect 3293 19144 3339 19164
rect 3339 19144 3342 19164
rect 3290 18950 3293 18978
rect 3293 18950 3339 18978
rect 3339 18950 3342 18978
rect 3290 18926 3342 18950
rect 3606 20460 3609 20502
rect 3609 20460 3655 20502
rect 3655 20460 3658 20502
rect 3606 20450 3658 20460
rect 3606 20232 3658 20284
rect 3606 20015 3658 20067
rect 3606 19835 3658 19849
rect 3606 19797 3609 19835
rect 3609 19797 3655 19835
rect 3655 19797 3658 19835
rect 3606 19621 3609 19631
rect 3609 19621 3655 19631
rect 3655 19621 3658 19631
rect 3606 19579 3658 19621
rect 3606 19361 3658 19413
rect 3606 19164 3658 19196
rect 3606 19144 3609 19164
rect 3609 19144 3655 19164
rect 3655 19144 3658 19164
rect 3606 18950 3609 18978
rect 3609 18950 3655 18978
rect 3655 18950 3658 18978
rect 3606 18926 3658 18950
rect 4061 20338 4113 20364
rect 4061 20312 4104 20338
rect 4104 20312 4113 20338
rect 4344 20329 4396 20364
rect 4344 20312 4347 20329
rect 4347 20312 4393 20329
rect 4393 20312 4396 20329
rect 4627 20338 4679 20364
rect 4627 20312 4636 20338
rect 4636 20312 4679 20338
rect 4061 20125 4104 20146
rect 4104 20125 4113 20146
rect 4061 20094 4113 20125
rect 4344 20120 4347 20146
rect 4347 20120 4393 20146
rect 4393 20120 4396 20146
rect 4344 20094 4396 20120
rect 4627 20125 4636 20146
rect 4636 20125 4679 20146
rect 4627 20094 4679 20125
rect 4061 19877 4113 19929
rect 4344 19877 4396 19929
rect 4627 19877 4679 19929
rect 4061 19667 4113 19711
rect 4061 19659 4104 19667
rect 4104 19659 4113 19667
rect 4344 19676 4396 19711
rect 4344 19659 4347 19676
rect 4347 19659 4393 19676
rect 4393 19659 4396 19676
rect 4627 19667 4679 19711
rect 4627 19659 4636 19667
rect 4636 19659 4679 19667
rect 4061 19453 4104 19494
rect 4104 19453 4113 19494
rect 4061 19442 4113 19453
rect 4344 19467 4347 19494
rect 4347 19467 4393 19494
rect 4393 19467 4396 19494
rect 4344 19442 4396 19467
rect 4627 19453 4636 19494
rect 4636 19453 4679 19494
rect 4627 19442 4679 19453
rect 4061 19224 4113 19276
rect 4344 19224 4396 19276
rect 4627 19224 4679 19276
rect 4061 19006 4113 19058
rect 4344 19023 4396 19058
rect 4344 19006 4347 19023
rect 4347 19006 4393 19023
rect 4393 19006 4396 19023
rect 4627 19006 4679 19058
rect 2269 18828 2321 18840
rect 2269 18788 2312 18828
rect 2312 18788 2321 18828
rect 2552 18814 2555 18840
rect 2555 18814 2601 18840
rect 2601 18814 2604 18840
rect 2552 18788 2604 18814
rect 2835 18828 2887 18840
rect 2835 18788 2844 18828
rect 2844 18788 2887 18828
rect 2269 18612 2312 18623
rect 2312 18612 2321 18623
rect 2269 18571 2321 18612
rect 2552 18571 2604 18623
rect 2835 18612 2844 18623
rect 2844 18612 2887 18623
rect 2835 18571 2887 18612
rect 2269 18353 2321 18405
rect 2552 18371 2604 18405
rect 2552 18353 2555 18371
rect 2555 18353 2601 18371
rect 2601 18353 2604 18371
rect 2835 18353 2887 18405
rect 2269 18136 2321 18188
rect 2552 18161 2555 18188
rect 2555 18161 2601 18188
rect 2601 18161 2604 18188
rect 2552 18136 2604 18161
rect 2835 18136 2887 18188
rect 5082 20460 5085 20502
rect 5085 20460 5131 20502
rect 5131 20460 5134 20502
rect 5082 20450 5134 20460
rect 5082 20232 5134 20284
rect 5082 20015 5134 20067
rect 9193 20460 9196 20502
rect 9196 20460 9242 20502
rect 9242 20460 9245 20502
rect 9193 20450 9245 20460
rect 9193 20232 9245 20284
rect 9193 20015 9245 20067
rect 5082 19835 5134 19849
rect 5082 19797 5085 19835
rect 5085 19797 5131 19835
rect 5131 19797 5134 19835
rect 5082 19621 5085 19631
rect 5085 19621 5131 19631
rect 5131 19621 5134 19631
rect 5082 19579 5134 19621
rect 5874 19785 5926 19837
rect 5874 19567 5926 19619
rect 7565 19785 7617 19837
rect 7565 19567 7617 19619
rect 9193 19835 9245 19849
rect 9193 19797 9196 19835
rect 9196 19797 9242 19835
rect 9242 19797 9245 19835
rect 9193 19621 9196 19631
rect 9196 19621 9242 19631
rect 9242 19621 9245 19631
rect 9193 19579 9245 19621
rect 5082 19361 5134 19413
rect 5082 19164 5134 19196
rect 5082 19144 5085 19164
rect 5085 19144 5131 19164
rect 5131 19144 5134 19164
rect 5082 18950 5085 18978
rect 5085 18950 5131 18978
rect 5131 18950 5134 18978
rect 5082 18926 5134 18950
rect 9193 19361 9245 19413
rect 9193 19164 9245 19196
rect 9193 19144 9196 19164
rect 9196 19144 9242 19164
rect 9242 19144 9245 19164
rect 9193 18950 9196 18978
rect 9196 18950 9242 18978
rect 9242 18950 9245 18978
rect 9193 18926 9245 18950
rect 9648 20338 9700 20364
rect 9648 20312 9691 20338
rect 9691 20312 9700 20338
rect 9931 20329 9983 20364
rect 9931 20312 9934 20329
rect 9934 20312 9980 20329
rect 9980 20312 9983 20329
rect 10214 20338 10266 20364
rect 10214 20312 10223 20338
rect 10223 20312 10266 20338
rect 9648 20125 9691 20146
rect 9691 20125 9700 20146
rect 9648 20094 9700 20125
rect 9931 20120 9934 20146
rect 9934 20120 9980 20146
rect 9980 20120 9983 20146
rect 9931 20094 9983 20120
rect 10214 20125 10223 20146
rect 10223 20125 10266 20146
rect 10214 20094 10266 20125
rect 9648 19877 9700 19929
rect 9931 19877 9983 19929
rect 10214 19877 10266 19929
rect 9648 19667 9700 19711
rect 9648 19659 9691 19667
rect 9691 19659 9700 19667
rect 9931 19676 9983 19711
rect 9931 19659 9934 19676
rect 9934 19659 9980 19676
rect 9980 19659 9983 19676
rect 10214 19667 10266 19711
rect 10214 19659 10223 19667
rect 10223 19659 10266 19667
rect 9648 19453 9691 19494
rect 9691 19453 9700 19494
rect 9648 19442 9700 19453
rect 9931 19467 9934 19494
rect 9934 19467 9980 19494
rect 9980 19467 9983 19494
rect 9931 19442 9983 19467
rect 10214 19453 10223 19494
rect 10223 19453 10266 19494
rect 10214 19442 10266 19453
rect 9648 19224 9700 19276
rect 9931 19224 9983 19276
rect 10214 19224 10266 19276
rect 9648 19006 9700 19058
rect 9931 19023 9983 19058
rect 9931 19006 9934 19023
rect 9934 19006 9980 19023
rect 9980 19006 9983 19023
rect 10214 19006 10266 19058
rect 4061 18828 4113 18840
rect 4061 18788 4104 18828
rect 4104 18788 4113 18828
rect 4344 18814 4347 18840
rect 4347 18814 4393 18840
rect 4393 18814 4396 18840
rect 4344 18788 4396 18814
rect 4627 18828 4679 18840
rect 4627 18788 4636 18828
rect 4636 18788 4679 18828
rect 4061 18612 4104 18623
rect 4104 18612 4113 18623
rect 4061 18571 4113 18612
rect 4344 18571 4396 18623
rect 4627 18612 4636 18623
rect 4636 18612 4679 18623
rect 4627 18571 4679 18612
rect 4061 18353 4113 18405
rect 4344 18371 4396 18405
rect 4344 18353 4347 18371
rect 4347 18353 4393 18371
rect 4393 18353 4396 18371
rect 4627 18353 4679 18405
rect 4061 18136 4113 18188
rect 4344 18161 4347 18188
rect 4347 18161 4393 18188
rect 4393 18161 4396 18188
rect 4344 18136 4396 18161
rect 4627 18136 4679 18188
rect 2269 17918 2321 17970
rect 2552 17918 2604 17970
rect 2835 17918 2887 17970
rect 10669 20460 10672 20502
rect 10672 20460 10718 20502
rect 10718 20460 10721 20502
rect 10669 20450 10721 20460
rect 10669 20232 10721 20284
rect 10669 20015 10721 20067
rect 10669 19835 10721 19849
rect 10669 19797 10672 19835
rect 10672 19797 10718 19835
rect 10718 19797 10721 19835
rect 10669 19621 10672 19631
rect 10672 19621 10718 19631
rect 10718 19621 10721 19631
rect 10669 19579 10721 19621
rect 10669 19361 10721 19413
rect 10669 19164 10721 19196
rect 10669 19144 10672 19164
rect 10672 19144 10718 19164
rect 10718 19144 10721 19164
rect 10669 18950 10672 18978
rect 10672 18950 10718 18978
rect 10718 18950 10721 18978
rect 10669 18926 10721 18950
rect 10985 20460 10988 20502
rect 10988 20460 11034 20502
rect 11034 20460 11037 20502
rect 10985 20450 11037 20460
rect 10985 20232 11037 20284
rect 10985 20015 11037 20067
rect 10985 19835 11037 19849
rect 10985 19797 10988 19835
rect 10988 19797 11034 19835
rect 11034 19797 11037 19835
rect 10985 19621 10988 19631
rect 10988 19621 11034 19631
rect 11034 19621 11037 19631
rect 10985 19579 11037 19621
rect 10985 19361 11037 19413
rect 10985 19164 11037 19196
rect 10985 19144 10988 19164
rect 10988 19144 11034 19164
rect 11034 19144 11037 19164
rect 10985 18950 10988 18978
rect 10988 18950 11034 18978
rect 11034 18950 11037 18978
rect 10985 18926 11037 18950
rect 11440 20338 11492 20364
rect 11440 20312 11483 20338
rect 11483 20312 11492 20338
rect 11723 20329 11775 20364
rect 11723 20312 11726 20329
rect 11726 20312 11772 20329
rect 11772 20312 11775 20329
rect 12006 20338 12058 20364
rect 12006 20312 12015 20338
rect 12015 20312 12058 20338
rect 11440 20125 11483 20146
rect 11483 20125 11492 20146
rect 11440 20094 11492 20125
rect 11723 20120 11726 20146
rect 11726 20120 11772 20146
rect 11772 20120 11775 20146
rect 11723 20094 11775 20120
rect 12006 20125 12015 20146
rect 12015 20125 12058 20146
rect 12006 20094 12058 20125
rect 11440 19877 11492 19929
rect 11723 19877 11775 19929
rect 12006 19877 12058 19929
rect 11440 19667 11492 19711
rect 11440 19659 11483 19667
rect 11483 19659 11492 19667
rect 11723 19676 11775 19711
rect 11723 19659 11726 19676
rect 11726 19659 11772 19676
rect 11772 19659 11775 19676
rect 12006 19667 12058 19711
rect 12006 19659 12015 19667
rect 12015 19659 12058 19667
rect 11440 19453 11483 19494
rect 11483 19453 11492 19494
rect 11440 19442 11492 19453
rect 11723 19467 11726 19494
rect 11726 19467 11772 19494
rect 11772 19467 11775 19494
rect 11723 19442 11775 19467
rect 12006 19453 12015 19494
rect 12015 19453 12058 19494
rect 12006 19442 12058 19453
rect 11440 19224 11492 19276
rect 11723 19224 11775 19276
rect 12006 19224 12058 19276
rect 11440 19006 11492 19058
rect 11723 19023 11775 19058
rect 11723 19006 11726 19023
rect 11726 19006 11772 19023
rect 11772 19006 11775 19023
rect 12006 19006 12058 19058
rect 9648 18828 9700 18840
rect 9648 18788 9691 18828
rect 9691 18788 9700 18828
rect 9931 18814 9934 18840
rect 9934 18814 9980 18840
rect 9980 18814 9983 18840
rect 9931 18788 9983 18814
rect 10214 18828 10266 18840
rect 10214 18788 10223 18828
rect 10223 18788 10266 18828
rect 9648 18612 9691 18623
rect 9691 18612 9700 18623
rect 9648 18571 9700 18612
rect 9931 18571 9983 18623
rect 10214 18612 10223 18623
rect 10223 18612 10266 18623
rect 10214 18571 10266 18612
rect 9648 18353 9700 18405
rect 9931 18371 9983 18405
rect 9931 18353 9934 18371
rect 9934 18353 9980 18371
rect 9980 18353 9983 18371
rect 10214 18353 10266 18405
rect 9648 18136 9700 18188
rect 9931 18161 9934 18188
rect 9934 18161 9980 18188
rect 9980 18161 9983 18188
rect 9931 18136 9983 18161
rect 10214 18136 10266 18188
rect 4061 17918 4113 17970
rect 4344 17918 4396 17970
rect 4627 17918 4679 17970
rect 12461 20460 12464 20502
rect 12464 20460 12510 20502
rect 12510 20460 12513 20502
rect 12461 20450 12513 20460
rect 12461 20232 12513 20284
rect 12461 20015 12513 20067
rect 16701 20446 16704 20489
rect 16704 20446 16750 20489
rect 16750 20446 16753 20489
rect 16701 20437 16753 20446
rect 18045 20446 18048 20489
rect 18048 20446 18094 20489
rect 18094 20446 18097 20489
rect 18045 20437 18097 20446
rect 16701 20219 16753 20271
rect 16701 20002 16753 20054
rect 12461 19835 12513 19849
rect 12461 19797 12464 19835
rect 12464 19797 12510 19835
rect 12510 19797 12513 19835
rect 12461 19621 12464 19631
rect 12464 19621 12510 19631
rect 12510 19621 12513 19631
rect 12461 19579 12513 19621
rect 13253 19785 13305 19837
rect 13253 19567 13305 19619
rect 14944 19785 14996 19837
rect 14944 19567 14996 19619
rect 16701 19821 16753 19836
rect 16701 19784 16704 19821
rect 16704 19784 16750 19821
rect 16750 19784 16753 19821
rect 16701 19608 16704 19618
rect 16704 19608 16750 19618
rect 16750 19608 16753 19618
rect 16701 19566 16753 19608
rect 12461 19361 12513 19413
rect 12461 19164 12513 19196
rect 12461 19144 12464 19164
rect 12464 19144 12510 19164
rect 12510 19144 12513 19164
rect 12461 18950 12464 18978
rect 12464 18950 12510 18978
rect 12510 18950 12513 18978
rect 12461 18926 12513 18950
rect 16701 19348 16753 19400
rect 16701 19150 16753 19183
rect 16701 19131 16704 19150
rect 16704 19131 16750 19150
rect 16750 19131 16753 19150
rect 16701 18936 16704 18965
rect 16704 18936 16750 18965
rect 16750 18936 16753 18965
rect 16701 18913 16753 18936
rect 11440 18828 11492 18840
rect 11440 18788 11483 18828
rect 11483 18788 11492 18828
rect 11723 18814 11726 18840
rect 11726 18814 11772 18840
rect 11772 18814 11775 18840
rect 11723 18788 11775 18814
rect 12006 18828 12058 18840
rect 12006 18788 12015 18828
rect 12015 18788 12058 18828
rect 11440 18612 11483 18623
rect 11483 18612 11492 18623
rect 11440 18571 11492 18612
rect 11723 18571 11775 18623
rect 12006 18612 12015 18623
rect 12015 18612 12058 18623
rect 12006 18571 12058 18612
rect 11440 18353 11492 18405
rect 11723 18371 11775 18405
rect 11723 18353 11726 18371
rect 11726 18353 11772 18371
rect 11772 18353 11775 18371
rect 12006 18353 12058 18405
rect 11440 18136 11492 18188
rect 11723 18161 11726 18188
rect 11726 18161 11772 18188
rect 11772 18161 11775 18188
rect 11723 18136 11775 18161
rect 12006 18136 12058 18188
rect 9648 17918 9700 17970
rect 9931 17918 9983 17970
rect 10214 17918 10266 17970
rect 17373 20333 17425 20385
rect 17373 20157 17425 20167
rect 17373 20115 17376 20157
rect 17376 20115 17422 20157
rect 17422 20115 17425 20157
rect 17373 19943 17376 19950
rect 17376 19943 17422 19950
rect 17422 19943 17425 19950
rect 17373 19898 17425 19943
rect 17373 19680 17425 19732
rect 17373 19486 17425 19514
rect 17373 19462 17376 19486
rect 17376 19462 17422 19486
rect 17422 19462 17425 19486
rect 17373 19272 17376 19297
rect 17376 19272 17422 19297
rect 17422 19272 17425 19297
rect 17373 19245 17425 19272
rect 17373 19027 17425 19079
rect 18045 20219 18097 20271
rect 18045 20002 18097 20054
rect 18045 19821 18097 19836
rect 18045 19784 18048 19821
rect 18048 19784 18094 19821
rect 18094 19784 18097 19821
rect 18045 19608 18048 19618
rect 18048 19608 18094 19618
rect 18094 19608 18097 19618
rect 18045 19566 18097 19608
rect 18045 19348 18097 19400
rect 18045 19150 18097 19183
rect 18045 19131 18048 19150
rect 18048 19131 18094 19150
rect 18094 19131 18097 19150
rect 18045 18936 18048 18965
rect 18048 18936 18094 18965
rect 18094 18936 18097 18965
rect 18045 18913 18097 18936
rect 18335 20446 18338 20489
rect 18338 20446 18384 20489
rect 18384 20446 18387 20489
rect 18335 20437 18387 20446
rect 19679 20446 19682 20489
rect 19682 20446 19728 20489
rect 19728 20446 19731 20489
rect 19679 20437 19731 20446
rect 18335 20219 18387 20271
rect 18335 20002 18387 20054
rect 18335 19821 18387 19836
rect 18335 19784 18338 19821
rect 18338 19784 18384 19821
rect 18384 19784 18387 19821
rect 18335 19608 18338 19618
rect 18338 19608 18384 19618
rect 18384 19608 18387 19618
rect 18335 19566 18387 19608
rect 18335 19348 18387 19400
rect 18335 19150 18387 19183
rect 18335 19131 18338 19150
rect 18338 19131 18384 19150
rect 18384 19131 18387 19150
rect 18335 18936 18338 18965
rect 18338 18936 18384 18965
rect 18384 18936 18387 18965
rect 18335 18913 18387 18936
rect 19007 20333 19059 20385
rect 19007 20157 19059 20167
rect 19007 20115 19010 20157
rect 19010 20115 19056 20157
rect 19056 20115 19059 20157
rect 19007 19943 19010 19950
rect 19010 19943 19056 19950
rect 19056 19943 19059 19950
rect 19007 19898 19059 19943
rect 19007 19680 19059 19732
rect 19007 19486 19059 19514
rect 19007 19462 19010 19486
rect 19010 19462 19056 19486
rect 19056 19462 19059 19486
rect 19007 19272 19010 19297
rect 19010 19272 19056 19297
rect 19056 19272 19059 19297
rect 19007 19245 19059 19272
rect 19007 19027 19059 19079
rect 17373 18815 17425 18861
rect 17373 18809 17376 18815
rect 17376 18809 17422 18815
rect 17422 18809 17425 18815
rect 17373 18599 17376 18644
rect 17376 18599 17422 18644
rect 17422 18599 17425 18644
rect 17373 18592 17425 18599
rect 17373 18374 17425 18426
rect 17373 18156 17425 18208
rect 11440 17918 11492 17970
rect 11723 17918 11775 17970
rect 12006 17918 12058 17970
rect 19679 20219 19731 20271
rect 19679 20002 19731 20054
rect 19679 19821 19731 19836
rect 19679 19784 19682 19821
rect 19682 19784 19728 19821
rect 19728 19784 19731 19821
rect 19679 19608 19682 19618
rect 19682 19608 19728 19618
rect 19728 19608 19731 19618
rect 19679 19566 19731 19608
rect 19679 19348 19731 19400
rect 19679 19150 19731 19183
rect 19679 19131 19682 19150
rect 19682 19131 19728 19150
rect 19728 19131 19731 19150
rect 19679 18936 19682 18965
rect 19682 18936 19728 18965
rect 19728 18936 19731 18965
rect 19679 18913 19731 18936
rect 19968 20446 19971 20489
rect 19971 20446 20017 20489
rect 20017 20446 20020 20489
rect 19968 20437 20020 20446
rect 21312 20446 21315 20489
rect 21315 20446 21361 20489
rect 21361 20446 21364 20489
rect 21312 20437 21364 20446
rect 19968 20219 20020 20271
rect 19968 20002 20020 20054
rect 19968 19821 20020 19836
rect 19968 19784 19971 19821
rect 19971 19784 20017 19821
rect 20017 19784 20020 19821
rect 19968 19608 19971 19618
rect 19971 19608 20017 19618
rect 20017 19608 20020 19618
rect 19968 19566 20020 19608
rect 19968 19348 20020 19400
rect 19968 19150 20020 19183
rect 19968 19131 19971 19150
rect 19971 19131 20017 19150
rect 20017 19131 20020 19150
rect 19968 18936 19971 18965
rect 19971 18936 20017 18965
rect 20017 18936 20020 18965
rect 19968 18913 20020 18936
rect 20640 20333 20692 20385
rect 20640 20157 20692 20167
rect 20640 20115 20643 20157
rect 20643 20115 20689 20157
rect 20689 20115 20692 20157
rect 20640 19943 20643 19950
rect 20643 19943 20689 19950
rect 20689 19943 20692 19950
rect 20640 19898 20692 19943
rect 20640 19680 20692 19732
rect 20640 19486 20692 19514
rect 20640 19462 20643 19486
rect 20643 19462 20689 19486
rect 20689 19462 20692 19486
rect 20640 19272 20643 19297
rect 20643 19272 20689 19297
rect 20689 19272 20692 19297
rect 20640 19245 20692 19272
rect 20640 19027 20692 19079
rect 19007 18815 19059 18861
rect 19007 18809 19010 18815
rect 19010 18809 19056 18815
rect 19056 18809 19059 18815
rect 19007 18599 19010 18644
rect 19010 18599 19056 18644
rect 19056 18599 19059 18644
rect 19007 18592 19059 18599
rect 19007 18374 19059 18426
rect 19007 18156 19059 18208
rect 17373 17939 17425 17991
rect 21312 20219 21364 20271
rect 21312 20002 21364 20054
rect 21312 19821 21364 19836
rect 21312 19784 21315 19821
rect 21315 19784 21361 19821
rect 21361 19784 21364 19821
rect 21312 19608 21315 19618
rect 21315 19608 21361 19618
rect 21361 19608 21364 19618
rect 21312 19566 21364 19608
rect 21312 19348 21364 19400
rect 21312 19150 21364 19183
rect 21312 19131 21315 19150
rect 21315 19131 21361 19150
rect 21361 19131 21364 19150
rect 21312 18936 21315 18965
rect 21315 18936 21361 18965
rect 21361 18936 21364 18965
rect 21312 18913 21364 18936
rect 21602 20446 21605 20489
rect 21605 20446 21651 20489
rect 21651 20446 21654 20489
rect 21602 20437 21654 20446
rect 22946 20446 22949 20489
rect 22949 20446 22995 20489
rect 22995 20446 22998 20489
rect 22946 20437 22998 20446
rect 21602 20219 21654 20271
rect 21602 20002 21654 20054
rect 21602 19821 21654 19836
rect 21602 19784 21605 19821
rect 21605 19784 21651 19821
rect 21651 19784 21654 19821
rect 21602 19608 21605 19618
rect 21605 19608 21651 19618
rect 21651 19608 21654 19618
rect 21602 19566 21654 19608
rect 21602 19348 21654 19400
rect 21602 19150 21654 19183
rect 21602 19131 21605 19150
rect 21605 19131 21651 19150
rect 21651 19131 21654 19150
rect 21602 18936 21605 18965
rect 21605 18936 21651 18965
rect 21651 18936 21654 18965
rect 21602 18913 21654 18936
rect 22274 20333 22326 20385
rect 22274 20157 22326 20167
rect 22274 20115 22277 20157
rect 22277 20115 22323 20157
rect 22323 20115 22326 20157
rect 22274 19943 22277 19950
rect 22277 19943 22323 19950
rect 22323 19943 22326 19950
rect 22274 19898 22326 19943
rect 22274 19680 22326 19732
rect 22274 19486 22326 19514
rect 22274 19462 22277 19486
rect 22277 19462 22323 19486
rect 22323 19462 22326 19486
rect 22274 19272 22277 19297
rect 22277 19272 22323 19297
rect 22323 19272 22326 19297
rect 22274 19245 22326 19272
rect 22274 19027 22326 19079
rect 20640 18815 20692 18861
rect 20640 18809 20643 18815
rect 20643 18809 20689 18815
rect 20689 18809 20692 18815
rect 20640 18599 20643 18644
rect 20643 18599 20689 18644
rect 20689 18599 20692 18644
rect 20640 18592 20692 18599
rect 20640 18374 20692 18426
rect 20640 18156 20692 18208
rect 19007 17939 19059 17991
rect 22946 20219 22998 20271
rect 22946 20002 22998 20054
rect 22946 19821 22998 19836
rect 22946 19784 22949 19821
rect 22949 19784 22995 19821
rect 22995 19784 22998 19821
rect 22946 19608 22949 19618
rect 22949 19608 22995 19618
rect 22995 19608 22998 19618
rect 22946 19566 22998 19608
rect 23739 19785 23791 19837
rect 23739 19567 23791 19619
rect 25429 19785 25481 19837
rect 25429 19567 25481 19619
rect 27120 19785 27172 19837
rect 27120 19567 27172 19619
rect 22946 19348 22998 19400
rect 22946 19150 22998 19183
rect 22946 19131 22949 19150
rect 22949 19131 22995 19150
rect 22995 19131 22998 19150
rect 22946 18936 22949 18965
rect 22949 18936 22995 18965
rect 22995 18936 22998 18965
rect 22946 18913 22998 18936
rect 22274 18815 22326 18861
rect 22274 18809 22277 18815
rect 22277 18809 22323 18815
rect 22323 18809 22326 18815
rect 22274 18599 22277 18644
rect 22277 18599 22323 18644
rect 22323 18599 22326 18644
rect 22274 18592 22326 18599
rect 22274 18374 22326 18426
rect 22274 18156 22326 18208
rect 20640 17939 20692 17991
rect 22274 17939 22326 17991
rect 17373 17721 17425 17773
rect 19007 17721 19059 17773
rect 20640 17721 20692 17773
rect 22274 17721 22326 17773
rect 1992 16887 2044 16902
rect 2664 16887 2716 16902
rect 3112 16887 3164 16902
rect 3784 16887 3836 16902
rect 4232 16887 4284 16902
rect 1992 16850 2012 16887
rect 2012 16850 2044 16887
rect 2664 16850 2691 16887
rect 2691 16850 2716 16887
rect 3112 16850 3119 16887
rect 3119 16850 3164 16887
rect 3784 16850 3798 16887
rect 3798 16850 3836 16887
rect 4232 16850 4272 16887
rect 4272 16850 4284 16887
rect 4904 16850 4956 16902
rect 5352 16887 5404 16902
rect 5352 16850 5379 16887
rect 5379 16850 5404 16887
rect 6024 16850 6076 16902
rect 6472 16887 6524 16902
rect 6472 16850 6486 16887
rect 6486 16850 6524 16887
rect 7144 16850 7196 16902
rect 7592 16850 7644 16902
rect 8264 16850 8316 16902
rect 8712 16850 8764 16902
rect 9384 16850 9436 16902
rect 9832 16850 9884 16902
rect 10504 16887 10556 16902
rect 10504 16850 10551 16887
rect 10551 16850 10556 16887
rect 10952 16850 11004 16902
rect 11624 16887 11676 16902
rect 11624 16850 11658 16887
rect 11658 16850 11676 16887
rect 12072 16850 12124 16902
rect 12744 16887 12796 16902
rect 13192 16887 13244 16902
rect 13864 16887 13916 16902
rect 14312 16887 14364 16902
rect 14984 16887 15036 16902
rect 15432 16887 15484 16902
rect 16104 16887 16156 16902
rect 16552 16887 16604 16902
rect 17224 16887 17276 16902
rect 17672 16887 17724 16902
rect 12744 16850 12764 16887
rect 12764 16850 12796 16887
rect 13192 16850 13239 16887
rect 13239 16850 13244 16887
rect 13864 16850 13871 16887
rect 13871 16850 13916 16887
rect 14312 16850 14345 16887
rect 14345 16850 14364 16887
rect 14984 16850 15024 16887
rect 15024 16850 15036 16887
rect 15432 16850 15452 16887
rect 15452 16850 15484 16887
rect 16104 16850 16131 16887
rect 16131 16850 16156 16887
rect 16552 16850 16559 16887
rect 16559 16850 16604 16887
rect 17224 16850 17238 16887
rect 17238 16850 17276 16887
rect 17672 16850 17712 16887
rect 17712 16850 17724 16887
rect 18344 16850 18396 16902
rect 18792 16887 18844 16902
rect 18792 16850 18819 16887
rect 18819 16850 18844 16887
rect 19464 16850 19516 16902
rect 19912 16887 19964 16902
rect 19912 16850 19925 16887
rect 19925 16850 19964 16887
rect 1992 16726 2044 16778
rect 2664 16726 2716 16778
rect 3112 16726 3164 16778
rect 3784 16726 3836 16778
rect 4232 16726 4284 16778
rect 4904 16726 4956 16778
rect 5352 16726 5404 16778
rect 6024 16726 6076 16778
rect 6472 16726 6524 16778
rect 7144 16726 7196 16778
rect 7592 16726 7644 16778
rect 8264 16726 8316 16778
rect 8712 16726 8764 16778
rect 9384 16726 9436 16778
rect 9832 16726 9884 16778
rect 10504 16726 10556 16778
rect 10952 16726 11004 16778
rect 11624 16726 11676 16778
rect 12072 16726 12124 16778
rect 12744 16726 12796 16778
rect 13192 16726 13244 16778
rect 13864 16726 13916 16778
rect 14312 16726 14364 16778
rect 14984 16726 15036 16778
rect 15432 16726 15484 16778
rect 16104 16726 16156 16778
rect 16552 16726 16604 16778
rect 17224 16726 17276 16778
rect 17672 16726 17724 16778
rect 18344 16726 18396 16778
rect 18792 16726 18844 16778
rect 19464 16726 19516 16778
rect 19912 16726 19964 16778
rect 1992 16602 2044 16654
rect 2664 16602 2716 16654
rect 1992 16478 1995 16530
rect 1995 16478 2041 16530
rect 2041 16478 2044 16530
rect 1992 16354 1995 16406
rect 1995 16354 2041 16406
rect 2041 16354 2044 16406
rect 1992 16230 1995 16282
rect 1995 16230 2041 16282
rect 2041 16230 2044 16282
rect 1992 16106 1995 16158
rect 1995 16106 2041 16158
rect 2041 16106 2044 16158
rect 1992 15982 1995 16034
rect 1995 15982 2041 16034
rect 2041 15982 2044 16034
rect 1992 15858 1995 15910
rect 1995 15858 2041 15910
rect 2041 15858 2044 15910
rect 1992 15734 1995 15786
rect 1995 15734 2041 15786
rect 2041 15734 2044 15786
rect 1992 15610 1995 15662
rect 1995 15610 2041 15662
rect 2041 15610 2044 15662
rect 1992 15486 1995 15538
rect 1995 15486 2041 15538
rect 2041 15486 2044 15538
rect 3112 16602 3164 16654
rect 2664 16478 2667 16530
rect 2667 16478 2713 16530
rect 2713 16478 2716 16530
rect 2664 16354 2667 16406
rect 2667 16354 2713 16406
rect 2713 16354 2716 16406
rect 2664 16230 2667 16282
rect 2667 16230 2713 16282
rect 2713 16230 2716 16282
rect 2664 16106 2667 16158
rect 2667 16106 2713 16158
rect 2713 16106 2716 16158
rect 2664 15982 2667 16034
rect 2667 15982 2713 16034
rect 2713 15982 2716 16034
rect 2664 15858 2667 15910
rect 2667 15858 2713 15910
rect 2713 15858 2716 15910
rect 2664 15734 2667 15786
rect 2667 15734 2713 15786
rect 2713 15734 2716 15786
rect 2664 15610 2667 15662
rect 2667 15610 2713 15662
rect 2713 15610 2716 15662
rect 2664 15486 2667 15538
rect 2667 15486 2713 15538
rect 2713 15486 2716 15538
rect 2440 14944 2443 14996
rect 2443 14944 2489 14996
rect 2489 14944 2492 14996
rect 2440 14820 2443 14872
rect 2443 14820 2489 14872
rect 2489 14820 2492 14872
rect 2440 14696 2443 14748
rect 2443 14696 2489 14748
rect 2489 14696 2492 14748
rect 2440 14572 2443 14624
rect 2443 14572 2489 14624
rect 2489 14572 2492 14624
rect 2440 14448 2443 14500
rect 2443 14448 2489 14500
rect 2489 14448 2492 14500
rect 2440 14324 2443 14376
rect 2443 14324 2489 14376
rect 2489 14324 2492 14376
rect 2440 14200 2443 14252
rect 2443 14200 2489 14252
rect 2489 14200 2492 14252
rect 2440 14076 2443 14128
rect 2443 14076 2489 14128
rect 2489 14076 2492 14128
rect 2440 13952 2443 14004
rect 2443 13952 2489 14004
rect 2489 13952 2492 14004
rect 2440 13828 2443 13880
rect 2443 13828 2489 13880
rect 2489 13828 2492 13880
rect 2440 13704 2443 13756
rect 2443 13704 2489 13756
rect 2489 13704 2492 13756
rect 2440 13580 2443 13632
rect 2443 13580 2489 13632
rect 2489 13580 2492 13632
rect 2440 13456 2443 13508
rect 2443 13456 2489 13508
rect 2489 13456 2492 13508
rect 2440 13332 2443 13384
rect 2443 13332 2489 13384
rect 2489 13332 2492 13384
rect 2440 13208 2443 13260
rect 2443 13208 2489 13260
rect 2489 13208 2492 13260
rect 2440 13084 2443 13136
rect 2443 13084 2489 13136
rect 2489 13084 2492 13136
rect 2440 12960 2443 13012
rect 2443 12960 2489 13012
rect 2489 12960 2492 13012
rect 2440 12836 2443 12888
rect 2443 12836 2489 12888
rect 2489 12836 2492 12888
rect 2008 11859 2060 11911
rect 3784 16602 3836 16654
rect 3112 16478 3115 16530
rect 3115 16478 3161 16530
rect 3161 16478 3164 16530
rect 3112 16354 3115 16406
rect 3115 16354 3161 16406
rect 3161 16354 3164 16406
rect 3112 16230 3115 16282
rect 3115 16230 3161 16282
rect 3161 16230 3164 16282
rect 3112 16106 3115 16158
rect 3115 16106 3161 16158
rect 3161 16106 3164 16158
rect 3112 15982 3115 16034
rect 3115 15982 3161 16034
rect 3161 15982 3164 16034
rect 3112 15858 3115 15910
rect 3115 15858 3161 15910
rect 3161 15858 3164 15910
rect 3112 15734 3115 15786
rect 3115 15734 3161 15786
rect 3161 15734 3164 15786
rect 3112 15610 3115 15662
rect 3115 15610 3161 15662
rect 3161 15610 3164 15662
rect 3112 15486 3115 15538
rect 3115 15486 3161 15538
rect 3161 15486 3164 15538
rect 2888 14944 2891 14996
rect 2891 14944 2937 14996
rect 2937 14944 2940 14996
rect 2888 14820 2891 14872
rect 2891 14820 2937 14872
rect 2937 14820 2940 14872
rect 2888 14696 2891 14748
rect 2891 14696 2937 14748
rect 2937 14696 2940 14748
rect 2888 14572 2891 14624
rect 2891 14572 2937 14624
rect 2937 14572 2940 14624
rect 2888 14448 2891 14500
rect 2891 14448 2937 14500
rect 2937 14448 2940 14500
rect 2888 14324 2891 14376
rect 2891 14324 2937 14376
rect 2937 14324 2940 14376
rect 2888 14200 2891 14252
rect 2891 14200 2937 14252
rect 2937 14200 2940 14252
rect 2888 14076 2891 14128
rect 2891 14076 2937 14128
rect 2937 14076 2940 14128
rect 2888 13952 2891 14004
rect 2891 13952 2937 14004
rect 2937 13952 2940 14004
rect 2888 13828 2891 13880
rect 2891 13828 2937 13880
rect 2937 13828 2940 13880
rect 2888 13704 2891 13756
rect 2891 13704 2937 13756
rect 2937 13704 2940 13756
rect 2888 13580 2891 13632
rect 2891 13580 2937 13632
rect 2937 13580 2940 13632
rect 2888 13456 2891 13508
rect 2891 13456 2937 13508
rect 2937 13456 2940 13508
rect 2888 13332 2891 13384
rect 2891 13332 2937 13384
rect 2937 13332 2940 13384
rect 2888 13208 2891 13260
rect 2891 13208 2937 13260
rect 2937 13208 2940 13260
rect 2888 13084 2891 13136
rect 2891 13084 2937 13136
rect 2937 13084 2940 13136
rect 2888 12960 2891 13012
rect 2891 12960 2937 13012
rect 2937 12960 2940 13012
rect 2888 12836 2891 12888
rect 2891 12836 2937 12888
rect 2937 12836 2940 12888
rect 4232 16602 4284 16654
rect 3784 16478 3787 16530
rect 3787 16478 3833 16530
rect 3833 16478 3836 16530
rect 3784 16354 3787 16406
rect 3787 16354 3833 16406
rect 3833 16354 3836 16406
rect 3784 16230 3787 16282
rect 3787 16230 3833 16282
rect 3833 16230 3836 16282
rect 3784 16106 3787 16158
rect 3787 16106 3833 16158
rect 3833 16106 3836 16158
rect 3784 15982 3787 16034
rect 3787 15982 3833 16034
rect 3833 15982 3836 16034
rect 3784 15858 3787 15910
rect 3787 15858 3833 15910
rect 3833 15858 3836 15910
rect 3784 15734 3787 15786
rect 3787 15734 3833 15786
rect 3833 15734 3836 15786
rect 3784 15610 3787 15662
rect 3787 15610 3833 15662
rect 3833 15610 3836 15662
rect 3784 15486 3787 15538
rect 3787 15486 3833 15538
rect 3833 15486 3836 15538
rect 3560 14944 3563 14996
rect 3563 14944 3609 14996
rect 3609 14944 3612 14996
rect 3560 14820 3563 14872
rect 3563 14820 3609 14872
rect 3609 14820 3612 14872
rect 3560 14696 3563 14748
rect 3563 14696 3609 14748
rect 3609 14696 3612 14748
rect 3560 14572 3563 14624
rect 3563 14572 3609 14624
rect 3609 14572 3612 14624
rect 3560 14448 3563 14500
rect 3563 14448 3609 14500
rect 3609 14448 3612 14500
rect 3560 14324 3563 14376
rect 3563 14324 3609 14376
rect 3609 14324 3612 14376
rect 3560 14200 3563 14252
rect 3563 14200 3609 14252
rect 3609 14200 3612 14252
rect 3560 14076 3563 14128
rect 3563 14076 3609 14128
rect 3609 14076 3612 14128
rect 3560 13952 3563 14004
rect 3563 13952 3609 14004
rect 3609 13952 3612 14004
rect 3560 13828 3563 13880
rect 3563 13828 3609 13880
rect 3609 13828 3612 13880
rect 3560 13704 3563 13756
rect 3563 13704 3609 13756
rect 3609 13704 3612 13756
rect 3560 13580 3563 13632
rect 3563 13580 3609 13632
rect 3609 13580 3612 13632
rect 3560 13456 3563 13508
rect 3563 13456 3609 13508
rect 3609 13456 3612 13508
rect 3560 13332 3563 13384
rect 3563 13332 3609 13384
rect 3609 13332 3612 13384
rect 3560 13208 3563 13260
rect 3563 13208 3609 13260
rect 3609 13208 3612 13260
rect 3560 13084 3563 13136
rect 3563 13084 3609 13136
rect 3609 13084 3612 13136
rect 3560 12960 3563 13012
rect 3563 12960 3609 13012
rect 3609 12960 3612 13012
rect 3560 12836 3563 12888
rect 3563 12836 3609 12888
rect 3609 12836 3612 12888
rect 444 1065 496 1117
rect 444 847 496 899
rect 1270 1065 1322 1117
rect 1270 847 1322 899
rect 1511 1065 1563 1117
rect 1511 847 1563 899
rect 3128 11859 3180 11911
rect 4904 16602 4956 16654
rect 4232 16478 4235 16530
rect 4235 16478 4281 16530
rect 4281 16478 4284 16530
rect 4232 16354 4235 16406
rect 4235 16354 4281 16406
rect 4281 16354 4284 16406
rect 4232 16230 4235 16282
rect 4235 16230 4281 16282
rect 4281 16230 4284 16282
rect 4232 16106 4235 16158
rect 4235 16106 4281 16158
rect 4281 16106 4284 16158
rect 4232 15982 4235 16034
rect 4235 15982 4281 16034
rect 4281 15982 4284 16034
rect 4232 15858 4235 15910
rect 4235 15858 4281 15910
rect 4281 15858 4284 15910
rect 4232 15734 4235 15786
rect 4235 15734 4281 15786
rect 4281 15734 4284 15786
rect 4232 15610 4235 15662
rect 4235 15610 4281 15662
rect 4281 15610 4284 15662
rect 4232 15486 4235 15538
rect 4235 15486 4281 15538
rect 4281 15486 4284 15538
rect 4008 14944 4011 14996
rect 4011 14944 4057 14996
rect 4057 14944 4060 14996
rect 4008 14820 4011 14872
rect 4011 14820 4057 14872
rect 4057 14820 4060 14872
rect 4008 14696 4011 14748
rect 4011 14696 4057 14748
rect 4057 14696 4060 14748
rect 4008 14572 4011 14624
rect 4011 14572 4057 14624
rect 4057 14572 4060 14624
rect 4008 14448 4011 14500
rect 4011 14448 4057 14500
rect 4057 14448 4060 14500
rect 4008 14324 4011 14376
rect 4011 14324 4057 14376
rect 4057 14324 4060 14376
rect 4008 14200 4011 14252
rect 4011 14200 4057 14252
rect 4057 14200 4060 14252
rect 4008 14076 4011 14128
rect 4011 14076 4057 14128
rect 4057 14076 4060 14128
rect 4008 13952 4011 14004
rect 4011 13952 4057 14004
rect 4057 13952 4060 14004
rect 4008 13828 4011 13880
rect 4011 13828 4057 13880
rect 4057 13828 4060 13880
rect 4008 13704 4011 13756
rect 4011 13704 4057 13756
rect 4057 13704 4060 13756
rect 4008 13580 4011 13632
rect 4011 13580 4057 13632
rect 4057 13580 4060 13632
rect 4008 13456 4011 13508
rect 4011 13456 4057 13508
rect 4057 13456 4060 13508
rect 4008 13332 4011 13384
rect 4011 13332 4057 13384
rect 4057 13332 4060 13384
rect 4008 13208 4011 13260
rect 4011 13208 4057 13260
rect 4057 13208 4060 13260
rect 4008 13084 4011 13136
rect 4011 13084 4057 13136
rect 4057 13084 4060 13136
rect 4008 12960 4011 13012
rect 4011 12960 4057 13012
rect 4057 12960 4060 13012
rect 4008 12836 4011 12888
rect 4011 12836 4057 12888
rect 4057 12836 4060 12888
rect 5352 16602 5404 16654
rect 4904 16478 4907 16530
rect 4907 16478 4953 16530
rect 4953 16478 4956 16530
rect 4904 16354 4907 16406
rect 4907 16354 4953 16406
rect 4953 16354 4956 16406
rect 4904 16230 4907 16282
rect 4907 16230 4953 16282
rect 4953 16230 4956 16282
rect 4904 16106 4907 16158
rect 4907 16106 4953 16158
rect 4953 16106 4956 16158
rect 4904 15982 4907 16034
rect 4907 15982 4953 16034
rect 4953 15982 4956 16034
rect 4904 15858 4907 15910
rect 4907 15858 4953 15910
rect 4953 15858 4956 15910
rect 4904 15734 4907 15786
rect 4907 15734 4953 15786
rect 4953 15734 4956 15786
rect 4904 15610 4907 15662
rect 4907 15610 4953 15662
rect 4953 15610 4956 15662
rect 4904 15486 4907 15538
rect 4907 15486 4953 15538
rect 4953 15486 4956 15538
rect 4680 14944 4683 14996
rect 4683 14944 4729 14996
rect 4729 14944 4732 14996
rect 4680 14820 4683 14872
rect 4683 14820 4729 14872
rect 4729 14820 4732 14872
rect 4680 14696 4683 14748
rect 4683 14696 4729 14748
rect 4729 14696 4732 14748
rect 4680 14572 4683 14624
rect 4683 14572 4729 14624
rect 4729 14572 4732 14624
rect 4680 14448 4683 14500
rect 4683 14448 4729 14500
rect 4729 14448 4732 14500
rect 4680 14324 4683 14376
rect 4683 14324 4729 14376
rect 4729 14324 4732 14376
rect 4680 14200 4683 14252
rect 4683 14200 4729 14252
rect 4729 14200 4732 14252
rect 4680 14076 4683 14128
rect 4683 14076 4729 14128
rect 4729 14076 4732 14128
rect 4680 13952 4683 14004
rect 4683 13952 4729 14004
rect 4729 13952 4732 14004
rect 4680 13828 4683 13880
rect 4683 13828 4729 13880
rect 4729 13828 4732 13880
rect 4680 13704 4683 13756
rect 4683 13704 4729 13756
rect 4729 13704 4732 13756
rect 4680 13580 4683 13632
rect 4683 13580 4729 13632
rect 4729 13580 4732 13632
rect 4680 13456 4683 13508
rect 4683 13456 4729 13508
rect 4729 13456 4732 13508
rect 4680 13332 4683 13384
rect 4683 13332 4729 13384
rect 4729 13332 4732 13384
rect 4680 13208 4683 13260
rect 4683 13208 4729 13260
rect 4729 13208 4732 13260
rect 4680 13084 4683 13136
rect 4683 13084 4729 13136
rect 4729 13084 4732 13136
rect 4680 12960 4683 13012
rect 4683 12960 4729 13012
rect 4729 12960 4732 13012
rect 4680 12836 4683 12888
rect 4683 12836 4729 12888
rect 4729 12836 4732 12888
rect 2440 11757 2492 11758
rect 2440 11706 2443 11757
rect 2443 11706 2489 11757
rect 2489 11706 2492 11757
rect 2440 11582 2443 11634
rect 2443 11582 2489 11634
rect 2489 11582 2492 11634
rect 2440 11458 2443 11510
rect 2443 11458 2489 11510
rect 2489 11458 2492 11510
rect 2888 11757 2940 11758
rect 2888 11706 2891 11757
rect 2891 11706 2937 11757
rect 2937 11706 2940 11757
rect 2888 11582 2891 11634
rect 2891 11582 2937 11634
rect 2937 11582 2940 11634
rect 2888 11458 2891 11510
rect 2891 11458 2937 11510
rect 2937 11458 2940 11510
rect 4248 11859 4300 11911
rect 6024 16602 6076 16654
rect 5352 16478 5355 16530
rect 5355 16478 5401 16530
rect 5401 16478 5404 16530
rect 5352 16354 5355 16406
rect 5355 16354 5401 16406
rect 5401 16354 5404 16406
rect 5352 16230 5355 16282
rect 5355 16230 5401 16282
rect 5401 16230 5404 16282
rect 5352 16106 5355 16158
rect 5355 16106 5401 16158
rect 5401 16106 5404 16158
rect 5352 15982 5355 16034
rect 5355 15982 5401 16034
rect 5401 15982 5404 16034
rect 5352 15858 5355 15910
rect 5355 15858 5401 15910
rect 5401 15858 5404 15910
rect 5352 15734 5355 15786
rect 5355 15734 5401 15786
rect 5401 15734 5404 15786
rect 5352 15610 5355 15662
rect 5355 15610 5401 15662
rect 5401 15610 5404 15662
rect 5352 15486 5355 15538
rect 5355 15486 5401 15538
rect 5401 15486 5404 15538
rect 5128 14944 5131 14996
rect 5131 14944 5177 14996
rect 5177 14944 5180 14996
rect 5128 14820 5131 14872
rect 5131 14820 5177 14872
rect 5177 14820 5180 14872
rect 5128 14696 5131 14748
rect 5131 14696 5177 14748
rect 5177 14696 5180 14748
rect 5128 14572 5131 14624
rect 5131 14572 5177 14624
rect 5177 14572 5180 14624
rect 5128 14448 5131 14500
rect 5131 14448 5177 14500
rect 5177 14448 5180 14500
rect 5128 14324 5131 14376
rect 5131 14324 5177 14376
rect 5177 14324 5180 14376
rect 5128 14200 5131 14252
rect 5131 14200 5177 14252
rect 5177 14200 5180 14252
rect 5128 14076 5131 14128
rect 5131 14076 5177 14128
rect 5177 14076 5180 14128
rect 5128 13952 5131 14004
rect 5131 13952 5177 14004
rect 5177 13952 5180 14004
rect 5128 13828 5131 13880
rect 5131 13828 5177 13880
rect 5177 13828 5180 13880
rect 5128 13704 5131 13756
rect 5131 13704 5177 13756
rect 5177 13704 5180 13756
rect 5128 13580 5131 13632
rect 5131 13580 5177 13632
rect 5177 13580 5180 13632
rect 5128 13456 5131 13508
rect 5131 13456 5177 13508
rect 5177 13456 5180 13508
rect 5128 13332 5131 13384
rect 5131 13332 5177 13384
rect 5177 13332 5180 13384
rect 5128 13208 5131 13260
rect 5131 13208 5177 13260
rect 5177 13208 5180 13260
rect 5128 13084 5131 13136
rect 5131 13084 5177 13136
rect 5177 13084 5180 13136
rect 5128 12960 5131 13012
rect 5131 12960 5177 13012
rect 5177 12960 5180 13012
rect 5128 12836 5131 12888
rect 5131 12836 5177 12888
rect 5177 12836 5180 12888
rect 6472 16602 6524 16654
rect 6024 16478 6027 16530
rect 6027 16478 6073 16530
rect 6073 16478 6076 16530
rect 6024 16354 6027 16406
rect 6027 16354 6073 16406
rect 6073 16354 6076 16406
rect 6024 16230 6027 16282
rect 6027 16230 6073 16282
rect 6073 16230 6076 16282
rect 6024 16106 6027 16158
rect 6027 16106 6073 16158
rect 6073 16106 6076 16158
rect 6024 15982 6027 16034
rect 6027 15982 6073 16034
rect 6073 15982 6076 16034
rect 6024 15858 6027 15910
rect 6027 15858 6073 15910
rect 6073 15858 6076 15910
rect 6024 15734 6027 15786
rect 6027 15734 6073 15786
rect 6073 15734 6076 15786
rect 6024 15610 6027 15662
rect 6027 15610 6073 15662
rect 6073 15610 6076 15662
rect 6024 15486 6027 15538
rect 6027 15486 6073 15538
rect 6073 15486 6076 15538
rect 5800 14944 5803 14996
rect 5803 14944 5849 14996
rect 5849 14944 5852 14996
rect 5800 14820 5803 14872
rect 5803 14820 5849 14872
rect 5849 14820 5852 14872
rect 5800 14696 5803 14748
rect 5803 14696 5849 14748
rect 5849 14696 5852 14748
rect 5800 14572 5803 14624
rect 5803 14572 5849 14624
rect 5849 14572 5852 14624
rect 5800 14448 5803 14500
rect 5803 14448 5849 14500
rect 5849 14448 5852 14500
rect 5800 14324 5803 14376
rect 5803 14324 5849 14376
rect 5849 14324 5852 14376
rect 5800 14200 5803 14252
rect 5803 14200 5849 14252
rect 5849 14200 5852 14252
rect 5800 14076 5803 14128
rect 5803 14076 5849 14128
rect 5849 14076 5852 14128
rect 5800 13952 5803 14004
rect 5803 13952 5849 14004
rect 5849 13952 5852 14004
rect 5800 13828 5803 13880
rect 5803 13828 5849 13880
rect 5849 13828 5852 13880
rect 5800 13704 5803 13756
rect 5803 13704 5849 13756
rect 5849 13704 5852 13756
rect 5800 13580 5803 13632
rect 5803 13580 5849 13632
rect 5849 13580 5852 13632
rect 5800 13456 5803 13508
rect 5803 13456 5849 13508
rect 5849 13456 5852 13508
rect 5800 13332 5803 13384
rect 5803 13332 5849 13384
rect 5849 13332 5852 13384
rect 5800 13208 5803 13260
rect 5803 13208 5849 13260
rect 5849 13208 5852 13260
rect 5800 13084 5803 13136
rect 5803 13084 5849 13136
rect 5849 13084 5852 13136
rect 5800 12960 5803 13012
rect 5803 12960 5849 13012
rect 5849 12960 5852 13012
rect 5800 12836 5803 12888
rect 5803 12836 5849 12888
rect 5849 12836 5852 12888
rect 3560 11757 3612 11758
rect 3560 11706 3563 11757
rect 3563 11706 3609 11757
rect 3609 11706 3612 11757
rect 3560 11582 3563 11634
rect 3563 11582 3609 11634
rect 3609 11582 3612 11634
rect 3560 11458 3563 11510
rect 3563 11458 3609 11510
rect 3609 11458 3612 11510
rect 4008 11757 4060 11758
rect 4008 11706 4011 11757
rect 4011 11706 4057 11757
rect 4057 11706 4060 11757
rect 4008 11582 4011 11634
rect 4011 11582 4057 11634
rect 4057 11582 4060 11634
rect 4008 11458 4011 11510
rect 4011 11458 4057 11510
rect 4057 11458 4060 11510
rect 5368 11859 5420 11911
rect 7144 16602 7196 16654
rect 6472 16478 6475 16530
rect 6475 16478 6521 16530
rect 6521 16478 6524 16530
rect 6472 16354 6475 16406
rect 6475 16354 6521 16406
rect 6521 16354 6524 16406
rect 6472 16230 6475 16282
rect 6475 16230 6521 16282
rect 6521 16230 6524 16282
rect 6472 16106 6475 16158
rect 6475 16106 6521 16158
rect 6521 16106 6524 16158
rect 6472 15982 6475 16034
rect 6475 15982 6521 16034
rect 6521 15982 6524 16034
rect 6472 15858 6475 15910
rect 6475 15858 6521 15910
rect 6521 15858 6524 15910
rect 6472 15734 6475 15786
rect 6475 15734 6521 15786
rect 6521 15734 6524 15786
rect 6472 15610 6475 15662
rect 6475 15610 6521 15662
rect 6521 15610 6524 15662
rect 6472 15486 6475 15538
rect 6475 15486 6521 15538
rect 6521 15486 6524 15538
rect 6248 14944 6251 14996
rect 6251 14944 6297 14996
rect 6297 14944 6300 14996
rect 6248 14820 6251 14872
rect 6251 14820 6297 14872
rect 6297 14820 6300 14872
rect 6248 14696 6251 14748
rect 6251 14696 6297 14748
rect 6297 14696 6300 14748
rect 6248 14572 6251 14624
rect 6251 14572 6297 14624
rect 6297 14572 6300 14624
rect 6248 14448 6251 14500
rect 6251 14448 6297 14500
rect 6297 14448 6300 14500
rect 6248 14324 6251 14376
rect 6251 14324 6297 14376
rect 6297 14324 6300 14376
rect 6248 14200 6251 14252
rect 6251 14200 6297 14252
rect 6297 14200 6300 14252
rect 6248 14076 6251 14128
rect 6251 14076 6297 14128
rect 6297 14076 6300 14128
rect 6248 13952 6251 14004
rect 6251 13952 6297 14004
rect 6297 13952 6300 14004
rect 6248 13828 6251 13880
rect 6251 13828 6297 13880
rect 6297 13828 6300 13880
rect 6248 13704 6251 13756
rect 6251 13704 6297 13756
rect 6297 13704 6300 13756
rect 6248 13580 6251 13632
rect 6251 13580 6297 13632
rect 6297 13580 6300 13632
rect 6248 13456 6251 13508
rect 6251 13456 6297 13508
rect 6297 13456 6300 13508
rect 6248 13332 6251 13384
rect 6251 13332 6297 13384
rect 6297 13332 6300 13384
rect 6248 13208 6251 13260
rect 6251 13208 6297 13260
rect 6297 13208 6300 13260
rect 6248 13084 6251 13136
rect 6251 13084 6297 13136
rect 6297 13084 6300 13136
rect 6248 12960 6251 13012
rect 6251 12960 6297 13012
rect 6297 12960 6300 13012
rect 6248 12836 6251 12888
rect 6251 12836 6297 12888
rect 6297 12836 6300 12888
rect 7592 16602 7644 16654
rect 7144 16478 7147 16530
rect 7147 16478 7193 16530
rect 7193 16478 7196 16530
rect 7144 16354 7147 16406
rect 7147 16354 7193 16406
rect 7193 16354 7196 16406
rect 7144 16230 7147 16282
rect 7147 16230 7193 16282
rect 7193 16230 7196 16282
rect 7144 16106 7147 16158
rect 7147 16106 7193 16158
rect 7193 16106 7196 16158
rect 7144 15982 7147 16034
rect 7147 15982 7193 16034
rect 7193 15982 7196 16034
rect 7144 15858 7147 15910
rect 7147 15858 7193 15910
rect 7193 15858 7196 15910
rect 7144 15734 7147 15786
rect 7147 15734 7193 15786
rect 7193 15734 7196 15786
rect 7144 15610 7147 15662
rect 7147 15610 7193 15662
rect 7193 15610 7196 15662
rect 7144 15486 7147 15538
rect 7147 15486 7193 15538
rect 7193 15486 7196 15538
rect 6920 14944 6923 14996
rect 6923 14944 6969 14996
rect 6969 14944 6972 14996
rect 6920 14820 6923 14872
rect 6923 14820 6969 14872
rect 6969 14820 6972 14872
rect 6920 14696 6923 14748
rect 6923 14696 6969 14748
rect 6969 14696 6972 14748
rect 6920 14572 6923 14624
rect 6923 14572 6969 14624
rect 6969 14572 6972 14624
rect 6920 14448 6923 14500
rect 6923 14448 6969 14500
rect 6969 14448 6972 14500
rect 6920 14324 6923 14376
rect 6923 14324 6969 14376
rect 6969 14324 6972 14376
rect 6920 14200 6923 14252
rect 6923 14200 6969 14252
rect 6969 14200 6972 14252
rect 6920 14076 6923 14128
rect 6923 14076 6969 14128
rect 6969 14076 6972 14128
rect 6920 13952 6923 14004
rect 6923 13952 6969 14004
rect 6969 13952 6972 14004
rect 6920 13828 6923 13880
rect 6923 13828 6969 13880
rect 6969 13828 6972 13880
rect 6920 13704 6923 13756
rect 6923 13704 6969 13756
rect 6969 13704 6972 13756
rect 6920 13580 6923 13632
rect 6923 13580 6969 13632
rect 6969 13580 6972 13632
rect 6920 13456 6923 13508
rect 6923 13456 6969 13508
rect 6969 13456 6972 13508
rect 6920 13332 6923 13384
rect 6923 13332 6969 13384
rect 6969 13332 6972 13384
rect 6920 13208 6923 13260
rect 6923 13208 6969 13260
rect 6969 13208 6972 13260
rect 6920 13084 6923 13136
rect 6923 13084 6969 13136
rect 6969 13084 6972 13136
rect 6920 12960 6923 13012
rect 6923 12960 6969 13012
rect 6969 12960 6972 13012
rect 6920 12836 6923 12888
rect 6923 12836 6969 12888
rect 6969 12836 6972 12888
rect 4680 11757 4732 11758
rect 4680 11706 4683 11757
rect 4683 11706 4729 11757
rect 4729 11706 4732 11757
rect 4680 11582 4683 11634
rect 4683 11582 4729 11634
rect 4729 11582 4732 11634
rect 4680 11458 4683 11510
rect 4683 11458 4729 11510
rect 4729 11458 4732 11510
rect 5128 11757 5180 11758
rect 5128 11706 5131 11757
rect 5131 11706 5177 11757
rect 5177 11706 5180 11757
rect 5128 11582 5131 11634
rect 5131 11582 5177 11634
rect 5177 11582 5180 11634
rect 5128 11458 5131 11510
rect 5131 11458 5177 11510
rect 5177 11458 5180 11510
rect 6488 11859 6540 11911
rect 8264 16602 8316 16654
rect 7592 16478 7595 16530
rect 7595 16478 7641 16530
rect 7641 16478 7644 16530
rect 7592 16354 7595 16406
rect 7595 16354 7641 16406
rect 7641 16354 7644 16406
rect 7592 16230 7595 16282
rect 7595 16230 7641 16282
rect 7641 16230 7644 16282
rect 7592 16106 7595 16158
rect 7595 16106 7641 16158
rect 7641 16106 7644 16158
rect 7592 15982 7595 16034
rect 7595 15982 7641 16034
rect 7641 15982 7644 16034
rect 7592 15858 7595 15910
rect 7595 15858 7641 15910
rect 7641 15858 7644 15910
rect 7592 15734 7595 15786
rect 7595 15734 7641 15786
rect 7641 15734 7644 15786
rect 7592 15610 7595 15662
rect 7595 15610 7641 15662
rect 7641 15610 7644 15662
rect 7592 15486 7595 15538
rect 7595 15486 7641 15538
rect 7641 15486 7644 15538
rect 7368 14944 7371 14996
rect 7371 14944 7417 14996
rect 7417 14944 7420 14996
rect 7368 14820 7371 14872
rect 7371 14820 7417 14872
rect 7417 14820 7420 14872
rect 7368 14696 7371 14748
rect 7371 14696 7417 14748
rect 7417 14696 7420 14748
rect 7368 14572 7371 14624
rect 7371 14572 7417 14624
rect 7417 14572 7420 14624
rect 7368 14448 7371 14500
rect 7371 14448 7417 14500
rect 7417 14448 7420 14500
rect 7368 14324 7371 14376
rect 7371 14324 7417 14376
rect 7417 14324 7420 14376
rect 7368 14200 7371 14252
rect 7371 14200 7417 14252
rect 7417 14200 7420 14252
rect 7368 14076 7371 14128
rect 7371 14076 7417 14128
rect 7417 14076 7420 14128
rect 7368 13952 7371 14004
rect 7371 13952 7417 14004
rect 7417 13952 7420 14004
rect 7368 13828 7371 13880
rect 7371 13828 7417 13880
rect 7417 13828 7420 13880
rect 7368 13704 7371 13756
rect 7371 13704 7417 13756
rect 7417 13704 7420 13756
rect 7368 13580 7371 13632
rect 7371 13580 7417 13632
rect 7417 13580 7420 13632
rect 7368 13456 7371 13508
rect 7371 13456 7417 13508
rect 7417 13456 7420 13508
rect 7368 13332 7371 13384
rect 7371 13332 7417 13384
rect 7417 13332 7420 13384
rect 7368 13208 7371 13260
rect 7371 13208 7417 13260
rect 7417 13208 7420 13260
rect 7368 13084 7371 13136
rect 7371 13084 7417 13136
rect 7417 13084 7420 13136
rect 7368 12960 7371 13012
rect 7371 12960 7417 13012
rect 7417 12960 7420 13012
rect 7368 12836 7371 12888
rect 7371 12836 7417 12888
rect 7417 12836 7420 12888
rect 8712 16602 8764 16654
rect 8264 16478 8267 16530
rect 8267 16478 8313 16530
rect 8313 16478 8316 16530
rect 8264 16354 8267 16406
rect 8267 16354 8313 16406
rect 8313 16354 8316 16406
rect 8264 16230 8267 16282
rect 8267 16230 8313 16282
rect 8313 16230 8316 16282
rect 8264 16106 8267 16158
rect 8267 16106 8313 16158
rect 8313 16106 8316 16158
rect 8264 15982 8267 16034
rect 8267 15982 8313 16034
rect 8313 15982 8316 16034
rect 8264 15858 8267 15910
rect 8267 15858 8313 15910
rect 8313 15858 8316 15910
rect 8264 15734 8267 15786
rect 8267 15734 8313 15786
rect 8313 15734 8316 15786
rect 8264 15610 8267 15662
rect 8267 15610 8313 15662
rect 8313 15610 8316 15662
rect 8264 15486 8267 15538
rect 8267 15486 8313 15538
rect 8313 15486 8316 15538
rect 8040 14944 8043 14996
rect 8043 14944 8089 14996
rect 8089 14944 8092 14996
rect 8040 14820 8043 14872
rect 8043 14820 8089 14872
rect 8089 14820 8092 14872
rect 8040 14696 8043 14748
rect 8043 14696 8089 14748
rect 8089 14696 8092 14748
rect 8040 14572 8043 14624
rect 8043 14572 8089 14624
rect 8089 14572 8092 14624
rect 8040 14448 8043 14500
rect 8043 14448 8089 14500
rect 8089 14448 8092 14500
rect 8040 14324 8043 14376
rect 8043 14324 8089 14376
rect 8089 14324 8092 14376
rect 8040 14200 8043 14252
rect 8043 14200 8089 14252
rect 8089 14200 8092 14252
rect 8040 14076 8043 14128
rect 8043 14076 8089 14128
rect 8089 14076 8092 14128
rect 8040 13952 8043 14004
rect 8043 13952 8089 14004
rect 8089 13952 8092 14004
rect 8040 13828 8043 13880
rect 8043 13828 8089 13880
rect 8089 13828 8092 13880
rect 8040 13704 8043 13756
rect 8043 13704 8089 13756
rect 8089 13704 8092 13756
rect 8040 13580 8043 13632
rect 8043 13580 8089 13632
rect 8089 13580 8092 13632
rect 8040 13456 8043 13508
rect 8043 13456 8089 13508
rect 8089 13456 8092 13508
rect 8040 13332 8043 13384
rect 8043 13332 8089 13384
rect 8089 13332 8092 13384
rect 8040 13208 8043 13260
rect 8043 13208 8089 13260
rect 8089 13208 8092 13260
rect 8040 13084 8043 13136
rect 8043 13084 8089 13136
rect 8089 13084 8092 13136
rect 8040 12960 8043 13012
rect 8043 12960 8089 13012
rect 8089 12960 8092 13012
rect 8040 12836 8043 12888
rect 8043 12836 8089 12888
rect 8089 12836 8092 12888
rect 5800 11757 5852 11758
rect 5800 11706 5803 11757
rect 5803 11706 5849 11757
rect 5849 11706 5852 11757
rect 5800 11582 5803 11634
rect 5803 11582 5849 11634
rect 5849 11582 5852 11634
rect 5800 11458 5803 11510
rect 5803 11458 5849 11510
rect 5849 11458 5852 11510
rect 6248 11757 6300 11758
rect 6248 11706 6251 11757
rect 6251 11706 6297 11757
rect 6297 11706 6300 11757
rect 6248 11582 6251 11634
rect 6251 11582 6297 11634
rect 6297 11582 6300 11634
rect 6248 11458 6251 11510
rect 6251 11458 6297 11510
rect 6297 11458 6300 11510
rect 7608 11859 7660 11911
rect 9384 16602 9436 16654
rect 8712 16478 8715 16530
rect 8715 16478 8761 16530
rect 8761 16478 8764 16530
rect 8712 16354 8715 16406
rect 8715 16354 8761 16406
rect 8761 16354 8764 16406
rect 8712 16230 8715 16282
rect 8715 16230 8761 16282
rect 8761 16230 8764 16282
rect 8712 16106 8715 16158
rect 8715 16106 8761 16158
rect 8761 16106 8764 16158
rect 8712 15982 8715 16034
rect 8715 15982 8761 16034
rect 8761 15982 8764 16034
rect 8712 15858 8715 15910
rect 8715 15858 8761 15910
rect 8761 15858 8764 15910
rect 8712 15734 8715 15786
rect 8715 15734 8761 15786
rect 8761 15734 8764 15786
rect 8712 15610 8715 15662
rect 8715 15610 8761 15662
rect 8761 15610 8764 15662
rect 8712 15486 8715 15538
rect 8715 15486 8761 15538
rect 8761 15486 8764 15538
rect 8488 14944 8491 14996
rect 8491 14944 8537 14996
rect 8537 14944 8540 14996
rect 8488 14820 8491 14872
rect 8491 14820 8537 14872
rect 8537 14820 8540 14872
rect 8488 14696 8491 14748
rect 8491 14696 8537 14748
rect 8537 14696 8540 14748
rect 8488 14572 8491 14624
rect 8491 14572 8537 14624
rect 8537 14572 8540 14624
rect 8488 14448 8491 14500
rect 8491 14448 8537 14500
rect 8537 14448 8540 14500
rect 8488 14324 8491 14376
rect 8491 14324 8537 14376
rect 8537 14324 8540 14376
rect 8488 14200 8491 14252
rect 8491 14200 8537 14252
rect 8537 14200 8540 14252
rect 8488 14076 8491 14128
rect 8491 14076 8537 14128
rect 8537 14076 8540 14128
rect 8488 13952 8491 14004
rect 8491 13952 8537 14004
rect 8537 13952 8540 14004
rect 8488 13828 8491 13880
rect 8491 13828 8537 13880
rect 8537 13828 8540 13880
rect 8488 13704 8491 13756
rect 8491 13704 8537 13756
rect 8537 13704 8540 13756
rect 8488 13580 8491 13632
rect 8491 13580 8537 13632
rect 8537 13580 8540 13632
rect 8488 13456 8491 13508
rect 8491 13456 8537 13508
rect 8537 13456 8540 13508
rect 8488 13332 8491 13384
rect 8491 13332 8537 13384
rect 8537 13332 8540 13384
rect 8488 13208 8491 13260
rect 8491 13208 8537 13260
rect 8537 13208 8540 13260
rect 8488 13084 8491 13136
rect 8491 13084 8537 13136
rect 8537 13084 8540 13136
rect 8488 12960 8491 13012
rect 8491 12960 8537 13012
rect 8537 12960 8540 13012
rect 8488 12836 8491 12888
rect 8491 12836 8537 12888
rect 8537 12836 8540 12888
rect 9832 16602 9884 16654
rect 9384 16478 9387 16530
rect 9387 16478 9433 16530
rect 9433 16478 9436 16530
rect 9384 16354 9387 16406
rect 9387 16354 9433 16406
rect 9433 16354 9436 16406
rect 9384 16230 9387 16282
rect 9387 16230 9433 16282
rect 9433 16230 9436 16282
rect 9384 16106 9387 16158
rect 9387 16106 9433 16158
rect 9433 16106 9436 16158
rect 9384 15982 9387 16034
rect 9387 15982 9433 16034
rect 9433 15982 9436 16034
rect 9384 15858 9387 15910
rect 9387 15858 9433 15910
rect 9433 15858 9436 15910
rect 9384 15734 9387 15786
rect 9387 15734 9433 15786
rect 9433 15734 9436 15786
rect 9384 15610 9387 15662
rect 9387 15610 9433 15662
rect 9433 15610 9436 15662
rect 9384 15486 9387 15538
rect 9387 15486 9433 15538
rect 9433 15486 9436 15538
rect 9160 14944 9163 14996
rect 9163 14944 9209 14996
rect 9209 14944 9212 14996
rect 9160 14820 9163 14872
rect 9163 14820 9209 14872
rect 9209 14820 9212 14872
rect 9160 14696 9163 14748
rect 9163 14696 9209 14748
rect 9209 14696 9212 14748
rect 9160 14572 9163 14624
rect 9163 14572 9209 14624
rect 9209 14572 9212 14624
rect 9160 14448 9163 14500
rect 9163 14448 9209 14500
rect 9209 14448 9212 14500
rect 9160 14324 9163 14376
rect 9163 14324 9209 14376
rect 9209 14324 9212 14376
rect 9160 14200 9163 14252
rect 9163 14200 9209 14252
rect 9209 14200 9212 14252
rect 9160 14076 9163 14128
rect 9163 14076 9209 14128
rect 9209 14076 9212 14128
rect 9160 13952 9163 14004
rect 9163 13952 9209 14004
rect 9209 13952 9212 14004
rect 9160 13828 9163 13880
rect 9163 13828 9209 13880
rect 9209 13828 9212 13880
rect 9160 13704 9163 13756
rect 9163 13704 9209 13756
rect 9209 13704 9212 13756
rect 9160 13580 9163 13632
rect 9163 13580 9209 13632
rect 9209 13580 9212 13632
rect 9160 13456 9163 13508
rect 9163 13456 9209 13508
rect 9209 13456 9212 13508
rect 9160 13332 9163 13384
rect 9163 13332 9209 13384
rect 9209 13332 9212 13384
rect 9160 13208 9163 13260
rect 9163 13208 9209 13260
rect 9209 13208 9212 13260
rect 9160 13084 9163 13136
rect 9163 13084 9209 13136
rect 9209 13084 9212 13136
rect 9160 12960 9163 13012
rect 9163 12960 9209 13012
rect 9209 12960 9212 13012
rect 9160 12836 9163 12888
rect 9163 12836 9209 12888
rect 9209 12836 9212 12888
rect 6920 11757 6972 11758
rect 6920 11706 6923 11757
rect 6923 11706 6969 11757
rect 6969 11706 6972 11757
rect 6920 11582 6923 11634
rect 6923 11582 6969 11634
rect 6969 11582 6972 11634
rect 6920 11458 6923 11510
rect 6923 11458 6969 11510
rect 6969 11458 6972 11510
rect 7368 11757 7420 11758
rect 7368 11706 7371 11757
rect 7371 11706 7417 11757
rect 7417 11706 7420 11757
rect 7368 11582 7371 11634
rect 7371 11582 7417 11634
rect 7417 11582 7420 11634
rect 7368 11458 7371 11510
rect 7371 11458 7417 11510
rect 7417 11458 7420 11510
rect 8728 11859 8780 11911
rect 10504 16602 10556 16654
rect 9832 16478 9835 16530
rect 9835 16478 9881 16530
rect 9881 16478 9884 16530
rect 9832 16354 9835 16406
rect 9835 16354 9881 16406
rect 9881 16354 9884 16406
rect 9832 16230 9835 16282
rect 9835 16230 9881 16282
rect 9881 16230 9884 16282
rect 9832 16106 9835 16158
rect 9835 16106 9881 16158
rect 9881 16106 9884 16158
rect 9832 15982 9835 16034
rect 9835 15982 9881 16034
rect 9881 15982 9884 16034
rect 9832 15858 9835 15910
rect 9835 15858 9881 15910
rect 9881 15858 9884 15910
rect 9832 15734 9835 15786
rect 9835 15734 9881 15786
rect 9881 15734 9884 15786
rect 9832 15610 9835 15662
rect 9835 15610 9881 15662
rect 9881 15610 9884 15662
rect 9832 15486 9835 15538
rect 9835 15486 9881 15538
rect 9881 15486 9884 15538
rect 9608 14944 9611 14996
rect 9611 14944 9657 14996
rect 9657 14944 9660 14996
rect 9608 14820 9611 14872
rect 9611 14820 9657 14872
rect 9657 14820 9660 14872
rect 9608 14696 9611 14748
rect 9611 14696 9657 14748
rect 9657 14696 9660 14748
rect 9608 14572 9611 14624
rect 9611 14572 9657 14624
rect 9657 14572 9660 14624
rect 9608 14448 9611 14500
rect 9611 14448 9657 14500
rect 9657 14448 9660 14500
rect 9608 14324 9611 14376
rect 9611 14324 9657 14376
rect 9657 14324 9660 14376
rect 9608 14200 9611 14252
rect 9611 14200 9657 14252
rect 9657 14200 9660 14252
rect 9608 14076 9611 14128
rect 9611 14076 9657 14128
rect 9657 14076 9660 14128
rect 9608 13952 9611 14004
rect 9611 13952 9657 14004
rect 9657 13952 9660 14004
rect 9608 13828 9611 13880
rect 9611 13828 9657 13880
rect 9657 13828 9660 13880
rect 9608 13704 9611 13756
rect 9611 13704 9657 13756
rect 9657 13704 9660 13756
rect 9608 13580 9611 13632
rect 9611 13580 9657 13632
rect 9657 13580 9660 13632
rect 9608 13456 9611 13508
rect 9611 13456 9657 13508
rect 9657 13456 9660 13508
rect 9608 13332 9611 13384
rect 9611 13332 9657 13384
rect 9657 13332 9660 13384
rect 9608 13208 9611 13260
rect 9611 13208 9657 13260
rect 9657 13208 9660 13260
rect 9608 13084 9611 13136
rect 9611 13084 9657 13136
rect 9657 13084 9660 13136
rect 9608 12960 9611 13012
rect 9611 12960 9657 13012
rect 9657 12960 9660 13012
rect 9608 12836 9611 12888
rect 9611 12836 9657 12888
rect 9657 12836 9660 12888
rect 10952 16602 11004 16654
rect 10504 16478 10507 16530
rect 10507 16478 10553 16530
rect 10553 16478 10556 16530
rect 10504 16354 10507 16406
rect 10507 16354 10553 16406
rect 10553 16354 10556 16406
rect 10504 16230 10507 16282
rect 10507 16230 10553 16282
rect 10553 16230 10556 16282
rect 10504 16106 10507 16158
rect 10507 16106 10553 16158
rect 10553 16106 10556 16158
rect 10504 15982 10507 16034
rect 10507 15982 10553 16034
rect 10553 15982 10556 16034
rect 10504 15858 10507 15910
rect 10507 15858 10553 15910
rect 10553 15858 10556 15910
rect 10504 15734 10507 15786
rect 10507 15734 10553 15786
rect 10553 15734 10556 15786
rect 10504 15610 10507 15662
rect 10507 15610 10553 15662
rect 10553 15610 10556 15662
rect 10504 15486 10507 15538
rect 10507 15486 10553 15538
rect 10553 15486 10556 15538
rect 10280 14944 10283 14996
rect 10283 14944 10329 14996
rect 10329 14944 10332 14996
rect 10280 14820 10283 14872
rect 10283 14820 10329 14872
rect 10329 14820 10332 14872
rect 10280 14696 10283 14748
rect 10283 14696 10329 14748
rect 10329 14696 10332 14748
rect 10280 14572 10283 14624
rect 10283 14572 10329 14624
rect 10329 14572 10332 14624
rect 10280 14448 10283 14500
rect 10283 14448 10329 14500
rect 10329 14448 10332 14500
rect 10280 14324 10283 14376
rect 10283 14324 10329 14376
rect 10329 14324 10332 14376
rect 10280 14200 10283 14252
rect 10283 14200 10329 14252
rect 10329 14200 10332 14252
rect 10280 14076 10283 14128
rect 10283 14076 10329 14128
rect 10329 14076 10332 14128
rect 10280 13952 10283 14004
rect 10283 13952 10329 14004
rect 10329 13952 10332 14004
rect 10280 13828 10283 13880
rect 10283 13828 10329 13880
rect 10329 13828 10332 13880
rect 10280 13704 10283 13756
rect 10283 13704 10329 13756
rect 10329 13704 10332 13756
rect 10280 13580 10283 13632
rect 10283 13580 10329 13632
rect 10329 13580 10332 13632
rect 10280 13456 10283 13508
rect 10283 13456 10329 13508
rect 10329 13456 10332 13508
rect 10280 13332 10283 13384
rect 10283 13332 10329 13384
rect 10329 13332 10332 13384
rect 10280 13208 10283 13260
rect 10283 13208 10329 13260
rect 10329 13208 10332 13260
rect 10280 13084 10283 13136
rect 10283 13084 10329 13136
rect 10329 13084 10332 13136
rect 10280 12960 10283 13012
rect 10283 12960 10329 13012
rect 10329 12960 10332 13012
rect 10280 12836 10283 12888
rect 10283 12836 10329 12888
rect 10329 12836 10332 12888
rect 8040 11757 8092 11758
rect 8040 11706 8043 11757
rect 8043 11706 8089 11757
rect 8089 11706 8092 11757
rect 8040 11582 8043 11634
rect 8043 11582 8089 11634
rect 8089 11582 8092 11634
rect 8040 11458 8043 11510
rect 8043 11458 8089 11510
rect 8089 11458 8092 11510
rect 8488 11757 8540 11758
rect 8488 11706 8491 11757
rect 8491 11706 8537 11757
rect 8537 11706 8540 11757
rect 8488 11582 8491 11634
rect 8491 11582 8537 11634
rect 8537 11582 8540 11634
rect 8488 11458 8491 11510
rect 8491 11458 8537 11510
rect 8537 11458 8540 11510
rect 9848 11859 9900 11911
rect 11624 16602 11676 16654
rect 10952 16478 10955 16530
rect 10955 16478 11001 16530
rect 11001 16478 11004 16530
rect 10952 16354 10955 16406
rect 10955 16354 11001 16406
rect 11001 16354 11004 16406
rect 10952 16230 10955 16282
rect 10955 16230 11001 16282
rect 11001 16230 11004 16282
rect 10952 16106 10955 16158
rect 10955 16106 11001 16158
rect 11001 16106 11004 16158
rect 10952 15982 10955 16034
rect 10955 15982 11001 16034
rect 11001 15982 11004 16034
rect 10952 15858 10955 15910
rect 10955 15858 11001 15910
rect 11001 15858 11004 15910
rect 10952 15734 10955 15786
rect 10955 15734 11001 15786
rect 11001 15734 11004 15786
rect 10952 15610 10955 15662
rect 10955 15610 11001 15662
rect 11001 15610 11004 15662
rect 10952 15486 10955 15538
rect 10955 15486 11001 15538
rect 11001 15486 11004 15538
rect 10728 14944 10731 14996
rect 10731 14944 10777 14996
rect 10777 14944 10780 14996
rect 10728 14820 10731 14872
rect 10731 14820 10777 14872
rect 10777 14820 10780 14872
rect 10728 14696 10731 14748
rect 10731 14696 10777 14748
rect 10777 14696 10780 14748
rect 10728 14572 10731 14624
rect 10731 14572 10777 14624
rect 10777 14572 10780 14624
rect 10728 14448 10731 14500
rect 10731 14448 10777 14500
rect 10777 14448 10780 14500
rect 10728 14324 10731 14376
rect 10731 14324 10777 14376
rect 10777 14324 10780 14376
rect 10728 14200 10731 14252
rect 10731 14200 10777 14252
rect 10777 14200 10780 14252
rect 10728 14076 10731 14128
rect 10731 14076 10777 14128
rect 10777 14076 10780 14128
rect 10728 13952 10731 14004
rect 10731 13952 10777 14004
rect 10777 13952 10780 14004
rect 10728 13828 10731 13880
rect 10731 13828 10777 13880
rect 10777 13828 10780 13880
rect 10728 13704 10731 13756
rect 10731 13704 10777 13756
rect 10777 13704 10780 13756
rect 10728 13580 10731 13632
rect 10731 13580 10777 13632
rect 10777 13580 10780 13632
rect 10728 13456 10731 13508
rect 10731 13456 10777 13508
rect 10777 13456 10780 13508
rect 10728 13332 10731 13384
rect 10731 13332 10777 13384
rect 10777 13332 10780 13384
rect 10728 13208 10731 13260
rect 10731 13208 10777 13260
rect 10777 13208 10780 13260
rect 10728 13084 10731 13136
rect 10731 13084 10777 13136
rect 10777 13084 10780 13136
rect 10728 12960 10731 13012
rect 10731 12960 10777 13012
rect 10777 12960 10780 13012
rect 10728 12836 10731 12888
rect 10731 12836 10777 12888
rect 10777 12836 10780 12888
rect 12072 16602 12124 16654
rect 11624 16478 11627 16530
rect 11627 16478 11673 16530
rect 11673 16478 11676 16530
rect 11624 16354 11627 16406
rect 11627 16354 11673 16406
rect 11673 16354 11676 16406
rect 11624 16230 11627 16282
rect 11627 16230 11673 16282
rect 11673 16230 11676 16282
rect 11624 16106 11627 16158
rect 11627 16106 11673 16158
rect 11673 16106 11676 16158
rect 11624 15982 11627 16034
rect 11627 15982 11673 16034
rect 11673 15982 11676 16034
rect 11624 15858 11627 15910
rect 11627 15858 11673 15910
rect 11673 15858 11676 15910
rect 11624 15734 11627 15786
rect 11627 15734 11673 15786
rect 11673 15734 11676 15786
rect 11624 15610 11627 15662
rect 11627 15610 11673 15662
rect 11673 15610 11676 15662
rect 11624 15486 11627 15538
rect 11627 15486 11673 15538
rect 11673 15486 11676 15538
rect 11400 14944 11403 14996
rect 11403 14944 11449 14996
rect 11449 14944 11452 14996
rect 11400 14820 11403 14872
rect 11403 14820 11449 14872
rect 11449 14820 11452 14872
rect 11400 14696 11403 14748
rect 11403 14696 11449 14748
rect 11449 14696 11452 14748
rect 11400 14572 11403 14624
rect 11403 14572 11449 14624
rect 11449 14572 11452 14624
rect 11400 14448 11403 14500
rect 11403 14448 11449 14500
rect 11449 14448 11452 14500
rect 11400 14324 11403 14376
rect 11403 14324 11449 14376
rect 11449 14324 11452 14376
rect 11400 14200 11403 14252
rect 11403 14200 11449 14252
rect 11449 14200 11452 14252
rect 11400 14076 11403 14128
rect 11403 14076 11449 14128
rect 11449 14076 11452 14128
rect 11400 13952 11403 14004
rect 11403 13952 11449 14004
rect 11449 13952 11452 14004
rect 11400 13828 11403 13880
rect 11403 13828 11449 13880
rect 11449 13828 11452 13880
rect 11400 13704 11403 13756
rect 11403 13704 11449 13756
rect 11449 13704 11452 13756
rect 11400 13580 11403 13632
rect 11403 13580 11449 13632
rect 11449 13580 11452 13632
rect 11400 13456 11403 13508
rect 11403 13456 11449 13508
rect 11449 13456 11452 13508
rect 11400 13332 11403 13384
rect 11403 13332 11449 13384
rect 11449 13332 11452 13384
rect 11400 13208 11403 13260
rect 11403 13208 11449 13260
rect 11449 13208 11452 13260
rect 11400 13084 11403 13136
rect 11403 13084 11449 13136
rect 11449 13084 11452 13136
rect 11400 12960 11403 13012
rect 11403 12960 11449 13012
rect 11449 12960 11452 13012
rect 11400 12836 11403 12888
rect 11403 12836 11449 12888
rect 11449 12836 11452 12888
rect 9160 11757 9212 11758
rect 9160 11706 9163 11757
rect 9163 11706 9209 11757
rect 9209 11706 9212 11757
rect 9160 11582 9163 11634
rect 9163 11582 9209 11634
rect 9209 11582 9212 11634
rect 9160 11458 9163 11510
rect 9163 11458 9209 11510
rect 9209 11458 9212 11510
rect 9608 11757 9660 11758
rect 9608 11706 9611 11757
rect 9611 11706 9657 11757
rect 9657 11706 9660 11757
rect 9608 11582 9611 11634
rect 9611 11582 9657 11634
rect 9657 11582 9660 11634
rect 9608 11458 9611 11510
rect 9611 11458 9657 11510
rect 9657 11458 9660 11510
rect 10968 11859 11020 11911
rect 12744 16602 12796 16654
rect 12072 16478 12075 16530
rect 12075 16478 12121 16530
rect 12121 16478 12124 16530
rect 12072 16354 12075 16406
rect 12075 16354 12121 16406
rect 12121 16354 12124 16406
rect 12072 16230 12075 16282
rect 12075 16230 12121 16282
rect 12121 16230 12124 16282
rect 12072 16106 12075 16158
rect 12075 16106 12121 16158
rect 12121 16106 12124 16158
rect 12072 15982 12075 16034
rect 12075 15982 12121 16034
rect 12121 15982 12124 16034
rect 12072 15858 12075 15910
rect 12075 15858 12121 15910
rect 12121 15858 12124 15910
rect 12072 15734 12075 15786
rect 12075 15734 12121 15786
rect 12121 15734 12124 15786
rect 12072 15610 12075 15662
rect 12075 15610 12121 15662
rect 12121 15610 12124 15662
rect 12072 15486 12075 15538
rect 12075 15486 12121 15538
rect 12121 15486 12124 15538
rect 11848 14944 11851 14996
rect 11851 14944 11897 14996
rect 11897 14944 11900 14996
rect 11848 14820 11851 14872
rect 11851 14820 11897 14872
rect 11897 14820 11900 14872
rect 11848 14696 11851 14748
rect 11851 14696 11897 14748
rect 11897 14696 11900 14748
rect 11848 14572 11851 14624
rect 11851 14572 11897 14624
rect 11897 14572 11900 14624
rect 11848 14448 11851 14500
rect 11851 14448 11897 14500
rect 11897 14448 11900 14500
rect 11848 14324 11851 14376
rect 11851 14324 11897 14376
rect 11897 14324 11900 14376
rect 11848 14200 11851 14252
rect 11851 14200 11897 14252
rect 11897 14200 11900 14252
rect 11848 14076 11851 14128
rect 11851 14076 11897 14128
rect 11897 14076 11900 14128
rect 11848 13952 11851 14004
rect 11851 13952 11897 14004
rect 11897 13952 11900 14004
rect 11848 13828 11851 13880
rect 11851 13828 11897 13880
rect 11897 13828 11900 13880
rect 11848 13704 11851 13756
rect 11851 13704 11897 13756
rect 11897 13704 11900 13756
rect 11848 13580 11851 13632
rect 11851 13580 11897 13632
rect 11897 13580 11900 13632
rect 11848 13456 11851 13508
rect 11851 13456 11897 13508
rect 11897 13456 11900 13508
rect 11848 13332 11851 13384
rect 11851 13332 11897 13384
rect 11897 13332 11900 13384
rect 11848 13208 11851 13260
rect 11851 13208 11897 13260
rect 11897 13208 11900 13260
rect 11848 13084 11851 13136
rect 11851 13084 11897 13136
rect 11897 13084 11900 13136
rect 11848 12960 11851 13012
rect 11851 12960 11897 13012
rect 11897 12960 11900 13012
rect 11848 12836 11851 12888
rect 11851 12836 11897 12888
rect 11897 12836 11900 12888
rect 13192 16602 13244 16654
rect 12744 16478 12747 16530
rect 12747 16478 12793 16530
rect 12793 16478 12796 16530
rect 12744 16354 12747 16406
rect 12747 16354 12793 16406
rect 12793 16354 12796 16406
rect 12744 16230 12747 16282
rect 12747 16230 12793 16282
rect 12793 16230 12796 16282
rect 12744 16106 12747 16158
rect 12747 16106 12793 16158
rect 12793 16106 12796 16158
rect 12744 15982 12747 16034
rect 12747 15982 12793 16034
rect 12793 15982 12796 16034
rect 12744 15858 12747 15910
rect 12747 15858 12793 15910
rect 12793 15858 12796 15910
rect 12744 15734 12747 15786
rect 12747 15734 12793 15786
rect 12793 15734 12796 15786
rect 12744 15610 12747 15662
rect 12747 15610 12793 15662
rect 12793 15610 12796 15662
rect 12744 15486 12747 15538
rect 12747 15486 12793 15538
rect 12793 15486 12796 15538
rect 12520 14944 12523 14996
rect 12523 14944 12569 14996
rect 12569 14944 12572 14996
rect 12520 14820 12523 14872
rect 12523 14820 12569 14872
rect 12569 14820 12572 14872
rect 12520 14696 12523 14748
rect 12523 14696 12569 14748
rect 12569 14696 12572 14748
rect 12520 14572 12523 14624
rect 12523 14572 12569 14624
rect 12569 14572 12572 14624
rect 12520 14448 12523 14500
rect 12523 14448 12569 14500
rect 12569 14448 12572 14500
rect 12520 14324 12523 14376
rect 12523 14324 12569 14376
rect 12569 14324 12572 14376
rect 12520 14200 12523 14252
rect 12523 14200 12569 14252
rect 12569 14200 12572 14252
rect 12520 14076 12523 14128
rect 12523 14076 12569 14128
rect 12569 14076 12572 14128
rect 12520 13952 12523 14004
rect 12523 13952 12569 14004
rect 12569 13952 12572 14004
rect 12520 13828 12523 13880
rect 12523 13828 12569 13880
rect 12569 13828 12572 13880
rect 12520 13704 12523 13756
rect 12523 13704 12569 13756
rect 12569 13704 12572 13756
rect 12520 13580 12523 13632
rect 12523 13580 12569 13632
rect 12569 13580 12572 13632
rect 12520 13456 12523 13508
rect 12523 13456 12569 13508
rect 12569 13456 12572 13508
rect 12520 13332 12523 13384
rect 12523 13332 12569 13384
rect 12569 13332 12572 13384
rect 12520 13208 12523 13260
rect 12523 13208 12569 13260
rect 12569 13208 12572 13260
rect 12520 13084 12523 13136
rect 12523 13084 12569 13136
rect 12569 13084 12572 13136
rect 12520 12960 12523 13012
rect 12523 12960 12569 13012
rect 12569 12960 12572 13012
rect 12520 12836 12523 12888
rect 12523 12836 12569 12888
rect 12569 12836 12572 12888
rect 10280 11757 10332 11758
rect 10280 11706 10283 11757
rect 10283 11706 10329 11757
rect 10329 11706 10332 11757
rect 10280 11582 10283 11634
rect 10283 11582 10329 11634
rect 10329 11582 10332 11634
rect 10280 11458 10283 11510
rect 10283 11458 10329 11510
rect 10329 11458 10332 11510
rect 10728 11757 10780 11758
rect 10728 11706 10731 11757
rect 10731 11706 10777 11757
rect 10777 11706 10780 11757
rect 10728 11582 10731 11634
rect 10731 11582 10777 11634
rect 10777 11582 10780 11634
rect 10728 11458 10731 11510
rect 10731 11458 10777 11510
rect 10777 11458 10780 11510
rect 12088 11859 12140 11911
rect 13864 16602 13916 16654
rect 13192 16478 13195 16530
rect 13195 16478 13241 16530
rect 13241 16478 13244 16530
rect 13192 16354 13195 16406
rect 13195 16354 13241 16406
rect 13241 16354 13244 16406
rect 13192 16230 13195 16282
rect 13195 16230 13241 16282
rect 13241 16230 13244 16282
rect 13192 16106 13195 16158
rect 13195 16106 13241 16158
rect 13241 16106 13244 16158
rect 13192 15982 13195 16034
rect 13195 15982 13241 16034
rect 13241 15982 13244 16034
rect 13192 15858 13195 15910
rect 13195 15858 13241 15910
rect 13241 15858 13244 15910
rect 13192 15734 13195 15786
rect 13195 15734 13241 15786
rect 13241 15734 13244 15786
rect 13192 15610 13195 15662
rect 13195 15610 13241 15662
rect 13241 15610 13244 15662
rect 13192 15486 13195 15538
rect 13195 15486 13241 15538
rect 13241 15486 13244 15538
rect 12968 14944 12971 14996
rect 12971 14944 13017 14996
rect 13017 14944 13020 14996
rect 12968 14820 12971 14872
rect 12971 14820 13017 14872
rect 13017 14820 13020 14872
rect 12968 14696 12971 14748
rect 12971 14696 13017 14748
rect 13017 14696 13020 14748
rect 12968 14572 12971 14624
rect 12971 14572 13017 14624
rect 13017 14572 13020 14624
rect 12968 14448 12971 14500
rect 12971 14448 13017 14500
rect 13017 14448 13020 14500
rect 12968 14324 12971 14376
rect 12971 14324 13017 14376
rect 13017 14324 13020 14376
rect 12968 14200 12971 14252
rect 12971 14200 13017 14252
rect 13017 14200 13020 14252
rect 12968 14076 12971 14128
rect 12971 14076 13017 14128
rect 13017 14076 13020 14128
rect 12968 13952 12971 14004
rect 12971 13952 13017 14004
rect 13017 13952 13020 14004
rect 12968 13828 12971 13880
rect 12971 13828 13017 13880
rect 13017 13828 13020 13880
rect 12968 13704 12971 13756
rect 12971 13704 13017 13756
rect 13017 13704 13020 13756
rect 12968 13580 12971 13632
rect 12971 13580 13017 13632
rect 13017 13580 13020 13632
rect 12968 13456 12971 13508
rect 12971 13456 13017 13508
rect 13017 13456 13020 13508
rect 12968 13332 12971 13384
rect 12971 13332 13017 13384
rect 13017 13332 13020 13384
rect 12968 13208 12971 13260
rect 12971 13208 13017 13260
rect 13017 13208 13020 13260
rect 12968 13084 12971 13136
rect 12971 13084 13017 13136
rect 13017 13084 13020 13136
rect 12968 12960 12971 13012
rect 12971 12960 13017 13012
rect 13017 12960 13020 13012
rect 12968 12836 12971 12888
rect 12971 12836 13017 12888
rect 13017 12836 13020 12888
rect 14312 16602 14364 16654
rect 13864 16478 13867 16530
rect 13867 16478 13913 16530
rect 13913 16478 13916 16530
rect 13864 16354 13867 16406
rect 13867 16354 13913 16406
rect 13913 16354 13916 16406
rect 13864 16230 13867 16282
rect 13867 16230 13913 16282
rect 13913 16230 13916 16282
rect 13864 16106 13867 16158
rect 13867 16106 13913 16158
rect 13913 16106 13916 16158
rect 13864 15982 13867 16034
rect 13867 15982 13913 16034
rect 13913 15982 13916 16034
rect 13864 15858 13867 15910
rect 13867 15858 13913 15910
rect 13913 15858 13916 15910
rect 13864 15734 13867 15786
rect 13867 15734 13913 15786
rect 13913 15734 13916 15786
rect 13864 15610 13867 15662
rect 13867 15610 13913 15662
rect 13913 15610 13916 15662
rect 13864 15486 13867 15538
rect 13867 15486 13913 15538
rect 13913 15486 13916 15538
rect 13640 14944 13643 14996
rect 13643 14944 13689 14996
rect 13689 14944 13692 14996
rect 13640 14820 13643 14872
rect 13643 14820 13689 14872
rect 13689 14820 13692 14872
rect 13640 14696 13643 14748
rect 13643 14696 13689 14748
rect 13689 14696 13692 14748
rect 13640 14572 13643 14624
rect 13643 14572 13689 14624
rect 13689 14572 13692 14624
rect 13640 14448 13643 14500
rect 13643 14448 13689 14500
rect 13689 14448 13692 14500
rect 13640 14324 13643 14376
rect 13643 14324 13689 14376
rect 13689 14324 13692 14376
rect 13640 14200 13643 14252
rect 13643 14200 13689 14252
rect 13689 14200 13692 14252
rect 13640 14076 13643 14128
rect 13643 14076 13689 14128
rect 13689 14076 13692 14128
rect 13640 13952 13643 14004
rect 13643 13952 13689 14004
rect 13689 13952 13692 14004
rect 13640 13828 13643 13880
rect 13643 13828 13689 13880
rect 13689 13828 13692 13880
rect 13640 13704 13643 13756
rect 13643 13704 13689 13756
rect 13689 13704 13692 13756
rect 13640 13580 13643 13632
rect 13643 13580 13689 13632
rect 13689 13580 13692 13632
rect 13640 13456 13643 13508
rect 13643 13456 13689 13508
rect 13689 13456 13692 13508
rect 13640 13332 13643 13384
rect 13643 13332 13689 13384
rect 13689 13332 13692 13384
rect 13640 13208 13643 13260
rect 13643 13208 13689 13260
rect 13689 13208 13692 13260
rect 13640 13084 13643 13136
rect 13643 13084 13689 13136
rect 13689 13084 13692 13136
rect 13640 12960 13643 13012
rect 13643 12960 13689 13012
rect 13689 12960 13692 13012
rect 13640 12836 13643 12888
rect 13643 12836 13689 12888
rect 13689 12836 13692 12888
rect 11400 11757 11452 11758
rect 11400 11706 11403 11757
rect 11403 11706 11449 11757
rect 11449 11706 11452 11757
rect 11400 11582 11403 11634
rect 11403 11582 11449 11634
rect 11449 11582 11452 11634
rect 11400 11458 11403 11510
rect 11403 11458 11449 11510
rect 11449 11458 11452 11510
rect 11848 11757 11900 11758
rect 11848 11706 11851 11757
rect 11851 11706 11897 11757
rect 11897 11706 11900 11757
rect 11848 11582 11851 11634
rect 11851 11582 11897 11634
rect 11897 11582 11900 11634
rect 11848 11458 11851 11510
rect 11851 11458 11897 11510
rect 11897 11458 11900 11510
rect 13208 11859 13260 11911
rect 14984 16602 15036 16654
rect 14312 16478 14315 16530
rect 14315 16478 14361 16530
rect 14361 16478 14364 16530
rect 14312 16354 14315 16406
rect 14315 16354 14361 16406
rect 14361 16354 14364 16406
rect 14312 16230 14315 16282
rect 14315 16230 14361 16282
rect 14361 16230 14364 16282
rect 14312 16106 14315 16158
rect 14315 16106 14361 16158
rect 14361 16106 14364 16158
rect 14312 15982 14315 16034
rect 14315 15982 14361 16034
rect 14361 15982 14364 16034
rect 14312 15858 14315 15910
rect 14315 15858 14361 15910
rect 14361 15858 14364 15910
rect 14312 15734 14315 15786
rect 14315 15734 14361 15786
rect 14361 15734 14364 15786
rect 14312 15610 14315 15662
rect 14315 15610 14361 15662
rect 14361 15610 14364 15662
rect 14312 15486 14315 15538
rect 14315 15486 14361 15538
rect 14361 15486 14364 15538
rect 14088 14944 14091 14996
rect 14091 14944 14137 14996
rect 14137 14944 14140 14996
rect 14088 14820 14091 14872
rect 14091 14820 14137 14872
rect 14137 14820 14140 14872
rect 14088 14696 14091 14748
rect 14091 14696 14137 14748
rect 14137 14696 14140 14748
rect 14088 14572 14091 14624
rect 14091 14572 14137 14624
rect 14137 14572 14140 14624
rect 14088 14448 14091 14500
rect 14091 14448 14137 14500
rect 14137 14448 14140 14500
rect 14088 14324 14091 14376
rect 14091 14324 14137 14376
rect 14137 14324 14140 14376
rect 14088 14200 14091 14252
rect 14091 14200 14137 14252
rect 14137 14200 14140 14252
rect 14088 14076 14091 14128
rect 14091 14076 14137 14128
rect 14137 14076 14140 14128
rect 14088 13952 14091 14004
rect 14091 13952 14137 14004
rect 14137 13952 14140 14004
rect 14088 13828 14091 13880
rect 14091 13828 14137 13880
rect 14137 13828 14140 13880
rect 14088 13704 14091 13756
rect 14091 13704 14137 13756
rect 14137 13704 14140 13756
rect 14088 13580 14091 13632
rect 14091 13580 14137 13632
rect 14137 13580 14140 13632
rect 14088 13456 14091 13508
rect 14091 13456 14137 13508
rect 14137 13456 14140 13508
rect 14088 13332 14091 13384
rect 14091 13332 14137 13384
rect 14137 13332 14140 13384
rect 14088 13208 14091 13260
rect 14091 13208 14137 13260
rect 14137 13208 14140 13260
rect 14088 13084 14091 13136
rect 14091 13084 14137 13136
rect 14137 13084 14140 13136
rect 14088 12960 14091 13012
rect 14091 12960 14137 13012
rect 14137 12960 14140 13012
rect 14088 12836 14091 12888
rect 14091 12836 14137 12888
rect 14137 12836 14140 12888
rect 15432 16602 15484 16654
rect 14984 16478 14987 16530
rect 14987 16478 15033 16530
rect 15033 16478 15036 16530
rect 14984 16354 14987 16406
rect 14987 16354 15033 16406
rect 15033 16354 15036 16406
rect 14984 16230 14987 16282
rect 14987 16230 15033 16282
rect 15033 16230 15036 16282
rect 14984 16106 14987 16158
rect 14987 16106 15033 16158
rect 15033 16106 15036 16158
rect 14984 15982 14987 16034
rect 14987 15982 15033 16034
rect 15033 15982 15036 16034
rect 14984 15858 14987 15910
rect 14987 15858 15033 15910
rect 15033 15858 15036 15910
rect 14984 15734 14987 15786
rect 14987 15734 15033 15786
rect 15033 15734 15036 15786
rect 14984 15610 14987 15662
rect 14987 15610 15033 15662
rect 15033 15610 15036 15662
rect 14984 15486 14987 15538
rect 14987 15486 15033 15538
rect 15033 15486 15036 15538
rect 14760 14944 14763 14996
rect 14763 14944 14809 14996
rect 14809 14944 14812 14996
rect 14760 14820 14763 14872
rect 14763 14820 14809 14872
rect 14809 14820 14812 14872
rect 14760 14696 14763 14748
rect 14763 14696 14809 14748
rect 14809 14696 14812 14748
rect 14760 14572 14763 14624
rect 14763 14572 14809 14624
rect 14809 14572 14812 14624
rect 14760 14448 14763 14500
rect 14763 14448 14809 14500
rect 14809 14448 14812 14500
rect 14760 14324 14763 14376
rect 14763 14324 14809 14376
rect 14809 14324 14812 14376
rect 14760 14200 14763 14252
rect 14763 14200 14809 14252
rect 14809 14200 14812 14252
rect 14760 14076 14763 14128
rect 14763 14076 14809 14128
rect 14809 14076 14812 14128
rect 14760 13952 14763 14004
rect 14763 13952 14809 14004
rect 14809 13952 14812 14004
rect 14760 13828 14763 13880
rect 14763 13828 14809 13880
rect 14809 13828 14812 13880
rect 14760 13704 14763 13756
rect 14763 13704 14809 13756
rect 14809 13704 14812 13756
rect 14760 13580 14763 13632
rect 14763 13580 14809 13632
rect 14809 13580 14812 13632
rect 14760 13456 14763 13508
rect 14763 13456 14809 13508
rect 14809 13456 14812 13508
rect 14760 13332 14763 13384
rect 14763 13332 14809 13384
rect 14809 13332 14812 13384
rect 14760 13208 14763 13260
rect 14763 13208 14809 13260
rect 14809 13208 14812 13260
rect 14760 13084 14763 13136
rect 14763 13084 14809 13136
rect 14809 13084 14812 13136
rect 14760 12960 14763 13012
rect 14763 12960 14809 13012
rect 14809 12960 14812 13012
rect 14760 12836 14763 12888
rect 14763 12836 14809 12888
rect 14809 12836 14812 12888
rect 12520 11757 12572 11758
rect 12520 11706 12523 11757
rect 12523 11706 12569 11757
rect 12569 11706 12572 11757
rect 12520 11582 12523 11634
rect 12523 11582 12569 11634
rect 12569 11582 12572 11634
rect 12520 11458 12523 11510
rect 12523 11458 12569 11510
rect 12569 11458 12572 11510
rect 12968 11757 13020 11758
rect 12968 11706 12971 11757
rect 12971 11706 13017 11757
rect 13017 11706 13020 11757
rect 12968 11582 12971 11634
rect 12971 11582 13017 11634
rect 13017 11582 13020 11634
rect 12968 11458 12971 11510
rect 12971 11458 13017 11510
rect 13017 11458 13020 11510
rect 14328 11859 14380 11911
rect 16104 16602 16156 16654
rect 15432 16478 15435 16530
rect 15435 16478 15481 16530
rect 15481 16478 15484 16530
rect 15432 16354 15435 16406
rect 15435 16354 15481 16406
rect 15481 16354 15484 16406
rect 15432 16230 15435 16282
rect 15435 16230 15481 16282
rect 15481 16230 15484 16282
rect 15432 16106 15435 16158
rect 15435 16106 15481 16158
rect 15481 16106 15484 16158
rect 15432 15982 15435 16034
rect 15435 15982 15481 16034
rect 15481 15982 15484 16034
rect 15432 15858 15435 15910
rect 15435 15858 15481 15910
rect 15481 15858 15484 15910
rect 15432 15734 15435 15786
rect 15435 15734 15481 15786
rect 15481 15734 15484 15786
rect 15432 15610 15435 15662
rect 15435 15610 15481 15662
rect 15481 15610 15484 15662
rect 15432 15486 15435 15538
rect 15435 15486 15481 15538
rect 15481 15486 15484 15538
rect 15208 14944 15211 14996
rect 15211 14944 15257 14996
rect 15257 14944 15260 14996
rect 15208 14820 15211 14872
rect 15211 14820 15257 14872
rect 15257 14820 15260 14872
rect 15208 14696 15211 14748
rect 15211 14696 15257 14748
rect 15257 14696 15260 14748
rect 15208 14572 15211 14624
rect 15211 14572 15257 14624
rect 15257 14572 15260 14624
rect 15208 14448 15211 14500
rect 15211 14448 15257 14500
rect 15257 14448 15260 14500
rect 15208 14324 15211 14376
rect 15211 14324 15257 14376
rect 15257 14324 15260 14376
rect 15208 14200 15211 14252
rect 15211 14200 15257 14252
rect 15257 14200 15260 14252
rect 15208 14076 15211 14128
rect 15211 14076 15257 14128
rect 15257 14076 15260 14128
rect 15208 13952 15211 14004
rect 15211 13952 15257 14004
rect 15257 13952 15260 14004
rect 15208 13828 15211 13880
rect 15211 13828 15257 13880
rect 15257 13828 15260 13880
rect 15208 13704 15211 13756
rect 15211 13704 15257 13756
rect 15257 13704 15260 13756
rect 15208 13580 15211 13632
rect 15211 13580 15257 13632
rect 15257 13580 15260 13632
rect 15208 13456 15211 13508
rect 15211 13456 15257 13508
rect 15257 13456 15260 13508
rect 15208 13332 15211 13384
rect 15211 13332 15257 13384
rect 15257 13332 15260 13384
rect 15208 13208 15211 13260
rect 15211 13208 15257 13260
rect 15257 13208 15260 13260
rect 15208 13084 15211 13136
rect 15211 13084 15257 13136
rect 15257 13084 15260 13136
rect 15208 12960 15211 13012
rect 15211 12960 15257 13012
rect 15257 12960 15260 13012
rect 15208 12836 15211 12888
rect 15211 12836 15257 12888
rect 15257 12836 15260 12888
rect 16552 16602 16604 16654
rect 16104 16478 16107 16530
rect 16107 16478 16153 16530
rect 16153 16478 16156 16530
rect 16104 16354 16107 16406
rect 16107 16354 16153 16406
rect 16153 16354 16156 16406
rect 16104 16230 16107 16282
rect 16107 16230 16153 16282
rect 16153 16230 16156 16282
rect 16104 16106 16107 16158
rect 16107 16106 16153 16158
rect 16153 16106 16156 16158
rect 16104 15982 16107 16034
rect 16107 15982 16153 16034
rect 16153 15982 16156 16034
rect 16104 15858 16107 15910
rect 16107 15858 16153 15910
rect 16153 15858 16156 15910
rect 16104 15734 16107 15786
rect 16107 15734 16153 15786
rect 16153 15734 16156 15786
rect 16104 15610 16107 15662
rect 16107 15610 16153 15662
rect 16153 15610 16156 15662
rect 16104 15486 16107 15538
rect 16107 15486 16153 15538
rect 16153 15486 16156 15538
rect 15880 14944 15883 14996
rect 15883 14944 15929 14996
rect 15929 14944 15932 14996
rect 15880 14820 15883 14872
rect 15883 14820 15929 14872
rect 15929 14820 15932 14872
rect 15880 14696 15883 14748
rect 15883 14696 15929 14748
rect 15929 14696 15932 14748
rect 15880 14572 15883 14624
rect 15883 14572 15929 14624
rect 15929 14572 15932 14624
rect 15880 14448 15883 14500
rect 15883 14448 15929 14500
rect 15929 14448 15932 14500
rect 15880 14324 15883 14376
rect 15883 14324 15929 14376
rect 15929 14324 15932 14376
rect 15880 14200 15883 14252
rect 15883 14200 15929 14252
rect 15929 14200 15932 14252
rect 15880 14076 15883 14128
rect 15883 14076 15929 14128
rect 15929 14076 15932 14128
rect 15880 13952 15883 14004
rect 15883 13952 15929 14004
rect 15929 13952 15932 14004
rect 15880 13828 15883 13880
rect 15883 13828 15929 13880
rect 15929 13828 15932 13880
rect 15880 13704 15883 13756
rect 15883 13704 15929 13756
rect 15929 13704 15932 13756
rect 15880 13580 15883 13632
rect 15883 13580 15929 13632
rect 15929 13580 15932 13632
rect 15880 13456 15883 13508
rect 15883 13456 15929 13508
rect 15929 13456 15932 13508
rect 15880 13332 15883 13384
rect 15883 13332 15929 13384
rect 15929 13332 15932 13384
rect 15880 13208 15883 13260
rect 15883 13208 15929 13260
rect 15929 13208 15932 13260
rect 15880 13084 15883 13136
rect 15883 13084 15929 13136
rect 15929 13084 15932 13136
rect 15880 12960 15883 13012
rect 15883 12960 15929 13012
rect 15929 12960 15932 13012
rect 15880 12836 15883 12888
rect 15883 12836 15929 12888
rect 15929 12836 15932 12888
rect 13640 11757 13692 11758
rect 13640 11706 13643 11757
rect 13643 11706 13689 11757
rect 13689 11706 13692 11757
rect 13640 11582 13643 11634
rect 13643 11582 13689 11634
rect 13689 11582 13692 11634
rect 13640 11458 13643 11510
rect 13643 11458 13689 11510
rect 13689 11458 13692 11510
rect 14088 11757 14140 11758
rect 14088 11706 14091 11757
rect 14091 11706 14137 11757
rect 14137 11706 14140 11757
rect 14088 11582 14091 11634
rect 14091 11582 14137 11634
rect 14137 11582 14140 11634
rect 14088 11458 14091 11510
rect 14091 11458 14137 11510
rect 14137 11458 14140 11510
rect 15448 11859 15500 11911
rect 17224 16602 17276 16654
rect 16552 16478 16555 16530
rect 16555 16478 16601 16530
rect 16601 16478 16604 16530
rect 16552 16354 16555 16406
rect 16555 16354 16601 16406
rect 16601 16354 16604 16406
rect 16552 16230 16555 16282
rect 16555 16230 16601 16282
rect 16601 16230 16604 16282
rect 16552 16106 16555 16158
rect 16555 16106 16601 16158
rect 16601 16106 16604 16158
rect 16552 15982 16555 16034
rect 16555 15982 16601 16034
rect 16601 15982 16604 16034
rect 16552 15858 16555 15910
rect 16555 15858 16601 15910
rect 16601 15858 16604 15910
rect 16552 15734 16555 15786
rect 16555 15734 16601 15786
rect 16601 15734 16604 15786
rect 16552 15610 16555 15662
rect 16555 15610 16601 15662
rect 16601 15610 16604 15662
rect 16552 15486 16555 15538
rect 16555 15486 16601 15538
rect 16601 15486 16604 15538
rect 16328 14944 16331 14996
rect 16331 14944 16377 14996
rect 16377 14944 16380 14996
rect 16328 14820 16331 14872
rect 16331 14820 16377 14872
rect 16377 14820 16380 14872
rect 16328 14696 16331 14748
rect 16331 14696 16377 14748
rect 16377 14696 16380 14748
rect 16328 14572 16331 14624
rect 16331 14572 16377 14624
rect 16377 14572 16380 14624
rect 16328 14448 16331 14500
rect 16331 14448 16377 14500
rect 16377 14448 16380 14500
rect 16328 14324 16331 14376
rect 16331 14324 16377 14376
rect 16377 14324 16380 14376
rect 16328 14200 16331 14252
rect 16331 14200 16377 14252
rect 16377 14200 16380 14252
rect 16328 14076 16331 14128
rect 16331 14076 16377 14128
rect 16377 14076 16380 14128
rect 16328 13952 16331 14004
rect 16331 13952 16377 14004
rect 16377 13952 16380 14004
rect 16328 13828 16331 13880
rect 16331 13828 16377 13880
rect 16377 13828 16380 13880
rect 16328 13704 16331 13756
rect 16331 13704 16377 13756
rect 16377 13704 16380 13756
rect 16328 13580 16331 13632
rect 16331 13580 16377 13632
rect 16377 13580 16380 13632
rect 16328 13456 16331 13508
rect 16331 13456 16377 13508
rect 16377 13456 16380 13508
rect 16328 13332 16331 13384
rect 16331 13332 16377 13384
rect 16377 13332 16380 13384
rect 16328 13208 16331 13260
rect 16331 13208 16377 13260
rect 16377 13208 16380 13260
rect 16328 13084 16331 13136
rect 16331 13084 16377 13136
rect 16377 13084 16380 13136
rect 16328 12960 16331 13012
rect 16331 12960 16377 13012
rect 16377 12960 16380 13012
rect 16328 12836 16331 12888
rect 16331 12836 16377 12888
rect 16377 12836 16380 12888
rect 17672 16602 17724 16654
rect 17224 16478 17227 16530
rect 17227 16478 17273 16530
rect 17273 16478 17276 16530
rect 17224 16354 17227 16406
rect 17227 16354 17273 16406
rect 17273 16354 17276 16406
rect 17224 16230 17227 16282
rect 17227 16230 17273 16282
rect 17273 16230 17276 16282
rect 17224 16106 17227 16158
rect 17227 16106 17273 16158
rect 17273 16106 17276 16158
rect 17224 15982 17227 16034
rect 17227 15982 17273 16034
rect 17273 15982 17276 16034
rect 17224 15858 17227 15910
rect 17227 15858 17273 15910
rect 17273 15858 17276 15910
rect 17224 15734 17227 15786
rect 17227 15734 17273 15786
rect 17273 15734 17276 15786
rect 17224 15610 17227 15662
rect 17227 15610 17273 15662
rect 17273 15610 17276 15662
rect 17224 15486 17227 15538
rect 17227 15486 17273 15538
rect 17273 15486 17276 15538
rect 17000 14944 17003 14996
rect 17003 14944 17049 14996
rect 17049 14944 17052 14996
rect 17000 14820 17003 14872
rect 17003 14820 17049 14872
rect 17049 14820 17052 14872
rect 17000 14696 17003 14748
rect 17003 14696 17049 14748
rect 17049 14696 17052 14748
rect 17000 14572 17003 14624
rect 17003 14572 17049 14624
rect 17049 14572 17052 14624
rect 17000 14448 17003 14500
rect 17003 14448 17049 14500
rect 17049 14448 17052 14500
rect 17000 14324 17003 14376
rect 17003 14324 17049 14376
rect 17049 14324 17052 14376
rect 17000 14200 17003 14252
rect 17003 14200 17049 14252
rect 17049 14200 17052 14252
rect 17000 14076 17003 14128
rect 17003 14076 17049 14128
rect 17049 14076 17052 14128
rect 17000 13952 17003 14004
rect 17003 13952 17049 14004
rect 17049 13952 17052 14004
rect 17000 13828 17003 13880
rect 17003 13828 17049 13880
rect 17049 13828 17052 13880
rect 17000 13704 17003 13756
rect 17003 13704 17049 13756
rect 17049 13704 17052 13756
rect 17000 13580 17003 13632
rect 17003 13580 17049 13632
rect 17049 13580 17052 13632
rect 17000 13456 17003 13508
rect 17003 13456 17049 13508
rect 17049 13456 17052 13508
rect 17000 13332 17003 13384
rect 17003 13332 17049 13384
rect 17049 13332 17052 13384
rect 17000 13208 17003 13260
rect 17003 13208 17049 13260
rect 17049 13208 17052 13260
rect 17000 13084 17003 13136
rect 17003 13084 17049 13136
rect 17049 13084 17052 13136
rect 17000 12960 17003 13012
rect 17003 12960 17049 13012
rect 17049 12960 17052 13012
rect 17000 12836 17003 12888
rect 17003 12836 17049 12888
rect 17049 12836 17052 12888
rect 14760 11757 14812 11758
rect 14760 11706 14763 11757
rect 14763 11706 14809 11757
rect 14809 11706 14812 11757
rect 14760 11582 14763 11634
rect 14763 11582 14809 11634
rect 14809 11582 14812 11634
rect 14760 11458 14763 11510
rect 14763 11458 14809 11510
rect 14809 11458 14812 11510
rect 15208 11757 15260 11758
rect 15208 11706 15211 11757
rect 15211 11706 15257 11757
rect 15257 11706 15260 11757
rect 15208 11582 15211 11634
rect 15211 11582 15257 11634
rect 15257 11582 15260 11634
rect 15208 11458 15211 11510
rect 15211 11458 15257 11510
rect 15257 11458 15260 11510
rect 16568 11859 16620 11911
rect 18344 16602 18396 16654
rect 17672 16478 17675 16530
rect 17675 16478 17721 16530
rect 17721 16478 17724 16530
rect 17672 16354 17675 16406
rect 17675 16354 17721 16406
rect 17721 16354 17724 16406
rect 17672 16230 17675 16282
rect 17675 16230 17721 16282
rect 17721 16230 17724 16282
rect 17672 16106 17675 16158
rect 17675 16106 17721 16158
rect 17721 16106 17724 16158
rect 17672 15982 17675 16034
rect 17675 15982 17721 16034
rect 17721 15982 17724 16034
rect 17672 15858 17675 15910
rect 17675 15858 17721 15910
rect 17721 15858 17724 15910
rect 17672 15734 17675 15786
rect 17675 15734 17721 15786
rect 17721 15734 17724 15786
rect 17672 15610 17675 15662
rect 17675 15610 17721 15662
rect 17721 15610 17724 15662
rect 17672 15486 17675 15538
rect 17675 15486 17721 15538
rect 17721 15486 17724 15538
rect 17448 14944 17451 14996
rect 17451 14944 17497 14996
rect 17497 14944 17500 14996
rect 17448 14820 17451 14872
rect 17451 14820 17497 14872
rect 17497 14820 17500 14872
rect 17448 14696 17451 14748
rect 17451 14696 17497 14748
rect 17497 14696 17500 14748
rect 17448 14572 17451 14624
rect 17451 14572 17497 14624
rect 17497 14572 17500 14624
rect 17448 14448 17451 14500
rect 17451 14448 17497 14500
rect 17497 14448 17500 14500
rect 17448 14324 17451 14376
rect 17451 14324 17497 14376
rect 17497 14324 17500 14376
rect 17448 14200 17451 14252
rect 17451 14200 17497 14252
rect 17497 14200 17500 14252
rect 17448 14076 17451 14128
rect 17451 14076 17497 14128
rect 17497 14076 17500 14128
rect 17448 13952 17451 14004
rect 17451 13952 17497 14004
rect 17497 13952 17500 14004
rect 17448 13828 17451 13880
rect 17451 13828 17497 13880
rect 17497 13828 17500 13880
rect 17448 13704 17451 13756
rect 17451 13704 17497 13756
rect 17497 13704 17500 13756
rect 17448 13580 17451 13632
rect 17451 13580 17497 13632
rect 17497 13580 17500 13632
rect 17448 13456 17451 13508
rect 17451 13456 17497 13508
rect 17497 13456 17500 13508
rect 17448 13332 17451 13384
rect 17451 13332 17497 13384
rect 17497 13332 17500 13384
rect 17448 13208 17451 13260
rect 17451 13208 17497 13260
rect 17497 13208 17500 13260
rect 17448 13084 17451 13136
rect 17451 13084 17497 13136
rect 17497 13084 17500 13136
rect 17448 12960 17451 13012
rect 17451 12960 17497 13012
rect 17497 12960 17500 13012
rect 17448 12836 17451 12888
rect 17451 12836 17497 12888
rect 17497 12836 17500 12888
rect 18792 16602 18844 16654
rect 18344 16478 18347 16530
rect 18347 16478 18393 16530
rect 18393 16478 18396 16530
rect 18344 16354 18347 16406
rect 18347 16354 18393 16406
rect 18393 16354 18396 16406
rect 18344 16230 18347 16282
rect 18347 16230 18393 16282
rect 18393 16230 18396 16282
rect 18344 16106 18347 16158
rect 18347 16106 18393 16158
rect 18393 16106 18396 16158
rect 18344 15982 18347 16034
rect 18347 15982 18393 16034
rect 18393 15982 18396 16034
rect 18344 15858 18347 15910
rect 18347 15858 18393 15910
rect 18393 15858 18396 15910
rect 18344 15734 18347 15786
rect 18347 15734 18393 15786
rect 18393 15734 18396 15786
rect 18344 15610 18347 15662
rect 18347 15610 18393 15662
rect 18393 15610 18396 15662
rect 18344 15486 18347 15538
rect 18347 15486 18393 15538
rect 18393 15486 18396 15538
rect 18120 14944 18123 14996
rect 18123 14944 18169 14996
rect 18169 14944 18172 14996
rect 18120 14820 18123 14872
rect 18123 14820 18169 14872
rect 18169 14820 18172 14872
rect 18120 14696 18123 14748
rect 18123 14696 18169 14748
rect 18169 14696 18172 14748
rect 18120 14572 18123 14624
rect 18123 14572 18169 14624
rect 18169 14572 18172 14624
rect 18120 14448 18123 14500
rect 18123 14448 18169 14500
rect 18169 14448 18172 14500
rect 18120 14324 18123 14376
rect 18123 14324 18169 14376
rect 18169 14324 18172 14376
rect 18120 14200 18123 14252
rect 18123 14200 18169 14252
rect 18169 14200 18172 14252
rect 18120 14076 18123 14128
rect 18123 14076 18169 14128
rect 18169 14076 18172 14128
rect 18120 13952 18123 14004
rect 18123 13952 18169 14004
rect 18169 13952 18172 14004
rect 18120 13828 18123 13880
rect 18123 13828 18169 13880
rect 18169 13828 18172 13880
rect 18120 13704 18123 13756
rect 18123 13704 18169 13756
rect 18169 13704 18172 13756
rect 18120 13580 18123 13632
rect 18123 13580 18169 13632
rect 18169 13580 18172 13632
rect 18120 13456 18123 13508
rect 18123 13456 18169 13508
rect 18169 13456 18172 13508
rect 18120 13332 18123 13384
rect 18123 13332 18169 13384
rect 18169 13332 18172 13384
rect 18120 13208 18123 13260
rect 18123 13208 18169 13260
rect 18169 13208 18172 13260
rect 18120 13084 18123 13136
rect 18123 13084 18169 13136
rect 18169 13084 18172 13136
rect 18120 12960 18123 13012
rect 18123 12960 18169 13012
rect 18169 12960 18172 13012
rect 18120 12836 18123 12888
rect 18123 12836 18169 12888
rect 18169 12836 18172 12888
rect 15880 11757 15932 11758
rect 15880 11706 15883 11757
rect 15883 11706 15929 11757
rect 15929 11706 15932 11757
rect 15880 11582 15883 11634
rect 15883 11582 15929 11634
rect 15929 11582 15932 11634
rect 15880 11458 15883 11510
rect 15883 11458 15929 11510
rect 15929 11458 15932 11510
rect 16328 11757 16380 11758
rect 16328 11706 16331 11757
rect 16331 11706 16377 11757
rect 16377 11706 16380 11757
rect 16328 11582 16331 11634
rect 16331 11582 16377 11634
rect 16377 11582 16380 11634
rect 16328 11458 16331 11510
rect 16331 11458 16377 11510
rect 16377 11458 16380 11510
rect 17688 11859 17740 11911
rect 19464 16602 19516 16654
rect 18792 16478 18795 16530
rect 18795 16478 18841 16530
rect 18841 16478 18844 16530
rect 18792 16354 18795 16406
rect 18795 16354 18841 16406
rect 18841 16354 18844 16406
rect 18792 16230 18795 16282
rect 18795 16230 18841 16282
rect 18841 16230 18844 16282
rect 18792 16106 18795 16158
rect 18795 16106 18841 16158
rect 18841 16106 18844 16158
rect 18792 15982 18795 16034
rect 18795 15982 18841 16034
rect 18841 15982 18844 16034
rect 18792 15858 18795 15910
rect 18795 15858 18841 15910
rect 18841 15858 18844 15910
rect 18792 15734 18795 15786
rect 18795 15734 18841 15786
rect 18841 15734 18844 15786
rect 18792 15610 18795 15662
rect 18795 15610 18841 15662
rect 18841 15610 18844 15662
rect 18792 15486 18795 15538
rect 18795 15486 18841 15538
rect 18841 15486 18844 15538
rect 18568 14944 18571 14996
rect 18571 14944 18617 14996
rect 18617 14944 18620 14996
rect 18568 14820 18571 14872
rect 18571 14820 18617 14872
rect 18617 14820 18620 14872
rect 18568 14696 18571 14748
rect 18571 14696 18617 14748
rect 18617 14696 18620 14748
rect 18568 14572 18571 14624
rect 18571 14572 18617 14624
rect 18617 14572 18620 14624
rect 18568 14448 18571 14500
rect 18571 14448 18617 14500
rect 18617 14448 18620 14500
rect 18568 14324 18571 14376
rect 18571 14324 18617 14376
rect 18617 14324 18620 14376
rect 18568 14200 18571 14252
rect 18571 14200 18617 14252
rect 18617 14200 18620 14252
rect 18568 14076 18571 14128
rect 18571 14076 18617 14128
rect 18617 14076 18620 14128
rect 18568 13952 18571 14004
rect 18571 13952 18617 14004
rect 18617 13952 18620 14004
rect 18568 13828 18571 13880
rect 18571 13828 18617 13880
rect 18617 13828 18620 13880
rect 18568 13704 18571 13756
rect 18571 13704 18617 13756
rect 18617 13704 18620 13756
rect 18568 13580 18571 13632
rect 18571 13580 18617 13632
rect 18617 13580 18620 13632
rect 18568 13456 18571 13508
rect 18571 13456 18617 13508
rect 18617 13456 18620 13508
rect 18568 13332 18571 13384
rect 18571 13332 18617 13384
rect 18617 13332 18620 13384
rect 18568 13208 18571 13260
rect 18571 13208 18617 13260
rect 18617 13208 18620 13260
rect 18568 13084 18571 13136
rect 18571 13084 18617 13136
rect 18617 13084 18620 13136
rect 18568 12960 18571 13012
rect 18571 12960 18617 13012
rect 18617 12960 18620 13012
rect 18568 12836 18571 12888
rect 18571 12836 18617 12888
rect 18617 12836 18620 12888
rect 19912 16602 19964 16654
rect 19464 16478 19467 16530
rect 19467 16478 19513 16530
rect 19513 16478 19516 16530
rect 19464 16354 19467 16406
rect 19467 16354 19513 16406
rect 19513 16354 19516 16406
rect 19464 16230 19467 16282
rect 19467 16230 19513 16282
rect 19513 16230 19516 16282
rect 19464 16106 19467 16158
rect 19467 16106 19513 16158
rect 19513 16106 19516 16158
rect 19464 15982 19467 16034
rect 19467 15982 19513 16034
rect 19513 15982 19516 16034
rect 19464 15858 19467 15910
rect 19467 15858 19513 15910
rect 19513 15858 19516 15910
rect 19464 15734 19467 15786
rect 19467 15734 19513 15786
rect 19513 15734 19516 15786
rect 19464 15610 19467 15662
rect 19467 15610 19513 15662
rect 19513 15610 19516 15662
rect 19464 15486 19467 15538
rect 19467 15486 19513 15538
rect 19513 15486 19516 15538
rect 19240 14944 19243 14996
rect 19243 14944 19289 14996
rect 19289 14944 19292 14996
rect 19240 14820 19243 14872
rect 19243 14820 19289 14872
rect 19289 14820 19292 14872
rect 19240 14696 19243 14748
rect 19243 14696 19289 14748
rect 19289 14696 19292 14748
rect 19240 14572 19243 14624
rect 19243 14572 19289 14624
rect 19289 14572 19292 14624
rect 19240 14448 19243 14500
rect 19243 14448 19289 14500
rect 19289 14448 19292 14500
rect 19240 14324 19243 14376
rect 19243 14324 19289 14376
rect 19289 14324 19292 14376
rect 19240 14200 19243 14252
rect 19243 14200 19289 14252
rect 19289 14200 19292 14252
rect 19240 14076 19243 14128
rect 19243 14076 19289 14128
rect 19289 14076 19292 14128
rect 19240 13952 19243 14004
rect 19243 13952 19289 14004
rect 19289 13952 19292 14004
rect 19240 13828 19243 13880
rect 19243 13828 19289 13880
rect 19289 13828 19292 13880
rect 19240 13704 19243 13756
rect 19243 13704 19289 13756
rect 19289 13704 19292 13756
rect 19240 13580 19243 13632
rect 19243 13580 19289 13632
rect 19289 13580 19292 13632
rect 19240 13456 19243 13508
rect 19243 13456 19289 13508
rect 19289 13456 19292 13508
rect 19240 13332 19243 13384
rect 19243 13332 19289 13384
rect 19289 13332 19292 13384
rect 19240 13208 19243 13260
rect 19243 13208 19289 13260
rect 19289 13208 19292 13260
rect 19240 13084 19243 13136
rect 19243 13084 19289 13136
rect 19289 13084 19292 13136
rect 19240 12960 19243 13012
rect 19243 12960 19289 13012
rect 19289 12960 19292 13012
rect 19240 12836 19243 12888
rect 19243 12836 19289 12888
rect 19289 12836 19292 12888
rect 17000 11757 17052 11758
rect 17000 11706 17003 11757
rect 17003 11706 17049 11757
rect 17049 11706 17052 11757
rect 17000 11582 17003 11634
rect 17003 11582 17049 11634
rect 17049 11582 17052 11634
rect 17000 11458 17003 11510
rect 17003 11458 17049 11510
rect 17049 11458 17052 11510
rect 17448 11757 17500 11758
rect 17448 11706 17451 11757
rect 17451 11706 17497 11757
rect 17497 11706 17500 11757
rect 17448 11582 17451 11634
rect 17451 11582 17497 11634
rect 17497 11582 17500 11634
rect 17448 11458 17451 11510
rect 17451 11458 17497 11510
rect 17497 11458 17500 11510
rect 18808 11859 18860 11911
rect 19912 16478 19915 16530
rect 19915 16478 19961 16530
rect 19961 16478 19964 16530
rect 19912 16354 19915 16406
rect 19915 16354 19961 16406
rect 19961 16354 19964 16406
rect 19912 16230 19915 16282
rect 19915 16230 19961 16282
rect 19961 16230 19964 16282
rect 19912 16106 19915 16158
rect 19915 16106 19961 16158
rect 19961 16106 19964 16158
rect 19912 15982 19915 16034
rect 19915 15982 19961 16034
rect 19961 15982 19964 16034
rect 19912 15858 19915 15910
rect 19915 15858 19961 15910
rect 19961 15858 19964 15910
rect 19912 15734 19915 15786
rect 19915 15734 19961 15786
rect 19961 15734 19964 15786
rect 19912 15610 19915 15662
rect 19915 15610 19961 15662
rect 19961 15610 19964 15662
rect 19912 15486 19915 15538
rect 19915 15486 19961 15538
rect 19961 15486 19964 15538
rect 19688 14944 19691 14996
rect 19691 14944 19737 14996
rect 19737 14944 19740 14996
rect 19688 14820 19691 14872
rect 19691 14820 19737 14872
rect 19737 14820 19740 14872
rect 19688 14696 19691 14748
rect 19691 14696 19737 14748
rect 19737 14696 19740 14748
rect 19688 14572 19691 14624
rect 19691 14572 19737 14624
rect 19737 14572 19740 14624
rect 19688 14448 19691 14500
rect 19691 14448 19737 14500
rect 19737 14448 19740 14500
rect 19688 14324 19691 14376
rect 19691 14324 19737 14376
rect 19737 14324 19740 14376
rect 19688 14200 19691 14252
rect 19691 14200 19737 14252
rect 19737 14200 19740 14252
rect 19688 14076 19691 14128
rect 19691 14076 19737 14128
rect 19737 14076 19740 14128
rect 19688 13952 19691 14004
rect 19691 13952 19737 14004
rect 19737 13952 19740 14004
rect 19688 13828 19691 13880
rect 19691 13828 19737 13880
rect 19737 13828 19740 13880
rect 19688 13704 19691 13756
rect 19691 13704 19737 13756
rect 19737 13704 19740 13756
rect 19688 13580 19691 13632
rect 19691 13580 19737 13632
rect 19737 13580 19740 13632
rect 19688 13456 19691 13508
rect 19691 13456 19737 13508
rect 19737 13456 19740 13508
rect 19688 13332 19691 13384
rect 19691 13332 19737 13384
rect 19737 13332 19740 13384
rect 19688 13208 19691 13260
rect 19691 13208 19737 13260
rect 19737 13208 19740 13260
rect 19688 13084 19691 13136
rect 19691 13084 19737 13136
rect 19737 13084 19740 13136
rect 19688 12960 19691 13012
rect 19691 12960 19737 13012
rect 19737 12960 19740 13012
rect 19688 12836 19691 12888
rect 19691 12836 19737 12888
rect 19737 12836 19740 12888
rect 18120 11757 18172 11758
rect 18120 11706 18123 11757
rect 18123 11706 18169 11757
rect 18169 11706 18172 11757
rect 18120 11582 18123 11634
rect 18123 11582 18169 11634
rect 18169 11582 18172 11634
rect 18120 11458 18123 11510
rect 18123 11458 18169 11510
rect 18169 11458 18172 11510
rect 18568 11757 18620 11758
rect 18568 11706 18571 11757
rect 18571 11706 18617 11757
rect 18617 11706 18620 11757
rect 18568 11582 18571 11634
rect 18571 11582 18617 11634
rect 18617 11582 18620 11634
rect 18568 11458 18571 11510
rect 18571 11458 18617 11510
rect 18617 11458 18620 11510
rect 19240 11757 19292 11758
rect 19240 11706 19243 11757
rect 19243 11706 19289 11757
rect 19289 11706 19292 11757
rect 19240 11582 19243 11634
rect 19243 11582 19289 11634
rect 19289 11582 19292 11634
rect 19240 11458 19243 11510
rect 19243 11458 19289 11510
rect 19289 11458 19292 11510
rect 19688 11757 19740 11758
rect 19688 11706 19691 11757
rect 19691 11706 19737 11757
rect 19737 11706 19740 11757
rect 19688 11582 19691 11634
rect 19691 11582 19737 11634
rect 19737 11582 19740 11634
rect 19688 11458 19691 11510
rect 19691 11458 19737 11510
rect 19737 11458 19740 11510
rect 2404 9312 2456 9364
rect 2611 9312 2663 9364
rect 3131 9312 3183 9364
rect 4095 9312 4147 9364
rect 4302 9312 4354 9364
rect 4822 9312 4874 9364
rect 5786 9312 5838 9364
rect 5993 9312 6045 9364
rect 6513 9312 6565 9364
rect 7671 9297 7716 9324
rect 7716 9297 7723 9324
rect 7671 9272 7723 9297
rect 8119 9272 8171 9324
rect 8567 9297 8574 9324
rect 8574 9297 8619 9324
rect 9304 9297 9349 9324
rect 9349 9297 9356 9324
rect 8567 9272 8619 9297
rect 9304 9272 9356 9297
rect 9752 9272 9804 9324
rect 10200 9297 10207 9324
rect 10207 9297 10252 9324
rect 10938 9297 10983 9324
rect 10983 9297 10990 9324
rect 10200 9272 10252 9297
rect 10938 9272 10990 9297
rect 11386 9272 11438 9324
rect 11834 9297 11841 9324
rect 11841 9297 11886 9324
rect 12572 9297 12617 9324
rect 12617 9297 12624 9324
rect 11834 9272 11886 9297
rect 12572 9272 12624 9297
rect 13020 9272 13072 9324
rect 13468 9297 13475 9324
rect 13475 9297 13520 9324
rect 13468 9272 13520 9297
rect 2404 9094 2456 9146
rect 2611 9106 2621 9146
rect 2621 9106 2663 9146
rect 2611 9094 2663 9106
rect 2404 8876 2456 8928
rect 2611 8898 2621 8928
rect 2621 8898 2663 8928
rect 2611 8876 2663 8898
rect 2404 8658 2456 8710
rect 2611 8690 2621 8710
rect 2621 8690 2663 8710
rect 2611 8658 2663 8690
rect 3131 9106 3135 9146
rect 3135 9106 3181 9146
rect 3181 9106 3183 9146
rect 3131 9094 3183 9106
rect 3131 8898 3135 8928
rect 3135 8898 3181 8928
rect 3181 8898 3183 8928
rect 3131 8876 3183 8898
rect 3131 8690 3135 8710
rect 3135 8690 3181 8710
rect 3181 8690 3183 8710
rect 3131 8658 3183 8690
rect 4095 9094 4147 9146
rect 4302 9106 4312 9146
rect 4312 9106 4354 9146
rect 4302 9094 4354 9106
rect 4095 8876 4147 8928
rect 4302 8898 4312 8928
rect 4312 8898 4354 8928
rect 4302 8876 4354 8898
rect 4095 8658 4147 8710
rect 4302 8690 4312 8710
rect 4312 8690 4354 8710
rect 4302 8658 4354 8690
rect 2404 8090 2456 8142
rect 2616 8139 2668 8142
rect 2616 8093 2642 8139
rect 2642 8093 2668 8139
rect 2616 8090 2668 8093
rect 2624 7827 2667 7879
rect 2667 7827 2676 7879
rect 2624 7610 2667 7662
rect 2667 7610 2676 7662
rect 2624 7392 2667 7444
rect 2667 7392 2676 7444
rect 2624 7174 2667 7226
rect 2667 7174 2676 7226
rect 2624 6956 2667 7008
rect 2667 6956 2676 7008
rect 2624 6739 2667 6791
rect 2667 6739 2676 6791
rect 4822 9106 4826 9146
rect 4826 9106 4872 9146
rect 4872 9106 4874 9146
rect 4822 9094 4874 9106
rect 4822 8898 4826 8928
rect 4826 8898 4872 8928
rect 4872 8898 4874 8928
rect 4822 8876 4874 8898
rect 4822 8690 4826 8710
rect 4826 8690 4872 8710
rect 4872 8690 4874 8710
rect 4822 8658 4874 8690
rect 5786 9094 5838 9146
rect 5993 9106 6003 9146
rect 6003 9106 6045 9146
rect 5993 9094 6045 9106
rect 5786 8876 5838 8928
rect 5993 8898 6003 8928
rect 6003 8898 6045 8928
rect 5993 8876 6045 8898
rect 5786 8658 5838 8710
rect 5993 8690 6003 8710
rect 6003 8690 6045 8710
rect 5993 8658 6045 8690
rect 4095 8090 4147 8142
rect 4307 8139 4359 8142
rect 4307 8093 4333 8139
rect 4333 8093 4359 8139
rect 4307 8090 4359 8093
rect 3138 7827 3181 7879
rect 3181 7827 3190 7879
rect 3138 7610 3181 7662
rect 3181 7610 3190 7662
rect 3138 7392 3181 7444
rect 3181 7392 3190 7444
rect 3138 7174 3181 7226
rect 3181 7174 3190 7226
rect 3138 6956 3181 7008
rect 3181 6956 3190 7008
rect 3138 6739 3181 6791
rect 3181 6739 3190 6791
rect 2841 5522 2845 5574
rect 2845 5522 2891 5574
rect 2891 5522 2893 5574
rect 2841 5304 2845 5356
rect 2845 5304 2891 5356
rect 2891 5304 2893 5356
rect 4315 7827 4358 7879
rect 4358 7827 4367 7879
rect 4315 7610 4358 7662
rect 4358 7610 4367 7662
rect 4315 7392 4358 7444
rect 4358 7392 4367 7444
rect 4315 7174 4358 7226
rect 4358 7174 4367 7226
rect 4315 6956 4358 7008
rect 4358 6956 4367 7008
rect 4315 6739 4358 6791
rect 4358 6739 4367 6791
rect 3355 5522 3359 5574
rect 3359 5522 3405 5574
rect 3405 5522 3407 5574
rect 3355 5304 3359 5356
rect 3359 5304 3405 5356
rect 3405 5304 3407 5356
rect 6513 9106 6517 9146
rect 6517 9106 6563 9146
rect 6563 9106 6565 9146
rect 6513 9094 6565 9106
rect 6513 8898 6517 8928
rect 6517 8898 6563 8928
rect 6563 8898 6565 8928
rect 6513 8876 6565 8898
rect 6513 8690 6517 8710
rect 6517 8690 6563 8710
rect 6563 8690 6565 8710
rect 6513 8658 6565 8690
rect 7671 9054 7723 9106
rect 8119 9054 8171 9106
rect 7671 8880 7723 8888
rect 7671 8836 7674 8880
rect 7674 8836 7720 8880
rect 7720 8836 7723 8880
rect 7671 8626 7723 8670
rect 7671 8618 7674 8626
rect 7674 8618 7720 8626
rect 7720 8618 7723 8626
rect 7897 8962 7898 8973
rect 7898 8962 7944 8973
rect 7944 8962 7949 8973
rect 7897 8921 7949 8962
rect 7897 8753 7949 8755
rect 7897 8707 7898 8753
rect 7898 8707 7944 8753
rect 7944 8707 7949 8753
rect 7897 8703 7949 8707
rect 8567 9054 8619 9106
rect 8119 8880 8171 8888
rect 8119 8836 8122 8880
rect 8122 8836 8168 8880
rect 8168 8836 8171 8880
rect 8119 8626 8171 8670
rect 8119 8618 8122 8626
rect 8122 8618 8168 8626
rect 8168 8618 8171 8626
rect 8341 8962 8346 8973
rect 8346 8962 8392 8973
rect 8392 8962 8393 8973
rect 8341 8921 8393 8962
rect 8341 8753 8393 8755
rect 8341 8707 8346 8753
rect 8346 8707 8392 8753
rect 8392 8707 8393 8753
rect 8341 8703 8393 8707
rect 7897 8485 7949 8537
rect 9304 9054 9356 9106
rect 8567 8880 8619 8888
rect 8567 8836 8570 8880
rect 8570 8836 8616 8880
rect 8616 8836 8619 8880
rect 8567 8626 8619 8670
rect 8567 8618 8570 8626
rect 8570 8618 8616 8626
rect 8616 8618 8619 8626
rect 9752 9054 9804 9106
rect 9304 8880 9356 8888
rect 9304 8836 9307 8880
rect 9307 8836 9353 8880
rect 9353 8836 9356 8880
rect 8341 8485 8393 8537
rect 5786 8090 5838 8142
rect 5998 8139 6050 8142
rect 5998 8093 6024 8139
rect 6024 8093 6050 8139
rect 5998 8090 6050 8093
rect 4829 7827 4872 7879
rect 4872 7827 4881 7879
rect 4829 7610 4872 7662
rect 4872 7610 4881 7662
rect 4829 7392 4872 7444
rect 4872 7392 4881 7444
rect 4829 7174 4872 7226
rect 4872 7174 4881 7226
rect 4829 6956 4872 7008
rect 4872 6956 4881 7008
rect 4829 6739 4872 6791
rect 4872 6739 4881 6791
rect 4532 5522 4536 5574
rect 4536 5522 4582 5574
rect 4582 5522 4584 5574
rect 4532 5304 4536 5356
rect 4536 5304 4582 5356
rect 4582 5304 4584 5356
rect 6006 7827 6049 7879
rect 6049 7827 6058 7879
rect 6006 7610 6049 7662
rect 6049 7610 6058 7662
rect 6006 7392 6049 7444
rect 6049 7392 6058 7444
rect 6006 7174 6049 7226
rect 6049 7174 6058 7226
rect 6006 6956 6049 7008
rect 6049 6956 6058 7008
rect 6006 6739 6049 6791
rect 6049 6739 6058 6791
rect 5046 5522 5050 5574
rect 5050 5522 5096 5574
rect 5096 5522 5098 5574
rect 5046 5304 5050 5356
rect 5050 5304 5096 5356
rect 5096 5304 5098 5356
rect 9304 8626 9356 8670
rect 9304 8618 9307 8626
rect 9307 8618 9353 8626
rect 9353 8618 9356 8626
rect 9530 8962 9531 8973
rect 9531 8962 9577 8973
rect 9577 8962 9582 8973
rect 9530 8921 9582 8962
rect 9530 8753 9582 8755
rect 9530 8707 9531 8753
rect 9531 8707 9577 8753
rect 9577 8707 9582 8753
rect 9530 8703 9582 8707
rect 10200 9054 10252 9106
rect 9752 8880 9804 8888
rect 9752 8836 9755 8880
rect 9755 8836 9801 8880
rect 9801 8836 9804 8880
rect 9752 8626 9804 8670
rect 9752 8618 9755 8626
rect 9755 8618 9801 8626
rect 9801 8618 9804 8626
rect 9974 8962 9979 8973
rect 9979 8962 10025 8973
rect 10025 8962 10026 8973
rect 9974 8921 10026 8962
rect 9974 8753 10026 8755
rect 9974 8707 9979 8753
rect 9979 8707 10025 8753
rect 10025 8707 10026 8753
rect 9974 8703 10026 8707
rect 9530 8485 9582 8537
rect 10938 9054 10990 9106
rect 10200 8880 10252 8888
rect 10200 8836 10203 8880
rect 10203 8836 10249 8880
rect 10249 8836 10252 8880
rect 10200 8626 10252 8670
rect 10200 8618 10203 8626
rect 10203 8618 10249 8626
rect 10249 8618 10252 8626
rect 11386 9054 11438 9106
rect 10938 8880 10990 8888
rect 10938 8836 10941 8880
rect 10941 8836 10987 8880
rect 10987 8836 10990 8880
rect 9974 8485 10026 8537
rect 10938 8626 10990 8670
rect 10938 8618 10941 8626
rect 10941 8618 10987 8626
rect 10987 8618 10990 8626
rect 11164 8962 11165 8973
rect 11165 8962 11211 8973
rect 11211 8962 11216 8973
rect 11164 8921 11216 8962
rect 11164 8753 11216 8755
rect 11164 8707 11165 8753
rect 11165 8707 11211 8753
rect 11211 8707 11216 8753
rect 11164 8703 11216 8707
rect 11834 9054 11886 9106
rect 11386 8880 11438 8888
rect 11386 8836 11389 8880
rect 11389 8836 11435 8880
rect 11435 8836 11438 8880
rect 11386 8626 11438 8670
rect 11386 8618 11389 8626
rect 11389 8618 11435 8626
rect 11435 8618 11438 8626
rect 11608 8962 11613 8973
rect 11613 8962 11659 8973
rect 11659 8962 11660 8973
rect 11608 8921 11660 8962
rect 11608 8753 11660 8755
rect 11608 8707 11613 8753
rect 11613 8707 11659 8753
rect 11659 8707 11660 8753
rect 11608 8703 11660 8707
rect 11164 8485 11216 8537
rect 12572 9054 12624 9106
rect 11834 8880 11886 8888
rect 11834 8836 11837 8880
rect 11837 8836 11883 8880
rect 11883 8836 11886 8880
rect 11834 8626 11886 8670
rect 11834 8618 11837 8626
rect 11837 8618 11883 8626
rect 11883 8618 11886 8626
rect 13020 9054 13072 9106
rect 12572 8880 12624 8888
rect 12572 8836 12575 8880
rect 12575 8836 12621 8880
rect 12621 8836 12624 8880
rect 11608 8485 11660 8537
rect 12572 8626 12624 8670
rect 12572 8618 12575 8626
rect 12575 8618 12621 8626
rect 12621 8618 12624 8626
rect 12798 8962 12799 8973
rect 12799 8962 12845 8973
rect 12845 8962 12850 8973
rect 12798 8921 12850 8962
rect 12798 8753 12850 8755
rect 12798 8707 12799 8753
rect 12799 8707 12845 8753
rect 12845 8707 12850 8753
rect 12798 8703 12850 8707
rect 13468 9054 13520 9106
rect 13020 8880 13072 8888
rect 13020 8836 13023 8880
rect 13023 8836 13069 8880
rect 13069 8836 13072 8880
rect 13020 8626 13072 8670
rect 13020 8618 13023 8626
rect 13023 8618 13069 8626
rect 13069 8618 13072 8626
rect 13242 8962 13247 8973
rect 13247 8962 13293 8973
rect 13293 8962 13294 8973
rect 13242 8921 13294 8962
rect 13242 8753 13294 8755
rect 13242 8707 13247 8753
rect 13247 8707 13293 8753
rect 13293 8707 13294 8753
rect 13242 8703 13294 8707
rect 12798 8485 12850 8537
rect 13468 8880 13520 8888
rect 13468 8836 13471 8880
rect 13471 8836 13517 8880
rect 13517 8836 13520 8880
rect 13468 8626 13520 8670
rect 13468 8618 13471 8626
rect 13471 8618 13517 8626
rect 13517 8618 13520 8626
rect 13242 8485 13294 8537
rect 6520 7827 6563 7879
rect 6563 7827 6572 7879
rect 6520 7610 6563 7662
rect 6563 7610 6572 7662
rect 6520 7392 6563 7444
rect 6563 7392 6572 7444
rect 6520 7174 6563 7226
rect 6563 7174 6572 7226
rect 6520 6956 6563 7008
rect 6563 6956 6572 7008
rect 6520 6739 6563 6791
rect 6563 6739 6572 6791
rect 6223 5522 6227 5574
rect 6227 5522 6273 5574
rect 6273 5522 6275 5574
rect 6223 5304 6227 5356
rect 6227 5304 6273 5356
rect 6273 5304 6275 5356
rect 7671 7793 7674 7819
rect 7674 7793 7720 7819
rect 7720 7793 7723 7819
rect 7671 7767 7723 7793
rect 7671 7577 7674 7601
rect 7674 7577 7720 7601
rect 7720 7577 7723 7601
rect 7671 7549 7723 7577
rect 7671 7361 7674 7383
rect 7674 7361 7720 7383
rect 7720 7361 7723 7383
rect 7671 7331 7723 7361
rect 8119 7793 8122 7819
rect 8122 7793 8168 7819
rect 8168 7793 8171 7819
rect 8119 7767 8171 7793
rect 8119 7577 8122 7601
rect 8122 7577 8168 7601
rect 8168 7577 8171 7601
rect 8119 7549 8171 7577
rect 8119 7361 8122 7383
rect 8122 7361 8168 7383
rect 8168 7361 8171 7383
rect 8119 7331 8171 7361
rect 8567 7793 8570 7819
rect 8570 7793 8616 7819
rect 8616 7793 8619 7819
rect 8567 7767 8619 7793
rect 8567 7577 8570 7601
rect 8570 7577 8616 7601
rect 8616 7577 8619 7601
rect 8567 7549 8619 7577
rect 8567 7361 8570 7383
rect 8570 7361 8616 7383
rect 8616 7361 8619 7383
rect 8567 7331 8619 7361
rect 9304 7793 9307 7819
rect 9307 7793 9353 7819
rect 9353 7793 9356 7819
rect 9304 7767 9356 7793
rect 9304 7577 9307 7601
rect 9307 7577 9353 7601
rect 9353 7577 9356 7601
rect 9304 7549 9356 7577
rect 9304 7361 9307 7383
rect 9307 7361 9353 7383
rect 9353 7361 9356 7383
rect 9304 7331 9356 7361
rect 9752 7793 9755 7819
rect 9755 7793 9801 7819
rect 9801 7793 9804 7819
rect 9752 7767 9804 7793
rect 9752 7577 9755 7601
rect 9755 7577 9801 7601
rect 9801 7577 9804 7601
rect 9752 7549 9804 7577
rect 9752 7361 9755 7383
rect 9755 7361 9801 7383
rect 9801 7361 9804 7383
rect 9752 7331 9804 7361
rect 10200 7793 10203 7819
rect 10203 7793 10249 7819
rect 10249 7793 10252 7819
rect 10200 7767 10252 7793
rect 10200 7577 10203 7601
rect 10203 7577 10249 7601
rect 10249 7577 10252 7601
rect 10200 7549 10252 7577
rect 10200 7361 10203 7383
rect 10203 7361 10249 7383
rect 10249 7361 10252 7383
rect 10200 7331 10252 7361
rect 10938 7793 10941 7819
rect 10941 7793 10987 7819
rect 10987 7793 10990 7819
rect 10938 7767 10990 7793
rect 10938 7577 10941 7601
rect 10941 7577 10987 7601
rect 10987 7577 10990 7601
rect 10938 7549 10990 7577
rect 10938 7361 10941 7383
rect 10941 7361 10987 7383
rect 10987 7361 10990 7383
rect 10938 7331 10990 7361
rect 11386 7793 11389 7819
rect 11389 7793 11435 7819
rect 11435 7793 11438 7819
rect 11386 7767 11438 7793
rect 11386 7577 11389 7601
rect 11389 7577 11435 7601
rect 11435 7577 11438 7601
rect 11386 7549 11438 7577
rect 11386 7361 11389 7383
rect 11389 7361 11435 7383
rect 11435 7361 11438 7383
rect 11386 7331 11438 7361
rect 11834 7793 11837 7819
rect 11837 7793 11883 7819
rect 11883 7793 11886 7819
rect 11834 7767 11886 7793
rect 11834 7577 11837 7601
rect 11837 7577 11883 7601
rect 11883 7577 11886 7601
rect 11834 7549 11886 7577
rect 11834 7361 11837 7383
rect 11837 7361 11883 7383
rect 11883 7361 11886 7383
rect 11834 7331 11886 7361
rect 12572 7793 12575 7819
rect 12575 7793 12621 7819
rect 12621 7793 12624 7819
rect 12572 7767 12624 7793
rect 12572 7577 12575 7601
rect 12575 7577 12621 7601
rect 12621 7577 12624 7601
rect 12572 7549 12624 7577
rect 12572 7361 12575 7383
rect 12575 7361 12621 7383
rect 12621 7361 12624 7383
rect 12572 7331 12624 7361
rect 13020 7793 13023 7819
rect 13023 7793 13069 7819
rect 13069 7793 13072 7819
rect 13020 7767 13072 7793
rect 13020 7577 13023 7601
rect 13023 7577 13069 7601
rect 13069 7577 13072 7601
rect 13020 7549 13072 7577
rect 13020 7361 13023 7383
rect 13023 7361 13069 7383
rect 13069 7361 13072 7383
rect 13020 7331 13072 7361
rect 13468 7793 13471 7819
rect 13471 7793 13517 7819
rect 13517 7793 13520 7819
rect 13468 7767 13520 7793
rect 13468 7577 13471 7601
rect 13471 7577 13517 7601
rect 13517 7577 13520 7601
rect 13468 7549 13520 7577
rect 13468 7361 13471 7383
rect 13471 7361 13517 7383
rect 13517 7361 13520 7383
rect 13468 7331 13520 7361
rect 7675 6657 7727 6709
rect 7675 6440 7727 6492
rect 8119 6658 8171 6710
rect 8119 6440 8171 6492
rect 7675 6254 7720 6274
rect 7720 6254 7727 6274
rect 7675 6222 7727 6254
rect 7675 6042 7720 6056
rect 7720 6042 7727 6056
rect 7675 6004 7727 6042
rect 7675 5830 7720 5839
rect 7720 5830 7727 5839
rect 7675 5787 7727 5830
rect 6737 5522 6741 5574
rect 6741 5522 6787 5574
rect 6787 5522 6789 5574
rect 6737 5304 6741 5356
rect 6741 5304 6787 5356
rect 6787 5304 6789 5356
rect 7447 5558 7499 5604
rect 7447 5552 7450 5558
rect 7450 5552 7496 5558
rect 7496 5552 7499 5558
rect 7447 5344 7499 5386
rect 7447 5334 7450 5344
rect 7450 5334 7496 5344
rect 7496 5334 7499 5344
rect 8563 6657 8615 6709
rect 8563 6440 8615 6492
rect 8119 6254 8122 6275
rect 8122 6254 8168 6275
rect 8168 6254 8171 6275
rect 8119 6223 8171 6254
rect 8119 6042 8122 6057
rect 8122 6042 8168 6057
rect 8168 6042 8171 6057
rect 8119 6005 8171 6042
rect 8119 5830 8122 5839
rect 8122 5830 8168 5839
rect 8168 5830 8171 5839
rect 8119 5787 8171 5830
rect 7895 5558 7947 5604
rect 7895 5552 7898 5558
rect 7898 5552 7944 5558
rect 7944 5552 7947 5558
rect 7895 5344 7947 5386
rect 7895 5334 7898 5344
rect 7898 5334 7944 5344
rect 7944 5334 7947 5344
rect 8563 6254 8570 6274
rect 8570 6254 8615 6274
rect 8563 6222 8615 6254
rect 8563 6042 8570 6056
rect 8570 6042 8615 6056
rect 8563 6004 8615 6042
rect 8563 5830 8570 5839
rect 8570 5830 8615 5839
rect 8563 5787 8615 5830
rect 8119 5618 8122 5622
rect 8122 5618 8168 5622
rect 8168 5618 8171 5622
rect 8119 5570 8171 5618
rect 8119 5352 8171 5404
rect 8343 5558 8395 5604
rect 8343 5552 8346 5558
rect 8346 5552 8392 5558
rect 8392 5552 8395 5558
rect 8343 5344 8395 5386
rect 8343 5334 8346 5344
rect 8346 5334 8392 5344
rect 8392 5334 8395 5344
rect 9308 6657 9360 6709
rect 9308 6440 9360 6492
rect 9752 6658 9804 6710
rect 9752 6440 9804 6492
rect 9308 6254 9353 6274
rect 9353 6254 9360 6274
rect 9308 6222 9360 6254
rect 9308 6042 9353 6056
rect 9353 6042 9360 6056
rect 9308 6004 9360 6042
rect 9308 5830 9353 5839
rect 9353 5830 9360 5839
rect 9308 5787 9360 5830
rect 8791 5558 8843 5604
rect 8791 5552 8794 5558
rect 8794 5552 8840 5558
rect 8840 5552 8843 5558
rect 8791 5344 8843 5386
rect 8791 5334 8794 5344
rect 8794 5334 8840 5344
rect 8840 5334 8843 5344
rect 9080 5558 9132 5604
rect 9080 5552 9083 5558
rect 9083 5552 9129 5558
rect 9129 5552 9132 5558
rect 9080 5344 9132 5386
rect 9080 5334 9083 5344
rect 9083 5334 9129 5344
rect 9129 5334 9132 5344
rect 10196 6657 10248 6709
rect 10196 6440 10248 6492
rect 9752 6254 9755 6275
rect 9755 6254 9801 6275
rect 9801 6254 9804 6275
rect 9752 6223 9804 6254
rect 9752 6042 9755 6057
rect 9755 6042 9801 6057
rect 9801 6042 9804 6057
rect 9752 6005 9804 6042
rect 9752 5830 9755 5839
rect 9755 5830 9801 5839
rect 9801 5830 9804 5839
rect 9752 5787 9804 5830
rect 9528 5558 9580 5604
rect 9528 5552 9531 5558
rect 9531 5552 9577 5558
rect 9577 5552 9580 5558
rect 9528 5344 9580 5386
rect 9528 5334 9531 5344
rect 9531 5334 9577 5344
rect 9577 5334 9580 5344
rect 10196 6254 10203 6274
rect 10203 6254 10248 6274
rect 10196 6222 10248 6254
rect 10196 6042 10203 6056
rect 10203 6042 10248 6056
rect 10196 6004 10248 6042
rect 10196 5830 10203 5839
rect 10203 5830 10248 5839
rect 10196 5787 10248 5830
rect 9752 5618 9755 5622
rect 9755 5618 9801 5622
rect 9801 5618 9804 5622
rect 9752 5570 9804 5618
rect 9752 5352 9804 5404
rect 9976 5558 10028 5604
rect 9976 5552 9979 5558
rect 9979 5552 10025 5558
rect 10025 5552 10028 5558
rect 9976 5344 10028 5386
rect 9976 5334 9979 5344
rect 9979 5334 10025 5344
rect 10025 5334 10028 5344
rect 10942 6657 10994 6709
rect 10942 6440 10994 6492
rect 11386 6658 11438 6710
rect 11386 6440 11438 6492
rect 10942 6254 10987 6274
rect 10987 6254 10994 6274
rect 10942 6222 10994 6254
rect 10942 6042 10987 6056
rect 10987 6042 10994 6056
rect 10942 6004 10994 6042
rect 10942 5830 10987 5839
rect 10987 5830 10994 5839
rect 10942 5787 10994 5830
rect 10424 5558 10476 5604
rect 10424 5552 10427 5558
rect 10427 5552 10473 5558
rect 10473 5552 10476 5558
rect 10424 5344 10476 5386
rect 10424 5334 10427 5344
rect 10427 5334 10473 5344
rect 10473 5334 10476 5344
rect 10714 5558 10766 5604
rect 10714 5552 10717 5558
rect 10717 5552 10763 5558
rect 10763 5552 10766 5558
rect 10714 5344 10766 5386
rect 10714 5334 10717 5344
rect 10717 5334 10763 5344
rect 10763 5334 10766 5344
rect 11830 6657 11882 6709
rect 11830 6440 11882 6492
rect 11386 6254 11389 6275
rect 11389 6254 11435 6275
rect 11435 6254 11438 6275
rect 11386 6223 11438 6254
rect 11386 6042 11389 6057
rect 11389 6042 11435 6057
rect 11435 6042 11438 6057
rect 11386 6005 11438 6042
rect 11386 5830 11389 5839
rect 11389 5830 11435 5839
rect 11435 5830 11438 5839
rect 11386 5787 11438 5830
rect 11162 5558 11214 5604
rect 11162 5552 11165 5558
rect 11165 5552 11211 5558
rect 11211 5552 11214 5558
rect 11162 5344 11214 5386
rect 11162 5334 11165 5344
rect 11165 5334 11211 5344
rect 11211 5334 11214 5344
rect 11830 6254 11837 6274
rect 11837 6254 11882 6274
rect 11830 6222 11882 6254
rect 11830 6042 11837 6056
rect 11837 6042 11882 6056
rect 11830 6004 11882 6042
rect 11830 5830 11837 5839
rect 11837 5830 11882 5839
rect 11830 5787 11882 5830
rect 11386 5618 11389 5622
rect 11389 5618 11435 5622
rect 11435 5618 11438 5622
rect 11386 5570 11438 5618
rect 11386 5352 11438 5404
rect 11610 5558 11662 5604
rect 11610 5552 11613 5558
rect 11613 5552 11659 5558
rect 11659 5552 11662 5558
rect 11610 5344 11662 5386
rect 11610 5334 11613 5344
rect 11613 5334 11659 5344
rect 11659 5334 11662 5344
rect 12576 6657 12628 6709
rect 12576 6440 12628 6492
rect 13020 6658 13072 6710
rect 13020 6440 13072 6492
rect 12576 6254 12621 6274
rect 12621 6254 12628 6274
rect 12576 6222 12628 6254
rect 12576 6042 12621 6056
rect 12621 6042 12628 6056
rect 12576 6004 12628 6042
rect 12576 5830 12621 5839
rect 12621 5830 12628 5839
rect 12576 5787 12628 5830
rect 12058 5558 12110 5604
rect 12058 5552 12061 5558
rect 12061 5552 12107 5558
rect 12107 5552 12110 5558
rect 12058 5344 12110 5386
rect 12058 5334 12061 5344
rect 12061 5334 12107 5344
rect 12107 5334 12110 5344
rect 12348 5558 12400 5604
rect 12348 5552 12351 5558
rect 12351 5552 12397 5558
rect 12397 5552 12400 5558
rect 12348 5344 12400 5386
rect 12348 5334 12351 5344
rect 12351 5334 12397 5344
rect 12397 5334 12400 5344
rect 13464 6657 13516 6709
rect 13464 6440 13516 6492
rect 13020 6254 13023 6275
rect 13023 6254 13069 6275
rect 13069 6254 13072 6275
rect 13020 6223 13072 6254
rect 13020 6042 13023 6057
rect 13023 6042 13069 6057
rect 13069 6042 13072 6057
rect 13020 6005 13072 6042
rect 13020 5830 13023 5839
rect 13023 5830 13069 5839
rect 13069 5830 13072 5839
rect 13020 5787 13072 5830
rect 12796 5558 12848 5604
rect 12796 5552 12799 5558
rect 12799 5552 12845 5558
rect 12845 5552 12848 5558
rect 12796 5344 12848 5386
rect 12796 5334 12799 5344
rect 12799 5334 12845 5344
rect 12845 5334 12848 5344
rect 13464 6254 13471 6274
rect 13471 6254 13516 6274
rect 13464 6222 13516 6254
rect 13464 6042 13471 6056
rect 13471 6042 13516 6056
rect 13464 6004 13516 6042
rect 13464 5830 13471 5839
rect 13471 5830 13516 5839
rect 13464 5787 13516 5830
rect 13020 5618 13023 5622
rect 13023 5618 13069 5622
rect 13069 5618 13072 5622
rect 13020 5570 13072 5618
rect 13020 5352 13072 5404
rect 13244 5558 13296 5604
rect 13244 5552 13247 5558
rect 13247 5552 13293 5558
rect 13293 5552 13296 5558
rect 13244 5344 13296 5386
rect 13244 5334 13247 5344
rect 13247 5334 13293 5344
rect 13293 5334 13296 5344
rect 13692 5558 13744 5604
rect 13692 5552 13695 5558
rect 13695 5552 13741 5558
rect 13741 5552 13744 5558
rect 13692 5344 13744 5386
rect 13692 5334 13695 5344
rect 13695 5334 13741 5344
rect 13741 5334 13744 5344
rect 4533 4887 4585 4939
rect 6223 4685 6275 4737
rect 3355 4483 3407 4535
rect 5046 4281 5098 4333
rect 6737 4080 6789 4132
rect 7447 3698 7499 3712
rect 7447 3660 7450 3698
rect 7450 3660 7496 3698
rect 7496 3660 7499 3698
rect 7447 3484 7450 3495
rect 7450 3484 7496 3495
rect 7496 3484 7499 3495
rect 7447 3443 7499 3484
rect 2404 3159 2456 3211
rect 2404 2941 2456 2993
rect 4095 3159 4147 3211
rect 4095 2941 4147 2993
rect 5786 3159 5838 3211
rect 5786 2941 5838 2993
rect 7447 3225 7499 3277
rect 7447 3027 7499 3059
rect 7447 3007 7450 3027
rect 7450 3007 7496 3027
rect 7496 3007 7499 3027
rect 7447 2813 7450 2842
rect 7450 2813 7496 2842
rect 7496 2813 7499 2842
rect 7447 2790 7499 2813
rect 1753 1065 1805 1117
rect 1753 847 1805 899
rect 8119 3530 8171 3584
rect 8119 3484 8122 3530
rect 8122 3484 8168 3530
rect 8168 3484 8171 3530
rect 8119 3363 8171 3484
rect 8119 3317 8122 3363
rect 8122 3317 8168 3363
rect 8168 3317 8171 3363
rect 8119 3195 8171 3317
rect 8119 3149 8122 3195
rect 8122 3149 8168 3195
rect 8168 3149 8171 3195
rect 8119 3027 8171 3149
rect 8119 2981 8122 3027
rect 8122 2981 8168 3027
rect 8168 2981 8171 3027
rect 8119 2859 8171 2981
rect 8119 2813 8122 2859
rect 8122 2813 8168 2859
rect 8168 2813 8171 2859
rect 8119 2692 8171 2813
rect 8119 2646 8122 2692
rect 8122 2646 8168 2692
rect 8168 2646 8171 2692
rect 8119 2596 8171 2646
rect 8791 3698 8843 3712
rect 8791 3660 8794 3698
rect 8794 3660 8840 3698
rect 8840 3660 8843 3698
rect 8791 3484 8794 3495
rect 8794 3484 8840 3495
rect 8840 3484 8843 3495
rect 8791 3443 8843 3484
rect 8791 3225 8843 3277
rect 8791 3027 8843 3059
rect 8791 3007 8794 3027
rect 8794 3007 8840 3027
rect 8840 3007 8843 3027
rect 8791 2813 8794 2842
rect 8794 2813 8840 2842
rect 8840 2813 8843 2842
rect 8791 2790 8843 2813
rect 9080 3698 9132 3712
rect 9080 3660 9083 3698
rect 9083 3660 9129 3698
rect 9129 3660 9132 3698
rect 9080 3484 9083 3495
rect 9083 3484 9129 3495
rect 9129 3484 9132 3495
rect 9080 3443 9132 3484
rect 9080 3225 9132 3277
rect 9080 3027 9132 3059
rect 9080 3007 9083 3027
rect 9083 3007 9129 3027
rect 9129 3007 9132 3027
rect 9080 2813 9083 2842
rect 9083 2813 9129 2842
rect 9129 2813 9132 2842
rect 9080 2790 9132 2813
rect 9753 3530 9805 3584
rect 9753 3484 9755 3530
rect 9755 3484 9801 3530
rect 9801 3484 9805 3530
rect 9753 3363 9805 3484
rect 9753 3317 9755 3363
rect 9755 3317 9801 3363
rect 9801 3317 9805 3363
rect 9753 3195 9805 3317
rect 9753 3149 9755 3195
rect 9755 3149 9801 3195
rect 9801 3149 9805 3195
rect 9753 3027 9805 3149
rect 9753 2981 9755 3027
rect 9755 2981 9801 3027
rect 9801 2981 9805 3027
rect 9753 2859 9805 2981
rect 9753 2813 9755 2859
rect 9755 2813 9801 2859
rect 9801 2813 9805 2859
rect 9753 2692 9805 2813
rect 9753 2646 9755 2692
rect 9755 2646 9801 2692
rect 9801 2646 9805 2692
rect 9753 2596 9805 2646
rect 10424 3698 10476 3712
rect 10424 3660 10427 3698
rect 10427 3660 10473 3698
rect 10473 3660 10476 3698
rect 10424 3484 10427 3495
rect 10427 3484 10473 3495
rect 10473 3484 10476 3495
rect 10424 3443 10476 3484
rect 10424 3225 10476 3277
rect 10424 3027 10476 3059
rect 10424 3007 10427 3027
rect 10427 3007 10473 3027
rect 10473 3007 10476 3027
rect 10424 2813 10427 2842
rect 10427 2813 10473 2842
rect 10473 2813 10476 2842
rect 10424 2790 10476 2813
rect 10714 3698 10766 3712
rect 10714 3660 10717 3698
rect 10717 3660 10763 3698
rect 10763 3660 10766 3698
rect 10714 3484 10717 3495
rect 10717 3484 10763 3495
rect 10763 3484 10766 3495
rect 10714 3443 10766 3484
rect 10714 3225 10766 3277
rect 10714 3027 10766 3059
rect 10714 3007 10717 3027
rect 10717 3007 10763 3027
rect 10763 3007 10766 3027
rect 10714 2813 10717 2842
rect 10717 2813 10763 2842
rect 10763 2813 10766 2842
rect 10714 2790 10766 2813
rect 11386 3530 11438 3584
rect 11386 3484 11389 3530
rect 11389 3484 11435 3530
rect 11435 3484 11438 3530
rect 11386 3363 11438 3484
rect 11386 3317 11389 3363
rect 11389 3317 11435 3363
rect 11435 3317 11438 3363
rect 11386 3195 11438 3317
rect 11386 3149 11389 3195
rect 11389 3149 11435 3195
rect 11435 3149 11438 3195
rect 11386 3027 11438 3149
rect 11386 2981 11389 3027
rect 11389 2981 11435 3027
rect 11435 2981 11438 3027
rect 11386 2859 11438 2981
rect 11386 2813 11389 2859
rect 11389 2813 11435 2859
rect 11435 2813 11438 2859
rect 11386 2692 11438 2813
rect 11386 2646 11389 2692
rect 11389 2646 11435 2692
rect 11435 2646 11438 2692
rect 11386 2596 11438 2646
rect 12058 3698 12110 3712
rect 12058 3660 12061 3698
rect 12061 3660 12107 3698
rect 12107 3660 12110 3698
rect 12058 3484 12061 3495
rect 12061 3484 12107 3495
rect 12107 3484 12110 3495
rect 12058 3443 12110 3484
rect 12058 3225 12110 3277
rect 12058 3027 12110 3059
rect 12058 3007 12061 3027
rect 12061 3007 12107 3027
rect 12107 3007 12110 3027
rect 12058 2813 12061 2842
rect 12061 2813 12107 2842
rect 12107 2813 12110 2842
rect 12058 2790 12110 2813
rect 12348 3698 12400 3712
rect 12348 3660 12351 3698
rect 12351 3660 12397 3698
rect 12397 3660 12400 3698
rect 12348 3484 12351 3495
rect 12351 3484 12397 3495
rect 12397 3484 12400 3495
rect 12348 3443 12400 3484
rect 12348 3225 12400 3277
rect 12348 3027 12400 3059
rect 12348 3007 12351 3027
rect 12351 3007 12397 3027
rect 12397 3007 12400 3027
rect 12348 2813 12351 2842
rect 12351 2813 12397 2842
rect 12397 2813 12400 2842
rect 12348 2790 12400 2813
rect 13020 3530 13072 3584
rect 13020 3484 13023 3530
rect 13023 3484 13069 3530
rect 13069 3484 13072 3530
rect 13020 3363 13072 3484
rect 13020 3317 13023 3363
rect 13023 3317 13069 3363
rect 13069 3317 13072 3363
rect 13020 3195 13072 3317
rect 13020 3149 13023 3195
rect 13023 3149 13069 3195
rect 13069 3149 13072 3195
rect 13020 3027 13072 3149
rect 13020 2981 13023 3027
rect 13023 2981 13069 3027
rect 13069 2981 13072 3027
rect 13020 2859 13072 2981
rect 13020 2813 13023 2859
rect 13023 2813 13069 2859
rect 13069 2813 13072 2859
rect 13020 2692 13072 2813
rect 13020 2646 13023 2692
rect 13023 2646 13069 2692
rect 13069 2646 13072 2692
rect 13020 2596 13072 2646
rect 13692 3698 13744 3712
rect 13692 3660 13695 3698
rect 13695 3660 13741 3698
rect 13741 3660 13744 3698
rect 13692 3484 13695 3495
rect 13695 3484 13741 3495
rect 13741 3484 13744 3495
rect 13692 3443 13744 3484
rect 13692 3225 13744 3277
rect 13692 3027 13744 3059
rect 13692 3007 13695 3027
rect 13695 3007 13741 3027
rect 13741 3007 13744 3027
rect 13692 2813 13695 2842
rect 13695 2813 13741 2842
rect 13741 2813 13744 2842
rect 13692 2790 13744 2813
rect 7838 1824 7890 1876
rect 9001 1874 9053 1926
rect 7838 1606 7884 1658
rect 7884 1606 7890 1658
rect 9001 1656 9009 1708
rect 9009 1656 9053 1708
rect 9900 1956 9952 2008
rect 10111 1956 10163 2008
rect 10321 1956 10373 2008
rect 10532 1956 10584 2008
rect 10743 1956 10795 2008
rect 10954 1956 11006 2008
rect 11165 1956 11217 2008
rect 11375 1956 11427 2008
rect 11586 1956 11638 2008
rect 11798 1956 11850 2008
rect 12009 1956 12061 2008
rect 12219 1956 12271 2008
rect 12430 1956 12482 2008
rect 12641 1956 12693 2008
rect 12852 1956 12904 2008
rect 13063 1956 13115 2008
rect 13273 1956 13325 2008
rect 13484 1956 13536 2008
rect 9900 1738 9952 1790
rect 10111 1784 10163 1790
rect 10321 1784 10373 1790
rect 10111 1738 10118 1784
rect 10118 1738 10163 1784
rect 10321 1738 10322 1784
rect 10322 1738 10373 1784
rect 10532 1738 10584 1790
rect 10743 1784 10795 1790
rect 10743 1738 10750 1784
rect 10750 1738 10795 1784
rect 10954 1738 11006 1790
rect 11165 1738 11217 1790
rect 11375 1784 11427 1790
rect 11586 1784 11638 1790
rect 11375 1738 11383 1784
rect 11383 1738 11427 1784
rect 11586 1738 11587 1784
rect 11587 1738 11638 1784
rect 11798 1738 11850 1790
rect 12009 1784 12061 1790
rect 12009 1738 12015 1784
rect 12015 1738 12061 1784
rect 12219 1738 12271 1790
rect 12430 1738 12482 1790
rect 12641 1784 12693 1790
rect 12641 1738 12648 1784
rect 12648 1738 12693 1784
rect 12852 1738 12904 1790
rect 13063 1738 13115 1790
rect 13273 1784 13325 1790
rect 13273 1738 13280 1784
rect 13280 1738 13325 1784
rect 13484 1738 13536 1790
rect 7218 1375 7270 1427
rect 8642 1432 8902 1451
rect 8642 1399 8754 1432
rect 8754 1399 8800 1432
rect 8800 1399 8902 1432
rect 9613 1448 9873 1451
rect 9613 1402 9642 1448
rect 9642 1402 9782 1448
rect 9782 1402 9873 1448
rect 9613 1399 9873 1402
rect 7218 1157 7270 1209
rect 7447 1108 7499 1160
rect 7447 890 7499 942
rect 8474 1126 8526 1178
rect 8474 908 8526 960
rect 9660 1123 9712 1173
rect 9660 1121 9703 1123
rect 9703 1121 9712 1123
rect 9871 1121 9923 1173
rect 10082 1121 10134 1173
rect 10293 1121 10345 1173
rect 10504 1121 10556 1173
rect 10714 1121 10766 1173
rect 10925 1121 10977 1173
rect 11136 1121 11188 1173
rect 11347 1121 11399 1173
rect 11558 1121 11610 1173
rect 11769 1121 11821 1173
rect 11980 1121 12032 1173
rect 12191 1121 12243 1173
rect 12402 1121 12454 1173
rect 12612 1121 12664 1173
rect 12823 1121 12875 1173
rect 13034 1121 13086 1173
rect 13245 1121 13297 1173
rect 13456 1121 13508 1173
rect 9660 919 9712 955
rect 9660 903 9703 919
rect 9703 903 9712 919
rect 9871 903 9923 955
rect 10082 943 10134 955
rect 10082 903 10089 943
rect 10089 903 10134 943
rect 10293 903 10345 955
rect 10504 903 10556 955
rect 10714 943 10766 955
rect 10714 903 10721 943
rect 10721 903 10766 943
rect 10925 903 10977 955
rect 11136 903 11188 955
rect 11347 943 11399 955
rect 11347 903 11354 943
rect 11354 903 11399 943
rect 11558 903 11610 955
rect 11769 903 11821 955
rect 11980 943 12032 955
rect 11980 903 11986 943
rect 11986 903 12032 943
rect 12191 903 12243 955
rect 12402 903 12454 955
rect 12612 943 12664 955
rect 12612 903 12619 943
rect 12619 903 12664 943
rect 12823 903 12875 955
rect 13034 903 13086 955
rect 13245 943 13297 955
rect 13245 903 13251 943
rect 13251 903 13297 943
rect 13456 903 13508 955
rect 28045 1078 28097 1130
rect 28045 860 28097 912
rect 28045 642 28097 694
rect 28287 1078 28339 1130
rect 28287 860 28339 912
rect 28287 642 28339 694
rect 28529 1078 28581 1130
rect 28529 860 28581 912
rect 28529 642 28581 694
rect 28770 1078 28822 1130
rect 28770 860 28822 912
rect 29561 1065 29613 1117
rect 29561 847 29613 899
rect 28770 642 28822 694
rect 8918 237 8970 289
rect 9130 237 9182 289
rect 733 185 785 237
rect 945 185 997 237
rect 29059 185 29111 237
rect 29271 185 29323 237
rect 8918 19 8970 71
rect 9130 19 9182 71
rect 733 -33 785 19
rect 945 -33 997 19
rect 29059 -33 29111 19
rect 29271 -33 29323 19
<< metal2 >>
rect 645 30026 1525 30125
rect 645 29970 740 30026
rect 796 29970 951 30026
rect 1007 29970 1163 30026
rect 1219 29970 1374 30026
rect 1430 29970 1525 30026
rect 645 29808 1525 29970
rect 645 29752 740 29808
rect 796 29752 951 29808
rect 1007 29752 1163 29808
rect 1219 29752 1374 29808
rect 1430 29752 1525 29808
rect 645 29590 1525 29752
rect 645 29534 740 29590
rect 796 29534 951 29590
rect 1007 29534 1163 29590
rect 1219 29534 1374 29590
rect 1430 29534 1525 29590
rect 645 29372 1525 29534
rect 645 29316 740 29372
rect 796 29316 951 29372
rect 1007 29316 1163 29372
rect 1219 29316 1374 29372
rect 1430 29316 1525 29372
rect 407 28998 532 29037
rect 407 28942 442 28998
rect 498 28942 532 28998
rect 407 28780 532 28942
rect 407 28724 442 28780
rect 498 28724 532 28780
rect 407 28686 532 28724
rect 645 1382 1525 29316
rect 5436 30026 5790 30064
rect 5436 29970 5479 30026
rect 5535 29970 5691 30026
rect 5747 29970 5790 30026
rect 5436 29808 5790 29970
rect 5436 29752 5479 29808
rect 5535 29752 5691 29808
rect 5747 29752 5790 29808
rect 5436 29590 5790 29752
rect 5436 29534 5479 29590
rect 5535 29534 5691 29590
rect 5747 29534 5790 29590
rect 5436 29372 5790 29534
rect 5436 29316 5479 29372
rect 5535 29316 5691 29372
rect 5747 29316 5790 29372
rect 1618 28502 1746 28539
rect 1618 28446 1654 28502
rect 1710 28446 1746 28502
rect 1618 28284 1746 28446
rect 1618 28228 1654 28284
rect 1710 28228 1746 28284
rect 1618 28066 1746 28228
rect 1618 28010 1654 28066
rect 1710 28010 1746 28066
rect 1618 27848 1746 28010
rect 1618 27792 1654 27848
rect 1710 27792 1746 27848
rect 1618 27754 1746 27792
rect 2058 28502 2186 28539
rect 2058 28446 2094 28502
rect 2150 28446 2186 28502
rect 2058 28284 2186 28446
rect 2058 28228 2094 28284
rect 2150 28228 2186 28284
rect 2058 28066 2186 28228
rect 2058 28010 2094 28066
rect 2150 28010 2186 28066
rect 2058 27848 2186 28010
rect 2058 27792 2094 27848
rect 2150 27792 2186 27848
rect 2058 27754 2186 27792
rect 2290 28500 2511 28772
rect 2290 28448 2328 28500
rect 2380 28448 2511 28500
rect 2290 28282 2511 28448
rect 2290 28230 2328 28282
rect 2380 28230 2511 28282
rect 2290 28064 2511 28230
rect 2290 28012 2328 28064
rect 2380 28012 2511 28064
rect 2290 27846 2511 28012
rect 2290 27794 2328 27846
rect 2380 27794 2511 27846
rect 2290 27754 2511 27794
rect 2645 28500 2866 28772
rect 2645 28448 2776 28500
rect 2828 28448 2866 28500
rect 2645 28282 2866 28448
rect 2645 28230 2776 28282
rect 2828 28230 2866 28282
rect 2645 28064 2866 28230
rect 2645 28012 2776 28064
rect 2828 28012 2866 28064
rect 2645 27846 2866 28012
rect 2645 27794 2776 27846
rect 2828 27794 2866 27846
rect 2645 27754 2866 27794
rect 2970 28502 3098 28539
rect 2970 28446 3006 28502
rect 3062 28446 3098 28502
rect 2970 28284 3098 28446
rect 2970 28228 3006 28284
rect 3062 28228 3098 28284
rect 2970 28066 3098 28228
rect 2970 28010 3006 28066
rect 3062 28010 3098 28066
rect 2970 27848 3098 28010
rect 2970 27792 3006 27848
rect 3062 27792 3098 27848
rect 2970 27754 3098 27792
rect 3410 28502 3538 28539
rect 3410 28446 3446 28502
rect 3502 28446 3538 28502
rect 3410 28284 3538 28446
rect 3410 28228 3446 28284
rect 3502 28228 3538 28284
rect 3410 28066 3538 28228
rect 3410 28010 3446 28066
rect 3502 28010 3538 28066
rect 3410 27848 3538 28010
rect 3410 27792 3446 27848
rect 3502 27792 3538 27848
rect 3410 27754 3538 27792
rect 3850 28502 3978 28539
rect 3850 28446 3886 28502
rect 3942 28446 3978 28502
rect 3850 28284 3978 28446
rect 3850 28228 3886 28284
rect 3942 28228 3978 28284
rect 3850 28066 3978 28228
rect 3850 28010 3886 28066
rect 3942 28010 3978 28066
rect 3850 27848 3978 28010
rect 3850 27792 3886 27848
rect 3942 27792 3978 27848
rect 3850 27754 3978 27792
rect 4082 28500 4303 28772
rect 4082 28448 4120 28500
rect 4172 28448 4303 28500
rect 4082 28282 4303 28448
rect 4082 28230 4120 28282
rect 4172 28230 4303 28282
rect 4082 28064 4303 28230
rect 4082 28012 4120 28064
rect 4172 28012 4303 28064
rect 4082 27846 4303 28012
rect 4082 27794 4120 27846
rect 4172 27794 4303 27846
rect 4082 27754 4303 27794
rect 4437 28500 4658 28772
rect 4437 28448 4568 28500
rect 4620 28448 4658 28500
rect 4437 28282 4658 28448
rect 4437 28230 4568 28282
rect 4620 28230 4658 28282
rect 4437 28064 4658 28230
rect 4437 28012 4568 28064
rect 4620 28012 4658 28064
rect 4437 27846 4658 28012
rect 4437 27794 4568 27846
rect 4620 27794 4658 27846
rect 4437 27754 4658 27794
rect 4762 28502 4890 28539
rect 4762 28446 4798 28502
rect 4854 28446 4890 28502
rect 4762 28284 4890 28446
rect 4762 28228 4798 28284
rect 4854 28228 4890 28284
rect 4762 28066 4890 28228
rect 4762 28010 4798 28066
rect 4854 28010 4890 28066
rect 4762 27848 4890 28010
rect 4762 27792 4798 27848
rect 4854 27792 4890 27848
rect 4762 27754 4890 27792
rect 5202 28502 5330 28539
rect 5202 28446 5238 28502
rect 5294 28446 5330 28502
rect 5202 28284 5330 28446
rect 5202 28228 5238 28284
rect 5294 28228 5330 28284
rect 5202 28066 5330 28228
rect 5202 28010 5238 28066
rect 5294 28010 5330 28066
rect 5202 27848 5330 28010
rect 5202 27792 5238 27848
rect 5294 27792 5330 27848
rect 5202 27754 5330 27792
rect 5436 27736 5790 29316
rect 16353 30026 16706 30125
rect 16353 29970 16395 30026
rect 16451 29970 16607 30026
rect 16663 29970 16706 30026
rect 16353 29808 16706 29970
rect 16353 29752 16395 29808
rect 16451 29752 16607 29808
rect 16663 29752 16706 29808
rect 16353 29590 16706 29752
rect 16353 29534 16395 29590
rect 16451 29534 16607 29590
rect 16663 29534 16706 29590
rect 16353 29372 16706 29534
rect 16353 29316 16395 29372
rect 16451 29316 16607 29372
rect 16663 29316 16706 29372
rect 6545 29037 6670 29038
rect 13923 29037 14048 29038
rect 6543 28999 6672 29037
rect 6543 28943 6580 28999
rect 6636 28943 6672 28999
rect 6543 28781 6672 28943
rect 6543 28725 6580 28781
rect 6636 28725 6672 28781
rect 13922 28999 14051 29037
rect 13922 28943 13958 28999
rect 14014 28943 14051 28999
rect 13922 28781 14051 28943
rect 16353 28860 16706 29316
rect 23301 30026 23654 30064
rect 23301 29970 23343 30026
rect 23399 29970 23555 30026
rect 23611 29970 23654 30026
rect 23301 29808 23654 29970
rect 23301 29752 23343 29808
rect 23399 29752 23555 29808
rect 23611 29752 23654 29808
rect 23301 29590 23654 29752
rect 23301 29534 23343 29590
rect 23399 29534 23555 29590
rect 23611 29534 23654 29590
rect 23301 29372 23654 29534
rect 23301 29316 23343 29372
rect 23399 29316 23555 29372
rect 23611 29316 23654 29372
rect 5885 28403 6013 28440
rect 5885 28347 5921 28403
rect 5977 28347 6013 28403
rect 5885 28185 6013 28347
rect 5885 28129 5921 28185
rect 5977 28129 6013 28185
rect 5885 27967 6013 28129
rect 5885 27911 5921 27967
rect 5977 27911 6013 27967
rect 5885 27873 6013 27911
rect 6324 28403 6452 28440
rect 6324 28347 6360 28403
rect 6416 28347 6452 28403
rect 6324 28185 6452 28347
rect 6324 28129 6360 28185
rect 6416 28129 6452 28185
rect 6324 27967 6452 28129
rect 6324 27911 6360 27967
rect 6416 27911 6452 27967
rect 6324 27873 6452 27911
rect 6543 28185 6672 28725
rect 8997 28502 9125 28539
rect 8997 28446 9033 28502
rect 9089 28446 9125 28502
rect 6543 28133 6582 28185
rect 6634 28133 6672 28185
rect 6543 27967 6672 28133
rect 6543 27915 6582 27967
rect 6634 27915 6672 27967
rect 6543 27874 6672 27915
rect 7708 28346 7836 28383
rect 7708 28290 7744 28346
rect 7800 28290 7836 28346
rect 7708 28128 7836 28290
rect 7708 28072 7744 28128
rect 7800 28072 7836 28128
rect 7708 27910 7836 28072
rect 7708 27854 7744 27910
rect 7800 27854 7836 27910
rect 7708 27816 7836 27854
rect 8997 28284 9125 28446
rect 8997 28228 9033 28284
rect 9089 28228 9125 28284
rect 8997 28066 9125 28228
rect 8997 28010 9033 28066
rect 9089 28010 9125 28066
rect 8997 27848 9125 28010
rect 8997 27792 9033 27848
rect 9089 27792 9125 27848
rect 8997 27754 9125 27792
rect 9437 28502 9565 28539
rect 9437 28446 9473 28502
rect 9529 28446 9565 28502
rect 9437 28284 9565 28446
rect 9437 28228 9473 28284
rect 9529 28228 9565 28284
rect 9437 28066 9565 28228
rect 9437 28010 9473 28066
rect 9529 28010 9565 28066
rect 9437 27848 9565 28010
rect 9437 27792 9473 27848
rect 9529 27792 9565 27848
rect 9437 27754 9565 27792
rect 9669 28500 9890 28772
rect 9669 28448 9707 28500
rect 9759 28448 9890 28500
rect 9669 28282 9890 28448
rect 9669 28230 9707 28282
rect 9759 28230 9890 28282
rect 9669 28064 9890 28230
rect 9669 28012 9707 28064
rect 9759 28012 9890 28064
rect 9669 27846 9890 28012
rect 9669 27794 9707 27846
rect 9759 27794 9890 27846
rect 9669 27754 9890 27794
rect 10024 28500 10245 28772
rect 10024 28448 10155 28500
rect 10207 28448 10245 28500
rect 10024 28282 10245 28448
rect 10024 28230 10155 28282
rect 10207 28230 10245 28282
rect 10024 28064 10245 28230
rect 10024 28012 10155 28064
rect 10207 28012 10245 28064
rect 10024 27846 10245 28012
rect 10024 27794 10155 27846
rect 10207 27794 10245 27846
rect 10024 27754 10245 27794
rect 10349 28502 10477 28539
rect 10349 28446 10385 28502
rect 10441 28446 10477 28502
rect 10349 28284 10477 28446
rect 10349 28228 10385 28284
rect 10441 28228 10477 28284
rect 10349 28066 10477 28228
rect 10349 28010 10385 28066
rect 10441 28010 10477 28066
rect 10349 27848 10477 28010
rect 10349 27792 10385 27848
rect 10441 27792 10477 27848
rect 10349 27754 10477 27792
rect 10789 28502 10917 28539
rect 10789 28446 10825 28502
rect 10881 28446 10917 28502
rect 10789 28284 10917 28446
rect 10789 28228 10825 28284
rect 10881 28228 10917 28284
rect 10789 28066 10917 28228
rect 10789 28010 10825 28066
rect 10881 28010 10917 28066
rect 10789 27848 10917 28010
rect 10789 27792 10825 27848
rect 10881 27792 10917 27848
rect 10789 27754 10917 27792
rect 11229 28502 11357 28539
rect 11229 28446 11265 28502
rect 11321 28446 11357 28502
rect 11229 28284 11357 28446
rect 11229 28228 11265 28284
rect 11321 28228 11357 28284
rect 11229 28066 11357 28228
rect 11229 28010 11265 28066
rect 11321 28010 11357 28066
rect 11229 27848 11357 28010
rect 11229 27792 11265 27848
rect 11321 27792 11357 27848
rect 11229 27754 11357 27792
rect 11461 28500 11682 28772
rect 11461 28448 11499 28500
rect 11551 28448 11682 28500
rect 11461 28282 11682 28448
rect 11461 28230 11499 28282
rect 11551 28230 11682 28282
rect 11461 28064 11682 28230
rect 11461 28012 11499 28064
rect 11551 28012 11682 28064
rect 11461 27846 11682 28012
rect 11461 27794 11499 27846
rect 11551 27794 11682 27846
rect 11461 27754 11682 27794
rect 11816 28500 12037 28772
rect 13922 28725 13958 28781
rect 14014 28725 14051 28781
rect 11816 28448 11947 28500
rect 11999 28448 12037 28500
rect 11816 28282 12037 28448
rect 11816 28230 11947 28282
rect 11999 28230 12037 28282
rect 11816 28064 12037 28230
rect 11816 28012 11947 28064
rect 11999 28012 12037 28064
rect 11816 27846 12037 28012
rect 11816 27794 11947 27846
rect 11999 27794 12037 27846
rect 11816 27754 12037 27794
rect 12141 28502 12269 28539
rect 12141 28446 12177 28502
rect 12233 28446 12269 28502
rect 12141 28284 12269 28446
rect 12141 28228 12177 28284
rect 12233 28228 12269 28284
rect 12141 28066 12269 28228
rect 12141 28010 12177 28066
rect 12233 28010 12269 28066
rect 12141 27848 12269 28010
rect 12141 27792 12177 27848
rect 12233 27792 12269 27848
rect 12141 27754 12269 27792
rect 12581 28502 12709 28539
rect 12581 28446 12617 28502
rect 12673 28446 12709 28502
rect 12581 28284 12709 28446
rect 12581 28228 12617 28284
rect 12673 28228 12709 28284
rect 12581 28066 12709 28228
rect 12581 28010 12617 28066
rect 12673 28010 12709 28066
rect 12581 27848 12709 28010
rect 13264 28403 13392 28440
rect 13264 28347 13300 28403
rect 13356 28347 13392 28403
rect 13264 28185 13392 28347
rect 13264 28129 13300 28185
rect 13356 28129 13392 28185
rect 13264 27967 13392 28129
rect 13264 27911 13300 27967
rect 13356 27911 13392 27967
rect 13264 27873 13392 27911
rect 13703 28403 13831 28440
rect 13703 28347 13739 28403
rect 13795 28347 13831 28403
rect 13703 28185 13831 28347
rect 13703 28129 13739 28185
rect 13795 28129 13831 28185
rect 13703 27967 13831 28129
rect 13703 27911 13739 27967
rect 13795 27911 13831 27967
rect 13703 27873 13831 27911
rect 13922 28185 14051 28725
rect 13922 28133 13961 28185
rect 14013 28133 14051 28185
rect 13922 27967 14051 28133
rect 13922 27915 13961 27967
rect 14013 27915 14051 27967
rect 13922 27874 14051 27915
rect 14225 28496 16706 28860
rect 12581 27792 12617 27848
rect 12673 27792 12709 27848
rect 12581 27754 12709 27792
rect 14225 27736 14578 28496
rect 16880 28394 17008 28431
rect 15087 28346 15215 28383
rect 15087 28290 15123 28346
rect 15179 28290 15215 28346
rect 15087 28128 15215 28290
rect 15087 28072 15123 28128
rect 15179 28072 15215 28128
rect 15087 27910 15215 28072
rect 15087 27854 15123 27910
rect 15179 27854 15215 27910
rect 15087 27816 15215 27854
rect 16880 28338 16916 28394
rect 16972 28338 17008 28394
rect 16880 28176 17008 28338
rect 17112 28305 17334 28998
rect 16880 28120 16916 28176
rect 16972 28120 17008 28176
rect 16880 27958 17008 28120
rect 16880 27902 16916 27958
rect 16972 27902 17008 27958
rect 5436 27683 6933 27736
rect 5436 27631 5837 27683
rect 5993 27631 6765 27683
rect 6921 27631 6933 27683
rect 5436 27602 6933 27631
rect 8742 27695 8866 27735
rect 8742 27643 8778 27695
rect 8830 27643 8866 27695
rect 8742 27555 8866 27643
rect 13074 27683 14578 27736
rect 16880 27740 17008 27902
rect 13074 27631 13216 27683
rect 13372 27631 14144 27683
rect 14300 27631 14578 27683
rect 13074 27602 14578 27631
rect 16121 27695 16245 27735
rect 16121 27643 16157 27695
rect 16209 27643 16245 27695
rect 16880 27684 16916 27740
rect 16972 27684 17008 27740
rect 16880 27646 17008 27684
rect 17113 28041 17334 28305
rect 17113 27989 17151 28041
rect 17203 27989 17334 28041
rect 17113 27823 17334 27989
rect 17113 27771 17151 27823
rect 17203 27771 17334 27823
rect 16121 27555 16245 27643
rect 17113 27605 17334 27771
rect 8739 27477 8868 27555
rect 8100 27431 8224 27432
rect 5611 27417 5735 27418
rect 5887 27417 6011 27418
rect 1618 27355 1746 27392
rect 1618 27299 1654 27355
rect 1710 27299 1746 27355
rect 1618 27137 1746 27299
rect 1618 27081 1654 27137
rect 1710 27081 1746 27137
rect 1618 26919 1746 27081
rect 1618 26863 1654 26919
rect 1710 26863 1746 26919
rect 1618 26825 1746 26863
rect 2066 27355 2194 27392
rect 2066 27299 2102 27355
rect 2158 27299 2194 27355
rect 2066 27137 2194 27299
rect 2066 27081 2102 27137
rect 2158 27081 2194 27137
rect 2066 26919 2194 27081
rect 2066 26863 2102 26919
rect 2158 26863 2194 26919
rect 2066 26825 2194 26863
rect 2514 27355 2642 27392
rect 2514 27299 2550 27355
rect 2606 27299 2642 27355
rect 2514 27137 2642 27299
rect 2514 27081 2550 27137
rect 2606 27081 2642 27137
rect 2514 26919 2642 27081
rect 2514 26863 2550 26919
rect 2606 26863 2642 26919
rect 2514 26825 2642 26863
rect 2962 27355 3090 27392
rect 2962 27299 2998 27355
rect 3054 27299 3090 27355
rect 2962 27137 3090 27299
rect 2962 27081 2998 27137
rect 3054 27081 3090 27137
rect 2962 26919 3090 27081
rect 2962 26863 2998 26919
rect 3054 26863 3090 26919
rect 2962 26825 3090 26863
rect 3410 27355 3538 27392
rect 3410 27299 3446 27355
rect 3502 27299 3538 27355
rect 3410 27137 3538 27299
rect 3410 27081 3446 27137
rect 3502 27081 3538 27137
rect 3410 26919 3538 27081
rect 3410 26863 3446 26919
rect 3502 26863 3538 26919
rect 3410 26825 3538 26863
rect 3858 27355 3986 27392
rect 3858 27299 3894 27355
rect 3950 27299 3986 27355
rect 3858 27137 3986 27299
rect 3858 27081 3894 27137
rect 3950 27081 3986 27137
rect 3858 26919 3986 27081
rect 3858 26863 3894 26919
rect 3950 26863 3986 26919
rect 3858 26825 3986 26863
rect 4306 27355 4434 27392
rect 4306 27299 4342 27355
rect 4398 27299 4434 27355
rect 4306 27137 4434 27299
rect 4306 27081 4342 27137
rect 4398 27081 4434 27137
rect 4306 26919 4434 27081
rect 4306 26863 4342 26919
rect 4398 26863 4434 26919
rect 4306 26825 4434 26863
rect 4754 27355 4882 27392
rect 4754 27299 4790 27355
rect 4846 27299 4882 27355
rect 4754 27137 4882 27299
rect 4754 27081 4790 27137
rect 4846 27081 4882 27137
rect 4754 26919 4882 27081
rect 4754 26863 4790 26919
rect 4846 26863 4882 26919
rect 4754 26825 4882 26863
rect 5202 27355 5330 27392
rect 5202 27299 5238 27355
rect 5294 27299 5330 27355
rect 5202 27137 5330 27299
rect 5202 27081 5238 27137
rect 5294 27081 5330 27137
rect 5202 26919 5330 27081
rect 5202 26863 5238 26919
rect 5294 26863 5330 26919
rect 5202 26825 5330 26863
rect 5609 27380 5737 27417
rect 5609 27324 5645 27380
rect 5701 27324 5737 27380
rect 5609 27162 5737 27324
rect 5609 27106 5645 27162
rect 5701 27106 5737 27162
rect 5609 26944 5737 27106
rect 5609 26888 5645 26944
rect 5701 26888 5737 26944
rect 5609 26850 5737 26888
rect 5885 27380 6013 27417
rect 5885 27324 5921 27380
rect 5977 27324 6013 27380
rect 5885 27162 6013 27324
rect 8098 27394 8226 27431
rect 8098 27338 8134 27394
rect 8190 27338 8226 27394
rect 5885 27106 5921 27162
rect 5977 27106 6013 27162
rect 6969 27212 7309 27251
rect 6969 27156 7005 27212
rect 7061 27156 7217 27212
rect 7273 27156 7309 27212
rect 6969 27117 7309 27156
rect 8098 27176 8226 27338
rect 8098 27120 8134 27176
rect 8190 27120 8226 27176
rect 5885 26944 6013 27106
rect 5885 26888 5921 26944
rect 5977 26888 6013 26944
rect 5885 26850 6013 26888
rect 6968 26974 7307 27015
rect 6968 26922 7005 26974
rect 7057 26922 7217 26974
rect 7269 26922 7307 26974
rect 6968 26882 7307 26922
rect 8098 26958 8226 27120
rect 8098 26902 8134 26958
rect 8190 26902 8226 26958
rect 7072 26881 7202 26882
rect 5836 26516 6171 26554
rect 5836 26460 5872 26516
rect 5928 26460 6079 26516
rect 6135 26460 6171 26516
rect 5836 26298 6171 26460
rect 5836 26242 5872 26298
rect 5928 26242 6079 26298
rect 6135 26242 6171 26298
rect 5836 26080 6171 26242
rect 5836 26024 5872 26080
rect 5928 26024 6079 26080
rect 6135 26024 6171 26080
rect 5836 25862 6171 26024
rect 5836 25806 5872 25862
rect 5928 25806 6079 25862
rect 6135 25806 6171 25862
rect 5836 25768 6171 25806
rect 6563 26493 6691 26530
rect 6563 26437 6599 26493
rect 6655 26437 6691 26493
rect 6563 26275 6691 26437
rect 6563 26219 6599 26275
rect 6655 26219 6691 26275
rect 6563 26057 6691 26219
rect 6563 26001 6599 26057
rect 6655 26001 6691 26057
rect 6563 25839 6691 26001
rect 6563 25783 6599 25839
rect 6655 25783 6691 25839
rect 6563 25745 6691 25783
rect 5836 25221 6176 25262
rect 5836 25169 5874 25221
rect 5926 25169 6086 25221
rect 6138 25169 6176 25221
rect 5836 25129 6176 25169
rect 1779 24775 1907 24813
rect 1779 24719 1815 24775
rect 1871 24719 1907 24775
rect 1779 24558 1907 24719
rect 1779 24502 1815 24558
rect 1871 24502 1907 24558
rect 1779 24340 1907 24502
rect 1779 24284 1815 24340
rect 1871 24284 1907 24340
rect 1779 24123 1907 24284
rect 1779 24067 1815 24123
rect 1871 24067 1907 24123
rect 1779 23905 1907 24067
rect 1779 23849 1815 23905
rect 1871 23849 1907 23905
rect 1779 23687 1907 23849
rect 1779 23631 1815 23687
rect 1871 23631 1907 23687
rect 1779 23469 1907 23631
rect 1779 23413 1815 23469
rect 1871 23413 1907 23469
rect 1779 23252 1907 23413
rect 1779 23196 1815 23252
rect 1871 23196 1907 23252
rect 1779 23034 1907 23196
rect 1779 22978 1815 23034
rect 1871 22978 1907 23034
rect 1779 22817 1907 22978
rect 1779 22761 1815 22817
rect 1871 22761 1907 22817
rect 1779 22722 1907 22761
rect 2230 24775 2926 24841
rect 2230 24719 2267 24775
rect 2323 24719 2550 24775
rect 2606 24719 2833 24775
rect 2889 24719 2926 24775
rect 2230 24558 2926 24719
rect 2230 24502 2267 24558
rect 2323 24502 2550 24558
rect 2606 24502 2833 24558
rect 2889 24502 2926 24558
rect 2230 24340 2926 24502
rect 2230 24284 2267 24340
rect 2323 24284 2550 24340
rect 2606 24284 2833 24340
rect 2889 24284 2926 24340
rect 2230 24123 2926 24284
rect 2230 24067 2267 24123
rect 2323 24067 2550 24123
rect 2606 24067 2833 24123
rect 2889 24067 2926 24123
rect 2230 23905 2926 24067
rect 2230 23849 2267 23905
rect 2323 23849 2550 23905
rect 2606 23849 2833 23905
rect 2889 23849 2926 23905
rect 2230 23687 2926 23849
rect 2230 23631 2267 23687
rect 2323 23631 2550 23687
rect 2606 23631 2833 23687
rect 2889 23631 2926 23687
rect 2230 23469 2926 23631
rect 2230 23413 2267 23469
rect 2323 23413 2550 23469
rect 2606 23413 2833 23469
rect 2889 23413 2926 23469
rect 2230 23252 2926 23413
rect 2230 23196 2267 23252
rect 2323 23196 2550 23252
rect 2606 23196 2833 23252
rect 2889 23196 2926 23252
rect 2230 23034 2926 23196
rect 2230 22978 2267 23034
rect 2323 22978 2550 23034
rect 2606 22978 2833 23034
rect 2889 22978 2926 23034
rect 2230 22817 2926 22978
rect 2230 22761 2267 22817
rect 2323 22761 2550 22817
rect 2606 22761 2833 22817
rect 2889 22761 2926 22817
rect 2230 22722 2926 22761
rect 3249 24775 3377 24813
rect 3249 24719 3285 24775
rect 3341 24719 3377 24775
rect 3249 24558 3377 24719
rect 3249 24502 3285 24558
rect 3341 24502 3377 24558
rect 3249 24340 3377 24502
rect 3249 24284 3285 24340
rect 3341 24284 3377 24340
rect 3249 24123 3377 24284
rect 3249 24067 3285 24123
rect 3341 24067 3377 24123
rect 3249 23905 3377 24067
rect 3249 23849 3285 23905
rect 3341 23849 3377 23905
rect 3249 23687 3377 23849
rect 3249 23631 3285 23687
rect 3341 23631 3377 23687
rect 3249 23469 3377 23631
rect 3249 23413 3285 23469
rect 3341 23413 3377 23469
rect 3249 23252 3377 23413
rect 3249 23196 3285 23252
rect 3341 23196 3377 23252
rect 3249 23034 3377 23196
rect 3249 22978 3285 23034
rect 3341 22978 3377 23034
rect 3249 22817 3377 22978
rect 3249 22761 3285 22817
rect 3341 22761 3377 22817
rect 3249 22722 3377 22761
rect 3571 24775 3699 24813
rect 3571 24719 3607 24775
rect 3663 24719 3699 24775
rect 3571 24558 3699 24719
rect 3571 24502 3607 24558
rect 3663 24502 3699 24558
rect 3571 24340 3699 24502
rect 3571 24284 3607 24340
rect 3663 24284 3699 24340
rect 3571 24123 3699 24284
rect 3571 24067 3607 24123
rect 3663 24067 3699 24123
rect 3571 23905 3699 24067
rect 3571 23849 3607 23905
rect 3663 23849 3699 23905
rect 3571 23687 3699 23849
rect 3571 23631 3607 23687
rect 3663 23631 3699 23687
rect 3571 23469 3699 23631
rect 3571 23413 3607 23469
rect 3663 23413 3699 23469
rect 3571 23252 3699 23413
rect 3571 23196 3607 23252
rect 3663 23196 3699 23252
rect 3571 23034 3699 23196
rect 3571 22978 3607 23034
rect 3663 22978 3699 23034
rect 3571 22817 3699 22978
rect 3571 22761 3607 22817
rect 3663 22761 3699 22817
rect 3571 22722 3699 22761
rect 4022 24775 4718 24841
rect 4022 24719 4059 24775
rect 4115 24719 4342 24775
rect 4398 24719 4625 24775
rect 4681 24719 4718 24775
rect 4022 24558 4718 24719
rect 4022 24502 4059 24558
rect 4115 24502 4342 24558
rect 4398 24502 4625 24558
rect 4681 24502 4718 24558
rect 4022 24340 4718 24502
rect 4022 24284 4059 24340
rect 4115 24284 4342 24340
rect 4398 24284 4625 24340
rect 4681 24284 4718 24340
rect 4022 24123 4718 24284
rect 4022 24067 4059 24123
rect 4115 24067 4342 24123
rect 4398 24067 4625 24123
rect 4681 24067 4718 24123
rect 4022 23905 4718 24067
rect 4022 23849 4059 23905
rect 4115 23849 4342 23905
rect 4398 23849 4625 23905
rect 4681 23849 4718 23905
rect 4022 23687 4718 23849
rect 4022 23631 4059 23687
rect 4115 23631 4342 23687
rect 4398 23631 4625 23687
rect 4681 23631 4718 23687
rect 4022 23469 4718 23631
rect 4022 23413 4059 23469
rect 4115 23413 4342 23469
rect 4398 23413 4625 23469
rect 4681 23413 4718 23469
rect 4022 23252 4718 23413
rect 4022 23196 4059 23252
rect 4115 23196 4342 23252
rect 4398 23196 4625 23252
rect 4681 23196 4718 23252
rect 4022 23034 4718 23196
rect 4022 22978 4059 23034
rect 4115 22978 4342 23034
rect 4398 22978 4625 23034
rect 4681 22978 4718 23034
rect 4022 22817 4718 22978
rect 4022 22761 4059 22817
rect 4115 22761 4342 22817
rect 4398 22761 4625 22817
rect 4681 22761 4718 22817
rect 4022 22722 4718 22761
rect 5041 24775 5169 24813
rect 5041 24719 5077 24775
rect 5133 24719 5169 24775
rect 5041 24558 5169 24719
rect 5041 24502 5077 24558
rect 5133 24502 5169 24558
rect 5041 24340 5169 24502
rect 5041 24284 5077 24340
rect 5133 24284 5169 24340
rect 5041 24123 5169 24284
rect 5041 24067 5077 24123
rect 5133 24067 5169 24123
rect 5041 23905 5169 24067
rect 5041 23849 5077 23905
rect 5133 23849 5169 23905
rect 5041 23687 5169 23849
rect 5041 23631 5077 23687
rect 5133 23631 5169 23687
rect 5041 23469 5169 23631
rect 5041 23413 5077 23469
rect 5133 23413 5169 23469
rect 5041 23252 5169 23413
rect 5041 23196 5077 23252
rect 5133 23196 5169 23252
rect 5041 23034 5169 23196
rect 5041 22978 5077 23034
rect 5133 22978 5169 23034
rect 5041 22817 5169 22978
rect 5041 22761 5077 22817
rect 5133 22761 5169 22817
rect 5041 22722 5169 22761
rect 1776 21842 2128 21882
rect 1776 21790 2039 21842
rect 2091 21790 2128 21842
rect 1776 21624 2128 21790
rect 1776 21572 2039 21624
rect 2091 21572 2128 21624
rect 1776 21531 2128 21572
rect 3028 21842 3380 21882
rect 3028 21790 3065 21842
rect 3117 21790 3380 21842
rect 3028 21624 3380 21790
rect 3028 21572 3065 21624
rect 3117 21572 3380 21624
rect 3028 21531 3380 21572
rect 1776 20502 1904 21531
rect 1776 20450 1814 20502
rect 1866 20450 1904 20502
rect 1776 20284 1904 20450
rect 1776 20232 1814 20284
rect 1866 20232 1904 20284
rect 1776 20196 1904 20232
rect 2230 20366 2926 20542
rect 2230 20310 2267 20366
rect 2323 20310 2550 20366
rect 2606 20310 2833 20366
rect 2889 20310 2926 20366
rect 1776 20067 1903 20196
rect 1776 20015 1814 20067
rect 1866 20015 1903 20067
rect 1776 19849 1903 20015
rect 1776 19797 1814 19849
rect 1866 19797 1903 19849
rect 1776 19631 1903 19797
rect 1776 19579 1814 19631
rect 1866 19579 1903 19631
rect 1776 19413 1903 19579
rect 1776 19361 1814 19413
rect 1866 19361 1903 19413
rect 1776 19196 1903 19361
rect 1776 19144 1814 19196
rect 1866 19144 1903 19196
rect 1776 18978 1903 19144
rect 1776 18926 1814 18978
rect 1866 18926 1903 18978
rect 1776 18886 1903 18926
rect 2230 20148 2926 20310
rect 3252 20502 3380 21531
rect 3252 20450 3290 20502
rect 3342 20450 3380 20502
rect 3252 20284 3380 20450
rect 3252 20232 3290 20284
rect 3342 20232 3380 20284
rect 3252 20196 3380 20232
rect 2230 20092 2267 20148
rect 2323 20092 2550 20148
rect 2606 20092 2833 20148
rect 2889 20092 2926 20148
rect 2230 19930 2926 20092
rect 2230 19874 2267 19930
rect 2323 19874 2550 19930
rect 2606 19874 2833 19930
rect 2889 19874 2926 19930
rect 2230 19711 2926 19874
rect 2230 19659 2269 19711
rect 2321 19659 2552 19711
rect 2604 19659 2835 19711
rect 2887 19659 2926 19711
rect 2230 19494 2926 19659
rect 2230 19442 2269 19494
rect 2321 19442 2552 19494
rect 2604 19442 2835 19494
rect 2887 19442 2926 19494
rect 2230 19276 2926 19442
rect 2230 19224 2269 19276
rect 2321 19224 2552 19276
rect 2604 19224 2835 19276
rect 2887 19224 2926 19276
rect 2230 19058 2926 19224
rect 2230 19006 2269 19058
rect 2321 19006 2552 19058
rect 2604 19006 2835 19058
rect 2887 19006 2926 19058
rect 2230 18840 2926 19006
rect 3253 20067 3380 20196
rect 3253 20015 3290 20067
rect 3342 20015 3380 20067
rect 3253 19849 3380 20015
rect 3253 19797 3290 19849
rect 3342 19797 3380 19849
rect 3253 19631 3380 19797
rect 3253 19579 3290 19631
rect 3342 19579 3380 19631
rect 3253 19413 3380 19579
rect 3253 19361 3290 19413
rect 3342 19361 3380 19413
rect 3253 19196 3380 19361
rect 3253 19144 3290 19196
rect 3342 19144 3380 19196
rect 3253 18978 3380 19144
rect 3253 18926 3290 18978
rect 3342 18926 3380 18978
rect 3253 18886 3380 18926
rect 3568 21842 3920 21882
rect 3568 21790 3831 21842
rect 3883 21790 3920 21842
rect 3568 21624 3920 21790
rect 3568 21572 3831 21624
rect 3883 21572 3920 21624
rect 3568 21531 3920 21572
rect 4820 21842 5172 21882
rect 4820 21790 4857 21842
rect 4909 21790 5172 21842
rect 4820 21624 5172 21790
rect 4820 21572 4857 21624
rect 4909 21572 5172 21624
rect 4820 21531 5172 21572
rect 3568 20502 3696 21531
rect 3568 20450 3606 20502
rect 3658 20450 3696 20502
rect 3568 20284 3696 20450
rect 3568 20232 3606 20284
rect 3658 20232 3696 20284
rect 3568 20196 3696 20232
rect 4022 20366 4718 20542
rect 4022 20310 4059 20366
rect 4115 20310 4342 20366
rect 4398 20310 4625 20366
rect 4681 20310 4718 20366
rect 3568 20067 3695 20196
rect 3568 20015 3606 20067
rect 3658 20015 3695 20067
rect 3568 19849 3695 20015
rect 3568 19797 3606 19849
rect 3658 19797 3695 19849
rect 3568 19631 3695 19797
rect 3568 19579 3606 19631
rect 3658 19579 3695 19631
rect 3568 19413 3695 19579
rect 3568 19361 3606 19413
rect 3658 19361 3695 19413
rect 3568 19196 3695 19361
rect 3568 19144 3606 19196
rect 3658 19144 3695 19196
rect 3568 18978 3695 19144
rect 3568 18926 3606 18978
rect 3658 18926 3695 18978
rect 3568 18886 3695 18926
rect 4022 20148 4718 20310
rect 5044 20502 5172 21531
rect 5044 20450 5082 20502
rect 5134 20450 5172 20502
rect 5044 20284 5172 20450
rect 5044 20232 5082 20284
rect 5134 20232 5172 20284
rect 5044 20196 5172 20232
rect 4022 20092 4059 20148
rect 4115 20092 4342 20148
rect 4398 20092 4625 20148
rect 4681 20092 4718 20148
rect 4022 19930 4718 20092
rect 4022 19874 4059 19930
rect 4115 19874 4342 19930
rect 4398 19874 4625 19930
rect 4681 19874 4718 19930
rect 4022 19711 4718 19874
rect 4022 19659 4061 19711
rect 4113 19659 4344 19711
rect 4396 19659 4627 19711
rect 4679 19659 4718 19711
rect 4022 19494 4718 19659
rect 4022 19442 4061 19494
rect 4113 19442 4344 19494
rect 4396 19442 4627 19494
rect 4679 19442 4718 19494
rect 4022 19276 4718 19442
rect 4022 19224 4061 19276
rect 4113 19224 4344 19276
rect 4396 19224 4627 19276
rect 4679 19224 4718 19276
rect 4022 19058 4718 19224
rect 4022 19006 4061 19058
rect 4113 19006 4344 19058
rect 4396 19006 4627 19058
rect 4679 19006 4718 19058
rect 2230 18788 2269 18840
rect 2321 18788 2552 18840
rect 2604 18788 2835 18840
rect 2887 18788 2926 18840
rect 2230 18623 2926 18788
rect 2230 18571 2269 18623
rect 2321 18571 2552 18623
rect 2604 18571 2835 18623
rect 2887 18571 2926 18623
rect 2230 18408 2926 18571
rect 2230 18352 2267 18408
rect 2323 18352 2550 18408
rect 2606 18352 2833 18408
rect 2889 18352 2926 18408
rect 2230 18190 2926 18352
rect 2230 18134 2267 18190
rect 2323 18134 2550 18190
rect 2606 18134 2833 18190
rect 2889 18134 2926 18190
rect 2230 17972 2926 18134
rect 2230 17916 2267 17972
rect 2323 17916 2550 17972
rect 2606 17916 2833 17972
rect 2889 17916 2926 17972
rect 2230 17754 2926 17916
rect 2230 17698 2267 17754
rect 2323 17698 2550 17754
rect 2606 17698 2833 17754
rect 2889 17698 2926 17754
rect 2230 17657 2926 17698
rect 4022 18840 4718 19006
rect 5045 20067 5172 20196
rect 5045 20015 5082 20067
rect 5134 20015 5172 20067
rect 5045 19849 5172 20015
rect 5045 19797 5082 19849
rect 5134 19797 5172 19849
rect 5045 19631 5172 19797
rect 5045 19579 5082 19631
rect 5134 19579 5172 19631
rect 5045 19413 5172 19579
rect 5836 19837 5965 25129
rect 6056 24804 6184 24842
rect 6056 24748 6092 24804
rect 6148 24748 6184 24804
rect 6056 24587 6184 24748
rect 6056 24531 6092 24587
rect 6148 24531 6184 24587
rect 6056 24369 6184 24531
rect 6056 24313 6092 24369
rect 6148 24313 6184 24369
rect 6056 24152 6184 24313
rect 6056 24096 6092 24152
rect 6148 24096 6184 24152
rect 6056 23934 6184 24096
rect 6056 23878 6092 23934
rect 6148 23878 6184 23934
rect 6056 23716 6184 23878
rect 6056 23660 6092 23716
rect 6148 23660 6184 23716
rect 6056 23498 6184 23660
rect 6056 23442 6092 23498
rect 6148 23442 6184 23498
rect 6056 23281 6184 23442
rect 6056 23225 6092 23281
rect 6148 23225 6184 23281
rect 6056 23063 6184 23225
rect 6570 24813 6698 24851
rect 6570 24757 6606 24813
rect 6662 24757 6698 24813
rect 6570 24595 6698 24757
rect 6570 24539 6606 24595
rect 6662 24539 6698 24595
rect 6570 24378 6698 24539
rect 6570 24322 6606 24378
rect 6662 24322 6698 24378
rect 6570 24160 6698 24322
rect 6570 24104 6606 24160
rect 6662 24104 6698 24160
rect 6570 23942 6698 24104
rect 6570 23886 6606 23942
rect 6662 23886 6698 23942
rect 6570 23724 6698 23886
rect 6570 23668 6606 23724
rect 6662 23668 6698 23724
rect 6570 23507 6698 23668
rect 6570 23451 6606 23507
rect 6662 23451 6698 23507
rect 6570 23289 6698 23451
rect 6570 23233 6606 23289
rect 6662 23233 6698 23289
rect 6570 23195 6698 23233
rect 6056 23007 6092 23063
rect 6148 23007 6184 23063
rect 7072 23054 7201 26881
rect 8098 26864 8226 26902
rect 8739 27425 8778 27477
rect 8830 27425 8868 27477
rect 16118 27477 16247 27555
rect 17113 27553 17151 27605
rect 17203 27553 17334 27605
rect 17113 27512 17334 27553
rect 17464 28041 17685 28998
rect 17464 27989 17595 28041
rect 17647 27989 17685 28041
rect 17464 27823 17685 27989
rect 17464 27771 17595 27823
rect 17647 27771 17685 27823
rect 17464 27605 17685 27771
rect 17790 28394 17918 28431
rect 17790 28338 17826 28394
rect 17882 28338 17918 28394
rect 17790 28176 17918 28338
rect 17790 28120 17826 28176
rect 17882 28120 17918 28176
rect 17790 27958 17918 28120
rect 17790 27902 17826 27958
rect 17882 27902 17918 27958
rect 17790 27740 17918 27902
rect 17790 27684 17826 27740
rect 17882 27684 17918 27740
rect 17790 27646 17918 27684
rect 18514 28394 18642 28431
rect 18514 28338 18550 28394
rect 18606 28338 18642 28394
rect 18514 28176 18642 28338
rect 18746 28305 18968 28998
rect 18514 28120 18550 28176
rect 18606 28120 18642 28176
rect 18514 27958 18642 28120
rect 18514 27902 18550 27958
rect 18606 27902 18642 27958
rect 18514 27740 18642 27902
rect 18514 27684 18550 27740
rect 18606 27684 18642 27740
rect 18514 27646 18642 27684
rect 18747 28041 18968 28305
rect 18747 27989 18785 28041
rect 18837 27989 18968 28041
rect 18747 27823 18968 27989
rect 18747 27771 18785 27823
rect 18837 27771 18968 27823
rect 17464 27553 17595 27605
rect 17647 27553 17685 27605
rect 17464 27512 17685 27553
rect 18747 27605 18968 27771
rect 18747 27553 18785 27605
rect 18837 27553 18968 27605
rect 18747 27512 18968 27553
rect 19098 28041 19319 28998
rect 19098 27989 19229 28041
rect 19281 27989 19319 28041
rect 19098 27823 19319 27989
rect 19098 27771 19229 27823
rect 19281 27771 19319 27823
rect 19098 27605 19319 27771
rect 19424 28394 19552 28431
rect 19424 28338 19460 28394
rect 19516 28338 19552 28394
rect 19424 28176 19552 28338
rect 19424 28120 19460 28176
rect 19516 28120 19552 28176
rect 19424 27958 19552 28120
rect 19424 27902 19460 27958
rect 19516 27902 19552 27958
rect 19424 27740 19552 27902
rect 19424 27684 19460 27740
rect 19516 27684 19552 27740
rect 19424 27646 19552 27684
rect 20147 28394 20275 28431
rect 20147 28338 20183 28394
rect 20239 28338 20275 28394
rect 20147 28176 20275 28338
rect 20147 28120 20183 28176
rect 20239 28120 20275 28176
rect 20147 27958 20275 28120
rect 20147 27902 20183 27958
rect 20239 27902 20275 27958
rect 20147 27740 20275 27902
rect 20147 27684 20183 27740
rect 20239 27684 20275 27740
rect 20147 27646 20275 27684
rect 20380 28305 20602 28998
rect 20731 28305 20953 28998
rect 21057 28394 21185 28431
rect 21057 28338 21093 28394
rect 21149 28338 21185 28394
rect 20380 28041 20601 28305
rect 20380 27989 20418 28041
rect 20470 27989 20601 28041
rect 20380 27823 20601 27989
rect 20380 27771 20418 27823
rect 20470 27771 20601 27823
rect 19098 27553 19229 27605
rect 19281 27553 19319 27605
rect 19098 27512 19319 27553
rect 20380 27605 20601 27771
rect 20380 27553 20418 27605
rect 20470 27553 20601 27605
rect 20380 27512 20601 27553
rect 20731 28041 20952 28305
rect 20731 27989 20862 28041
rect 20914 27989 20952 28041
rect 20731 27823 20952 27989
rect 20731 27771 20862 27823
rect 20914 27771 20952 27823
rect 20731 27605 20952 27771
rect 21057 28176 21185 28338
rect 21057 28120 21093 28176
rect 21149 28120 21185 28176
rect 21057 27958 21185 28120
rect 21057 27902 21093 27958
rect 21149 27902 21185 27958
rect 21057 27740 21185 27902
rect 21057 27684 21093 27740
rect 21149 27684 21185 27740
rect 21057 27646 21185 27684
rect 21781 28394 21909 28431
rect 21781 28338 21817 28394
rect 21873 28338 21909 28394
rect 21781 28176 21909 28338
rect 21781 28120 21817 28176
rect 21873 28120 21909 28176
rect 21781 27958 21909 28120
rect 21781 27902 21817 27958
rect 21873 27902 21909 27958
rect 21781 27740 21909 27902
rect 21781 27684 21817 27740
rect 21873 27684 21909 27740
rect 21781 27646 21909 27684
rect 22014 28041 22235 28998
rect 22014 27989 22052 28041
rect 22104 27989 22235 28041
rect 22014 27823 22235 27989
rect 22014 27771 22052 27823
rect 22104 27771 22235 27823
rect 20731 27553 20862 27605
rect 20914 27553 20952 27605
rect 20731 27512 20952 27553
rect 22014 27605 22235 27771
rect 22014 27553 22052 27605
rect 22104 27553 22235 27605
rect 22014 27512 22235 27553
rect 22365 28305 22587 28998
rect 22691 28394 22819 28431
rect 22691 28338 22727 28394
rect 22783 28338 22819 28394
rect 22365 28041 22586 28305
rect 22365 27989 22496 28041
rect 22548 27989 22586 28041
rect 22365 27823 22586 27989
rect 22365 27771 22496 27823
rect 22548 27771 22586 27823
rect 22365 27605 22586 27771
rect 22691 28176 22819 28338
rect 22691 28120 22727 28176
rect 22783 28120 22819 28176
rect 22691 27958 22819 28120
rect 22691 27902 22727 27958
rect 22783 27902 22819 27958
rect 22691 27740 22819 27902
rect 22691 27684 22727 27740
rect 22783 27684 22819 27740
rect 22691 27646 22819 27684
rect 23301 27736 23654 29316
rect 28532 30026 29412 30125
rect 28532 29970 28627 30026
rect 28683 29970 28838 30026
rect 28894 29970 29050 30026
rect 29106 29970 29261 30026
rect 29317 29970 29412 30026
rect 28532 29808 29412 29970
rect 28532 29752 28627 29808
rect 28683 29752 28838 29808
rect 28894 29752 29050 29808
rect 29106 29752 29261 29808
rect 29317 29752 29412 29808
rect 28532 29590 29412 29752
rect 28532 29534 28627 29590
rect 28683 29534 28838 29590
rect 28894 29534 29050 29590
rect 29106 29534 29261 29590
rect 29317 29534 29412 29590
rect 28532 29372 29412 29534
rect 28532 29316 28627 29372
rect 28683 29316 28838 29372
rect 28894 29316 29050 29372
rect 29106 29316 29261 29372
rect 29317 29316 29412 29372
rect 24409 29037 24534 29038
rect 24408 28999 24537 29037
rect 24408 28943 24444 28999
rect 24500 28943 24537 28999
rect 24408 28781 24537 28943
rect 24408 28725 24444 28781
rect 24500 28725 24537 28781
rect 23749 28403 23877 28440
rect 23749 28347 23785 28403
rect 23841 28347 23877 28403
rect 23749 28185 23877 28347
rect 23749 28129 23785 28185
rect 23841 28129 23877 28185
rect 23749 27967 23877 28129
rect 23749 27911 23785 27967
rect 23841 27911 23877 27967
rect 23749 27873 23877 27911
rect 24188 28403 24316 28440
rect 24188 28347 24224 28403
rect 24280 28347 24316 28403
rect 24188 28185 24316 28347
rect 24188 28129 24224 28185
rect 24280 28129 24316 28185
rect 24188 27967 24316 28129
rect 24188 27911 24224 27967
rect 24280 27911 24316 27967
rect 24188 27873 24316 27911
rect 24408 28185 24537 28725
rect 24408 28133 24446 28185
rect 24498 28133 24537 28185
rect 24408 27967 24537 28133
rect 24408 27915 24446 27967
rect 24498 27915 24537 27967
rect 24408 27874 24537 27915
rect 25572 28346 25700 28383
rect 25572 28290 25608 28346
rect 25664 28290 25700 28346
rect 25572 28128 25700 28290
rect 25572 28072 25608 28128
rect 25664 28072 25700 28128
rect 25572 27910 25700 28072
rect 25572 27854 25608 27910
rect 25664 27854 25700 27910
rect 25572 27816 25700 27854
rect 23301 27695 24791 27736
rect 22365 27553 22496 27605
rect 22548 27553 22586 27605
rect 23301 27643 23598 27695
rect 23650 27643 23810 27695
rect 23862 27673 24791 27695
rect 23862 27643 24572 27673
rect 23301 27621 24572 27643
rect 24728 27621 24791 27673
rect 23301 27602 24791 27621
rect 26606 27686 26730 27726
rect 26606 27634 26642 27686
rect 26694 27634 26730 27686
rect 22365 27512 22586 27553
rect 26606 27545 26730 27634
rect 15479 27431 15603 27432
rect 7527 26516 7862 26554
rect 7527 26460 7563 26516
rect 7619 26460 7770 26516
rect 7826 26460 7862 26516
rect 7527 26298 7862 26460
rect 7527 26242 7563 26298
rect 7619 26242 7770 26298
rect 7826 26242 7862 26298
rect 7527 26080 7862 26242
rect 7527 26024 7563 26080
rect 7619 26024 7770 26080
rect 7826 26024 7862 26080
rect 7527 25862 7862 26024
rect 7527 25806 7563 25862
rect 7619 25806 7770 25862
rect 7826 25806 7862 25862
rect 7527 25768 7862 25806
rect 8254 26493 8382 26530
rect 8254 26437 8290 26493
rect 8346 26437 8382 26493
rect 8254 26275 8382 26437
rect 8254 26219 8290 26275
rect 8346 26219 8382 26275
rect 8254 26057 8382 26219
rect 8254 26001 8290 26057
rect 8346 26001 8382 26057
rect 8254 25839 8382 26001
rect 8254 25783 8290 25839
rect 8346 25783 8382 25839
rect 8254 25745 8382 25783
rect 6056 22846 6184 23007
rect 6056 22790 6092 22846
rect 6148 22790 6184 22846
rect 6056 22751 6184 22790
rect 6558 22921 7201 23054
rect 7527 25221 7867 25262
rect 7527 25169 7565 25221
rect 7617 25169 7777 25221
rect 7829 25169 7867 25221
rect 7527 25129 7867 25169
rect 6275 21796 6399 21836
rect 6275 21744 6311 21796
rect 6363 21744 6399 21796
rect 6275 21578 6399 21744
rect 6275 21526 6311 21578
rect 6363 21526 6399 21578
rect 6275 21486 6399 21526
rect 6558 21567 6687 22921
rect 6558 21511 6595 21567
rect 6651 21511 6687 21567
rect 5836 19785 5874 19837
rect 5926 19785 5965 19837
rect 5836 19619 5965 19785
rect 5836 19572 5874 19619
rect 5838 19567 5874 19572
rect 5926 19572 5965 19619
rect 6558 21349 6687 21511
rect 6558 21293 6595 21349
rect 6651 21293 6687 21349
rect 6558 19626 6687 21293
rect 6787 22703 6916 22744
rect 6787 22651 6825 22703
rect 6877 22651 6916 22703
rect 6787 22485 6916 22651
rect 6787 22433 6825 22485
rect 6877 22433 6916 22485
rect 6787 21162 6916 22433
rect 7050 22043 7175 22082
rect 7050 21987 7085 22043
rect 7141 21987 7175 22043
rect 7050 21866 7175 21987
rect 6787 21110 6825 21162
rect 6877 21110 6916 21162
rect 6787 21069 6916 21110
rect 7048 21825 7177 21866
rect 7048 21769 7085 21825
rect 7141 21769 7177 21825
rect 7048 19828 7177 21769
rect 7527 19837 7656 25129
rect 7747 24804 7875 24842
rect 7747 24748 7783 24804
rect 7839 24748 7875 24804
rect 7747 24587 7875 24748
rect 7747 24531 7783 24587
rect 7839 24531 7875 24587
rect 7747 24369 7875 24531
rect 7747 24313 7783 24369
rect 7839 24313 7875 24369
rect 7747 24152 7875 24313
rect 7747 24096 7783 24152
rect 7839 24096 7875 24152
rect 7747 23934 7875 24096
rect 7747 23878 7783 23934
rect 7839 23878 7875 23934
rect 7747 23716 7875 23878
rect 7747 23660 7783 23716
rect 7839 23660 7875 23716
rect 7747 23498 7875 23660
rect 7747 23442 7783 23498
rect 7839 23442 7875 23498
rect 7747 23281 7875 23442
rect 7747 23225 7783 23281
rect 7839 23225 7875 23281
rect 7747 23063 7875 23225
rect 8261 24813 8389 24851
rect 8261 24757 8297 24813
rect 8353 24757 8389 24813
rect 8261 24595 8389 24757
rect 8261 24539 8297 24595
rect 8353 24539 8389 24595
rect 8261 24378 8389 24539
rect 8261 24322 8297 24378
rect 8353 24322 8389 24378
rect 8261 24160 8389 24322
rect 8261 24104 8297 24160
rect 8353 24104 8389 24160
rect 8261 23942 8389 24104
rect 8261 23886 8297 23942
rect 8353 23886 8389 23942
rect 8261 23724 8389 23886
rect 8261 23668 8297 23724
rect 8353 23668 8389 23724
rect 8261 23507 8389 23668
rect 8261 23451 8297 23507
rect 8353 23451 8389 23507
rect 8261 23289 8389 23451
rect 8261 23233 8297 23289
rect 8353 23233 8389 23289
rect 8261 23195 8389 23233
rect 7747 23007 7783 23063
rect 7839 23007 7875 23063
rect 7747 22846 7875 23007
rect 7747 22790 7783 22846
rect 7839 22790 7875 22846
rect 7747 22751 7875 22790
rect 8478 22703 8607 22744
rect 8478 22651 8516 22703
rect 8568 22651 8607 22703
rect 8478 22485 8607 22651
rect 8478 22433 8516 22485
rect 8568 22433 8607 22485
rect 7964 21796 8093 21837
rect 7964 21744 8002 21796
rect 8054 21744 8093 21796
rect 7964 21578 8093 21744
rect 8251 21605 8376 21606
rect 7964 21526 8002 21578
rect 8054 21526 8093 21578
rect 7964 20960 8093 21526
rect 7964 20908 8002 20960
rect 8054 20908 8093 20960
rect 7964 20867 8093 20908
rect 8249 21567 8378 21605
rect 8249 21511 8286 21567
rect 8342 21511 8378 21567
rect 8249 21349 8378 21511
rect 8249 21293 8286 21349
rect 8342 21293 8378 21349
rect 7527 19785 7565 19837
rect 7617 19785 7656 19837
rect 5926 19567 5962 19572
rect 5838 19527 5962 19567
rect 6558 19493 7177 19626
rect 7527 19619 7656 19785
rect 7527 19572 7565 19619
rect 7529 19567 7565 19572
rect 7617 19572 7656 19619
rect 8249 19626 8378 21293
rect 8478 20758 8607 22433
rect 8478 20706 8516 20758
rect 8568 20706 8607 20758
rect 8478 20665 8607 20706
rect 8739 22043 8868 27425
rect 12990 27417 13114 27418
rect 13266 27417 13390 27418
rect 8997 27355 9125 27392
rect 8997 27299 9033 27355
rect 9089 27299 9125 27355
rect 8997 27137 9125 27299
rect 8997 27081 9033 27137
rect 9089 27081 9125 27137
rect 8997 26919 9125 27081
rect 8997 26863 9033 26919
rect 9089 26863 9125 26919
rect 8997 26825 9125 26863
rect 9445 27355 9573 27392
rect 9445 27299 9481 27355
rect 9537 27299 9573 27355
rect 9445 27137 9573 27299
rect 9445 27081 9481 27137
rect 9537 27081 9573 27137
rect 9445 26919 9573 27081
rect 9445 26863 9481 26919
rect 9537 26863 9573 26919
rect 9445 26825 9573 26863
rect 9893 27355 10021 27392
rect 9893 27299 9929 27355
rect 9985 27299 10021 27355
rect 9893 27137 10021 27299
rect 9893 27081 9929 27137
rect 9985 27081 10021 27137
rect 9893 26919 10021 27081
rect 9893 26863 9929 26919
rect 9985 26863 10021 26919
rect 9893 26825 10021 26863
rect 10341 27355 10469 27392
rect 10341 27299 10377 27355
rect 10433 27299 10469 27355
rect 10341 27137 10469 27299
rect 10341 27081 10377 27137
rect 10433 27081 10469 27137
rect 10341 26919 10469 27081
rect 10341 26863 10377 26919
rect 10433 26863 10469 26919
rect 10341 26825 10469 26863
rect 10789 27355 10917 27392
rect 10789 27299 10825 27355
rect 10881 27299 10917 27355
rect 10789 27137 10917 27299
rect 10789 27081 10825 27137
rect 10881 27081 10917 27137
rect 10789 26919 10917 27081
rect 10789 26863 10825 26919
rect 10881 26863 10917 26919
rect 10789 26825 10917 26863
rect 11237 27355 11365 27392
rect 11237 27299 11273 27355
rect 11329 27299 11365 27355
rect 11237 27137 11365 27299
rect 11237 27081 11273 27137
rect 11329 27081 11365 27137
rect 11237 26919 11365 27081
rect 11237 26863 11273 26919
rect 11329 26863 11365 26919
rect 11237 26825 11365 26863
rect 11685 27355 11813 27392
rect 11685 27299 11721 27355
rect 11777 27299 11813 27355
rect 11685 27137 11813 27299
rect 11685 27081 11721 27137
rect 11777 27081 11813 27137
rect 11685 26919 11813 27081
rect 11685 26863 11721 26919
rect 11777 26863 11813 26919
rect 11685 26825 11813 26863
rect 12133 27355 12261 27392
rect 12133 27299 12169 27355
rect 12225 27299 12261 27355
rect 12133 27137 12261 27299
rect 12133 27081 12169 27137
rect 12225 27081 12261 27137
rect 12133 26919 12261 27081
rect 12133 26863 12169 26919
rect 12225 26863 12261 26919
rect 12133 26825 12261 26863
rect 12581 27355 12709 27392
rect 12581 27299 12617 27355
rect 12673 27299 12709 27355
rect 12581 27137 12709 27299
rect 12581 27081 12617 27137
rect 12673 27081 12709 27137
rect 12581 26919 12709 27081
rect 12581 26863 12617 26919
rect 12673 26863 12709 26919
rect 12581 26825 12709 26863
rect 12988 27380 13116 27417
rect 12988 27324 13024 27380
rect 13080 27324 13116 27380
rect 12988 27162 13116 27324
rect 12988 27106 13024 27162
rect 13080 27106 13116 27162
rect 12988 26944 13116 27106
rect 12988 26888 13024 26944
rect 13080 26888 13116 26944
rect 12988 26850 13116 26888
rect 13264 27380 13392 27417
rect 13264 27324 13300 27380
rect 13356 27324 13392 27380
rect 13264 27162 13392 27324
rect 15477 27394 15605 27431
rect 15477 27338 15513 27394
rect 15569 27338 15605 27394
rect 13264 27106 13300 27162
rect 13356 27106 13392 27162
rect 14348 27212 14688 27251
rect 14348 27156 14384 27212
rect 14440 27156 14596 27212
rect 14652 27156 14688 27212
rect 14348 27117 14688 27156
rect 15477 27176 15605 27338
rect 15477 27120 15513 27176
rect 15569 27120 15605 27176
rect 13264 26944 13392 27106
rect 13264 26888 13300 26944
rect 13356 26888 13392 26944
rect 13264 26850 13392 26888
rect 14347 26974 14686 27015
rect 14347 26922 14384 26974
rect 14436 26922 14596 26974
rect 14648 26922 14686 26974
rect 14347 26882 14686 26922
rect 15477 26958 15605 27120
rect 15477 26902 15513 26958
rect 15569 26902 15605 26958
rect 14451 26881 14581 26882
rect 13215 26516 13550 26554
rect 13215 26460 13251 26516
rect 13307 26460 13458 26516
rect 13514 26460 13550 26516
rect 13215 26298 13550 26460
rect 13215 26242 13251 26298
rect 13307 26242 13458 26298
rect 13514 26242 13550 26298
rect 13215 26080 13550 26242
rect 13215 26024 13251 26080
rect 13307 26024 13458 26080
rect 13514 26024 13550 26080
rect 13215 25862 13550 26024
rect 13215 25806 13251 25862
rect 13307 25806 13458 25862
rect 13514 25806 13550 25862
rect 13215 25768 13550 25806
rect 13942 26493 14070 26530
rect 13942 26437 13978 26493
rect 14034 26437 14070 26493
rect 13942 26275 14070 26437
rect 13942 26219 13978 26275
rect 14034 26219 14070 26275
rect 13942 26057 14070 26219
rect 13942 26001 13978 26057
rect 14034 26001 14070 26057
rect 13942 25839 14070 26001
rect 13942 25783 13978 25839
rect 14034 25783 14070 25839
rect 13942 25745 14070 25783
rect 13215 25221 13555 25262
rect 13215 25169 13253 25221
rect 13305 25169 13465 25221
rect 13517 25169 13555 25221
rect 13215 25129 13555 25169
rect 9158 24775 9286 24813
rect 9158 24719 9194 24775
rect 9250 24719 9286 24775
rect 9158 24558 9286 24719
rect 9158 24502 9194 24558
rect 9250 24502 9286 24558
rect 9158 24340 9286 24502
rect 9158 24284 9194 24340
rect 9250 24284 9286 24340
rect 9158 24123 9286 24284
rect 9158 24067 9194 24123
rect 9250 24067 9286 24123
rect 9158 23905 9286 24067
rect 9158 23849 9194 23905
rect 9250 23849 9286 23905
rect 9158 23687 9286 23849
rect 9158 23631 9194 23687
rect 9250 23631 9286 23687
rect 9158 23469 9286 23631
rect 9158 23413 9194 23469
rect 9250 23413 9286 23469
rect 9158 23252 9286 23413
rect 9158 23196 9194 23252
rect 9250 23196 9286 23252
rect 9158 23034 9286 23196
rect 9158 22978 9194 23034
rect 9250 22978 9286 23034
rect 9158 22817 9286 22978
rect 9158 22761 9194 22817
rect 9250 22761 9286 22817
rect 9158 22722 9286 22761
rect 9609 24775 10305 24841
rect 9609 24719 9646 24775
rect 9702 24719 9929 24775
rect 9985 24719 10212 24775
rect 10268 24719 10305 24775
rect 9609 24558 10305 24719
rect 9609 24502 9646 24558
rect 9702 24502 9929 24558
rect 9985 24502 10212 24558
rect 10268 24502 10305 24558
rect 9609 24340 10305 24502
rect 9609 24284 9646 24340
rect 9702 24284 9929 24340
rect 9985 24284 10212 24340
rect 10268 24284 10305 24340
rect 9609 24123 10305 24284
rect 9609 24067 9646 24123
rect 9702 24067 9929 24123
rect 9985 24067 10212 24123
rect 10268 24067 10305 24123
rect 9609 23905 10305 24067
rect 9609 23849 9646 23905
rect 9702 23849 9929 23905
rect 9985 23849 10212 23905
rect 10268 23849 10305 23905
rect 9609 23687 10305 23849
rect 9609 23631 9646 23687
rect 9702 23631 9929 23687
rect 9985 23631 10212 23687
rect 10268 23631 10305 23687
rect 9609 23469 10305 23631
rect 9609 23413 9646 23469
rect 9702 23413 9929 23469
rect 9985 23413 10212 23469
rect 10268 23413 10305 23469
rect 9609 23252 10305 23413
rect 9609 23196 9646 23252
rect 9702 23196 9929 23252
rect 9985 23196 10212 23252
rect 10268 23196 10305 23252
rect 9609 23034 10305 23196
rect 9609 22978 9646 23034
rect 9702 22978 9929 23034
rect 9985 22978 10212 23034
rect 10268 22978 10305 23034
rect 9609 22817 10305 22978
rect 9609 22761 9646 22817
rect 9702 22761 9929 22817
rect 9985 22761 10212 22817
rect 10268 22761 10305 22817
rect 9609 22722 10305 22761
rect 10628 24775 10756 24813
rect 10628 24719 10664 24775
rect 10720 24719 10756 24775
rect 10628 24558 10756 24719
rect 10628 24502 10664 24558
rect 10720 24502 10756 24558
rect 10628 24340 10756 24502
rect 10628 24284 10664 24340
rect 10720 24284 10756 24340
rect 10628 24123 10756 24284
rect 10628 24067 10664 24123
rect 10720 24067 10756 24123
rect 10628 23905 10756 24067
rect 10628 23849 10664 23905
rect 10720 23849 10756 23905
rect 10628 23687 10756 23849
rect 10628 23631 10664 23687
rect 10720 23631 10756 23687
rect 10628 23469 10756 23631
rect 10628 23413 10664 23469
rect 10720 23413 10756 23469
rect 10628 23252 10756 23413
rect 10628 23196 10664 23252
rect 10720 23196 10756 23252
rect 10628 23034 10756 23196
rect 10628 22978 10664 23034
rect 10720 22978 10756 23034
rect 10628 22817 10756 22978
rect 10628 22761 10664 22817
rect 10720 22761 10756 22817
rect 10628 22722 10756 22761
rect 10950 24775 11078 24813
rect 10950 24719 10986 24775
rect 11042 24719 11078 24775
rect 10950 24558 11078 24719
rect 10950 24502 10986 24558
rect 11042 24502 11078 24558
rect 10950 24340 11078 24502
rect 10950 24284 10986 24340
rect 11042 24284 11078 24340
rect 10950 24123 11078 24284
rect 10950 24067 10986 24123
rect 11042 24067 11078 24123
rect 10950 23905 11078 24067
rect 10950 23849 10986 23905
rect 11042 23849 11078 23905
rect 10950 23687 11078 23849
rect 10950 23631 10986 23687
rect 11042 23631 11078 23687
rect 10950 23469 11078 23631
rect 10950 23413 10986 23469
rect 11042 23413 11078 23469
rect 10950 23252 11078 23413
rect 10950 23196 10986 23252
rect 11042 23196 11078 23252
rect 10950 23034 11078 23196
rect 10950 22978 10986 23034
rect 11042 22978 11078 23034
rect 10950 22817 11078 22978
rect 10950 22761 10986 22817
rect 11042 22761 11078 22817
rect 10950 22722 11078 22761
rect 11401 24775 12097 24841
rect 11401 24719 11438 24775
rect 11494 24719 11721 24775
rect 11777 24719 12004 24775
rect 12060 24719 12097 24775
rect 11401 24558 12097 24719
rect 11401 24502 11438 24558
rect 11494 24502 11721 24558
rect 11777 24502 12004 24558
rect 12060 24502 12097 24558
rect 11401 24340 12097 24502
rect 11401 24284 11438 24340
rect 11494 24284 11721 24340
rect 11777 24284 12004 24340
rect 12060 24284 12097 24340
rect 11401 24123 12097 24284
rect 11401 24067 11438 24123
rect 11494 24067 11721 24123
rect 11777 24067 12004 24123
rect 12060 24067 12097 24123
rect 11401 23905 12097 24067
rect 11401 23849 11438 23905
rect 11494 23849 11721 23905
rect 11777 23849 12004 23905
rect 12060 23849 12097 23905
rect 11401 23687 12097 23849
rect 11401 23631 11438 23687
rect 11494 23631 11721 23687
rect 11777 23631 12004 23687
rect 12060 23631 12097 23687
rect 11401 23469 12097 23631
rect 11401 23413 11438 23469
rect 11494 23413 11721 23469
rect 11777 23413 12004 23469
rect 12060 23413 12097 23469
rect 11401 23252 12097 23413
rect 11401 23196 11438 23252
rect 11494 23196 11721 23252
rect 11777 23196 12004 23252
rect 12060 23196 12097 23252
rect 11401 23034 12097 23196
rect 11401 22978 11438 23034
rect 11494 22978 11721 23034
rect 11777 22978 12004 23034
rect 12060 22978 12097 23034
rect 11401 22817 12097 22978
rect 11401 22761 11438 22817
rect 11494 22761 11721 22817
rect 11777 22761 12004 22817
rect 12060 22761 12097 22817
rect 11401 22722 12097 22761
rect 12420 24775 12548 24813
rect 12420 24719 12456 24775
rect 12512 24719 12548 24775
rect 12420 24558 12548 24719
rect 12420 24502 12456 24558
rect 12512 24502 12548 24558
rect 12420 24340 12548 24502
rect 12420 24284 12456 24340
rect 12512 24284 12548 24340
rect 12420 24123 12548 24284
rect 12420 24067 12456 24123
rect 12512 24067 12548 24123
rect 12420 23905 12548 24067
rect 12420 23849 12456 23905
rect 12512 23849 12548 23905
rect 12420 23687 12548 23849
rect 12420 23631 12456 23687
rect 12512 23631 12548 23687
rect 12420 23469 12548 23631
rect 12420 23413 12456 23469
rect 12512 23413 12548 23469
rect 12420 23252 12548 23413
rect 12420 23196 12456 23252
rect 12512 23196 12548 23252
rect 12420 23034 12548 23196
rect 12420 22978 12456 23034
rect 12512 22978 12548 23034
rect 12420 22817 12548 22978
rect 12420 22761 12456 22817
rect 12512 22761 12548 22817
rect 12420 22722 12548 22761
rect 8739 21987 8776 22043
rect 8832 21987 8868 22043
rect 8739 21825 8868 21987
rect 8739 21769 8776 21825
rect 8832 21769 8868 21825
rect 8739 19828 8868 21769
rect 9155 21842 9507 21882
rect 9155 21790 9418 21842
rect 9470 21790 9507 21842
rect 9155 21624 9507 21790
rect 9155 21572 9418 21624
rect 9470 21572 9507 21624
rect 9155 21531 9507 21572
rect 10407 21842 10759 21882
rect 10407 21790 10444 21842
rect 10496 21790 10759 21842
rect 10407 21624 10759 21790
rect 10407 21572 10444 21624
rect 10496 21572 10759 21624
rect 10407 21531 10759 21572
rect 9155 20502 9283 21531
rect 9155 20450 9193 20502
rect 9245 20450 9283 20502
rect 9155 20284 9283 20450
rect 9155 20232 9193 20284
rect 9245 20232 9283 20284
rect 9155 20196 9283 20232
rect 9609 20366 10305 20542
rect 9609 20310 9646 20366
rect 9702 20310 9929 20366
rect 9985 20310 10212 20366
rect 10268 20310 10305 20366
rect 9155 20067 9282 20196
rect 9155 20015 9193 20067
rect 9245 20015 9282 20067
rect 9155 19849 9282 20015
rect 9155 19797 9193 19849
rect 9245 19797 9282 19849
rect 9155 19631 9282 19797
rect 7617 19567 7653 19572
rect 7529 19527 7653 19567
rect 8249 19493 8868 19626
rect 9155 19579 9193 19631
rect 9245 19579 9282 19631
rect 5045 19361 5082 19413
rect 5134 19361 5172 19413
rect 5045 19196 5172 19361
rect 5045 19144 5082 19196
rect 5134 19144 5172 19196
rect 5045 18978 5172 19144
rect 5045 18926 5082 18978
rect 5134 18926 5172 18978
rect 5045 18886 5172 18926
rect 9155 19413 9282 19579
rect 9155 19361 9193 19413
rect 9245 19361 9282 19413
rect 9155 19196 9282 19361
rect 9155 19144 9193 19196
rect 9245 19144 9282 19196
rect 9155 18978 9282 19144
rect 9155 18926 9193 18978
rect 9245 18926 9282 18978
rect 9155 18886 9282 18926
rect 9609 20148 10305 20310
rect 10631 20502 10759 21531
rect 10631 20450 10669 20502
rect 10721 20450 10759 20502
rect 10631 20284 10759 20450
rect 10631 20232 10669 20284
rect 10721 20232 10759 20284
rect 10631 20196 10759 20232
rect 9609 20092 9646 20148
rect 9702 20092 9929 20148
rect 9985 20092 10212 20148
rect 10268 20092 10305 20148
rect 9609 19930 10305 20092
rect 9609 19874 9646 19930
rect 9702 19874 9929 19930
rect 9985 19874 10212 19930
rect 10268 19874 10305 19930
rect 9609 19711 10305 19874
rect 9609 19659 9648 19711
rect 9700 19659 9931 19711
rect 9983 19659 10214 19711
rect 10266 19659 10305 19711
rect 9609 19494 10305 19659
rect 9609 19442 9648 19494
rect 9700 19442 9931 19494
rect 9983 19442 10214 19494
rect 10266 19442 10305 19494
rect 9609 19276 10305 19442
rect 9609 19224 9648 19276
rect 9700 19224 9931 19276
rect 9983 19224 10214 19276
rect 10266 19224 10305 19276
rect 9609 19058 10305 19224
rect 9609 19006 9648 19058
rect 9700 19006 9931 19058
rect 9983 19006 10214 19058
rect 10266 19006 10305 19058
rect 4022 18788 4061 18840
rect 4113 18788 4344 18840
rect 4396 18788 4627 18840
rect 4679 18788 4718 18840
rect 4022 18623 4718 18788
rect 4022 18571 4061 18623
rect 4113 18571 4344 18623
rect 4396 18571 4627 18623
rect 4679 18571 4718 18623
rect 4022 18408 4718 18571
rect 4022 18352 4059 18408
rect 4115 18352 4342 18408
rect 4398 18352 4625 18408
rect 4681 18352 4718 18408
rect 4022 18190 4718 18352
rect 4022 18134 4059 18190
rect 4115 18134 4342 18190
rect 4398 18134 4625 18190
rect 4681 18134 4718 18190
rect 4022 17972 4718 18134
rect 4022 17916 4059 17972
rect 4115 17916 4342 17972
rect 4398 17916 4625 17972
rect 4681 17916 4718 17972
rect 9609 18840 10305 19006
rect 10632 20067 10759 20196
rect 10632 20015 10669 20067
rect 10721 20015 10759 20067
rect 10632 19849 10759 20015
rect 10632 19797 10669 19849
rect 10721 19797 10759 19849
rect 10632 19631 10759 19797
rect 10632 19579 10669 19631
rect 10721 19579 10759 19631
rect 10632 19413 10759 19579
rect 10632 19361 10669 19413
rect 10721 19361 10759 19413
rect 10632 19196 10759 19361
rect 10632 19144 10669 19196
rect 10721 19144 10759 19196
rect 10632 18978 10759 19144
rect 10632 18926 10669 18978
rect 10721 18926 10759 18978
rect 10632 18886 10759 18926
rect 10947 21842 11299 21882
rect 10947 21790 11210 21842
rect 11262 21790 11299 21842
rect 10947 21624 11299 21790
rect 10947 21572 11210 21624
rect 11262 21572 11299 21624
rect 10947 21531 11299 21572
rect 12199 21842 12551 21882
rect 12199 21790 12236 21842
rect 12288 21790 12551 21842
rect 12199 21624 12551 21790
rect 12199 21572 12236 21624
rect 12288 21572 12551 21624
rect 12199 21531 12551 21572
rect 10947 20502 11075 21531
rect 10947 20450 10985 20502
rect 11037 20450 11075 20502
rect 10947 20284 11075 20450
rect 10947 20232 10985 20284
rect 11037 20232 11075 20284
rect 10947 20196 11075 20232
rect 11401 20366 12097 20542
rect 11401 20310 11438 20366
rect 11494 20310 11721 20366
rect 11777 20310 12004 20366
rect 12060 20310 12097 20366
rect 10947 20067 11074 20196
rect 10947 20015 10985 20067
rect 11037 20015 11074 20067
rect 10947 19849 11074 20015
rect 10947 19797 10985 19849
rect 11037 19797 11074 19849
rect 10947 19631 11074 19797
rect 10947 19579 10985 19631
rect 11037 19579 11074 19631
rect 10947 19413 11074 19579
rect 10947 19361 10985 19413
rect 11037 19361 11074 19413
rect 10947 19196 11074 19361
rect 10947 19144 10985 19196
rect 11037 19144 11074 19196
rect 10947 18978 11074 19144
rect 10947 18926 10985 18978
rect 11037 18926 11074 18978
rect 10947 18886 11074 18926
rect 11401 20148 12097 20310
rect 12423 20502 12551 21531
rect 12423 20450 12461 20502
rect 12513 20450 12551 20502
rect 12423 20284 12551 20450
rect 12423 20232 12461 20284
rect 12513 20232 12551 20284
rect 12423 20196 12551 20232
rect 11401 20092 11438 20148
rect 11494 20092 11721 20148
rect 11777 20092 12004 20148
rect 12060 20092 12097 20148
rect 11401 19930 12097 20092
rect 11401 19874 11438 19930
rect 11494 19874 11721 19930
rect 11777 19874 12004 19930
rect 12060 19874 12097 19930
rect 11401 19711 12097 19874
rect 11401 19659 11440 19711
rect 11492 19659 11723 19711
rect 11775 19659 12006 19711
rect 12058 19659 12097 19711
rect 11401 19494 12097 19659
rect 11401 19442 11440 19494
rect 11492 19442 11723 19494
rect 11775 19442 12006 19494
rect 12058 19442 12097 19494
rect 11401 19276 12097 19442
rect 11401 19224 11440 19276
rect 11492 19224 11723 19276
rect 11775 19224 12006 19276
rect 12058 19224 12097 19276
rect 11401 19058 12097 19224
rect 11401 19006 11440 19058
rect 11492 19006 11723 19058
rect 11775 19006 12006 19058
rect 12058 19006 12097 19058
rect 9609 18788 9648 18840
rect 9700 18788 9931 18840
rect 9983 18788 10214 18840
rect 10266 18788 10305 18840
rect 9609 18623 10305 18788
rect 9609 18571 9648 18623
rect 9700 18571 9931 18623
rect 9983 18571 10214 18623
rect 10266 18571 10305 18623
rect 9609 18408 10305 18571
rect 9609 18352 9646 18408
rect 9702 18352 9929 18408
rect 9985 18352 10212 18408
rect 10268 18352 10305 18408
rect 9609 18190 10305 18352
rect 9609 18134 9646 18190
rect 9702 18134 9929 18190
rect 9985 18134 10212 18190
rect 10268 18134 10305 18190
rect 9609 17972 10305 18134
rect 4022 17754 4718 17916
rect 6842 17793 6971 17927
rect 8533 17793 8662 17927
rect 9609 17916 9646 17972
rect 9702 17916 9929 17972
rect 9985 17916 10212 17972
rect 10268 17916 10305 17972
rect 4022 17698 4059 17754
rect 4115 17698 4342 17754
rect 4398 17698 4625 17754
rect 4681 17698 4718 17754
rect 4022 17657 4718 17698
rect 9609 17754 10305 17916
rect 9609 17698 9646 17754
rect 9702 17698 9929 17754
rect 9985 17698 10212 17754
rect 10268 17698 10305 17754
rect 9609 17657 10305 17698
rect 11401 18840 12097 19006
rect 12424 20067 12551 20196
rect 12424 20015 12461 20067
rect 12513 20015 12551 20067
rect 12424 19849 12551 20015
rect 12424 19797 12461 19849
rect 12513 19797 12551 19849
rect 12424 19631 12551 19797
rect 12424 19579 12461 19631
rect 12513 19579 12551 19631
rect 12424 19413 12551 19579
rect 13215 19837 13344 25129
rect 13435 24804 13563 24842
rect 13435 24748 13471 24804
rect 13527 24748 13563 24804
rect 13435 24587 13563 24748
rect 13435 24531 13471 24587
rect 13527 24531 13563 24587
rect 13435 24369 13563 24531
rect 13435 24313 13471 24369
rect 13527 24313 13563 24369
rect 13435 24152 13563 24313
rect 13435 24096 13471 24152
rect 13527 24096 13563 24152
rect 13435 23934 13563 24096
rect 13435 23878 13471 23934
rect 13527 23878 13563 23934
rect 13435 23716 13563 23878
rect 13435 23660 13471 23716
rect 13527 23660 13563 23716
rect 13435 23498 13563 23660
rect 13435 23442 13471 23498
rect 13527 23442 13563 23498
rect 13435 23281 13563 23442
rect 13435 23225 13471 23281
rect 13527 23225 13563 23281
rect 13435 23063 13563 23225
rect 13949 24813 14077 24851
rect 13949 24757 13985 24813
rect 14041 24757 14077 24813
rect 13949 24595 14077 24757
rect 13949 24539 13985 24595
rect 14041 24539 14077 24595
rect 13949 24378 14077 24539
rect 13949 24322 13985 24378
rect 14041 24322 14077 24378
rect 13949 24160 14077 24322
rect 13949 24104 13985 24160
rect 14041 24104 14077 24160
rect 13949 23942 14077 24104
rect 13949 23886 13985 23942
rect 14041 23886 14077 23942
rect 13949 23724 14077 23886
rect 13949 23668 13985 23724
rect 14041 23668 14077 23724
rect 13949 23507 14077 23668
rect 13949 23451 13985 23507
rect 14041 23451 14077 23507
rect 13949 23289 14077 23451
rect 13949 23233 13985 23289
rect 14041 23233 14077 23289
rect 13949 23195 14077 23233
rect 13435 23007 13471 23063
rect 13527 23007 13563 23063
rect 14451 23054 14580 26881
rect 15477 26864 15605 26902
rect 16118 27425 16157 27477
rect 16209 27425 16247 27477
rect 14906 26516 15241 26554
rect 14906 26460 14942 26516
rect 14998 26460 15149 26516
rect 15205 26460 15241 26516
rect 14906 26298 15241 26460
rect 14906 26242 14942 26298
rect 14998 26242 15149 26298
rect 15205 26242 15241 26298
rect 14906 26080 15241 26242
rect 14906 26024 14942 26080
rect 14998 26024 15149 26080
rect 15205 26024 15241 26080
rect 14906 25862 15241 26024
rect 14906 25806 14942 25862
rect 14998 25806 15149 25862
rect 15205 25806 15241 25862
rect 14906 25768 15241 25806
rect 15633 26493 15761 26530
rect 15633 26437 15669 26493
rect 15725 26437 15761 26493
rect 15633 26275 15761 26437
rect 15633 26219 15669 26275
rect 15725 26219 15761 26275
rect 15633 26057 15761 26219
rect 15633 26001 15669 26057
rect 15725 26001 15761 26057
rect 15633 25839 15761 26001
rect 15633 25783 15669 25839
rect 15725 25783 15761 25839
rect 15633 25745 15761 25783
rect 13435 22846 13563 23007
rect 13435 22790 13471 22846
rect 13527 22790 13563 22846
rect 13435 22751 13563 22790
rect 13937 22921 14580 23054
rect 14906 25221 15246 25262
rect 14906 25169 14944 25221
rect 14996 25169 15156 25221
rect 15208 25169 15246 25221
rect 14906 25129 15246 25169
rect 13654 21796 13778 21836
rect 13654 21744 13690 21796
rect 13742 21744 13778 21796
rect 13654 21578 13778 21744
rect 13654 21526 13690 21578
rect 13742 21526 13778 21578
rect 13654 21486 13778 21526
rect 13937 21567 14066 22921
rect 13937 21511 13974 21567
rect 14030 21511 14066 21567
rect 13215 19785 13253 19837
rect 13305 19785 13344 19837
rect 13215 19619 13344 19785
rect 13215 19572 13253 19619
rect 13217 19567 13253 19572
rect 13305 19572 13344 19619
rect 13937 21349 14066 21511
rect 13937 21293 13974 21349
rect 14030 21293 14066 21349
rect 13937 19626 14066 21293
rect 14166 22703 14295 22744
rect 14166 22651 14204 22703
rect 14256 22651 14295 22703
rect 14166 22485 14295 22651
rect 14166 22433 14204 22485
rect 14256 22433 14295 22485
rect 14166 21162 14295 22433
rect 14429 22043 14554 22082
rect 14429 21987 14464 22043
rect 14520 21987 14554 22043
rect 14429 21866 14554 21987
rect 14166 21110 14204 21162
rect 14256 21110 14295 21162
rect 14166 21069 14295 21110
rect 14427 21825 14556 21866
rect 14427 21769 14464 21825
rect 14520 21769 14556 21825
rect 14427 19828 14556 21769
rect 14906 19837 15035 25129
rect 15126 24804 15254 24842
rect 15126 24748 15162 24804
rect 15218 24748 15254 24804
rect 15126 24587 15254 24748
rect 15126 24531 15162 24587
rect 15218 24531 15254 24587
rect 15126 24369 15254 24531
rect 15126 24313 15162 24369
rect 15218 24313 15254 24369
rect 15126 24152 15254 24313
rect 15126 24096 15162 24152
rect 15218 24096 15254 24152
rect 15126 23934 15254 24096
rect 15126 23878 15162 23934
rect 15218 23878 15254 23934
rect 15126 23716 15254 23878
rect 15126 23660 15162 23716
rect 15218 23660 15254 23716
rect 15126 23498 15254 23660
rect 15126 23442 15162 23498
rect 15218 23442 15254 23498
rect 15126 23281 15254 23442
rect 15126 23225 15162 23281
rect 15218 23225 15254 23281
rect 15126 23063 15254 23225
rect 15640 24813 15768 24851
rect 15640 24757 15676 24813
rect 15732 24757 15768 24813
rect 15640 24595 15768 24757
rect 15640 24539 15676 24595
rect 15732 24539 15768 24595
rect 15640 24378 15768 24539
rect 15640 24322 15676 24378
rect 15732 24322 15768 24378
rect 15640 24160 15768 24322
rect 15640 24104 15676 24160
rect 15732 24104 15768 24160
rect 15640 23942 15768 24104
rect 15640 23886 15676 23942
rect 15732 23886 15768 23942
rect 15640 23724 15768 23886
rect 15640 23668 15676 23724
rect 15732 23668 15768 23724
rect 15640 23507 15768 23668
rect 15640 23451 15676 23507
rect 15732 23451 15768 23507
rect 15640 23289 15768 23451
rect 15640 23233 15676 23289
rect 15732 23233 15768 23289
rect 15640 23195 15768 23233
rect 15126 23007 15162 23063
rect 15218 23007 15254 23063
rect 15126 22846 15254 23007
rect 15126 22790 15162 22846
rect 15218 22790 15254 22846
rect 15126 22751 15254 22790
rect 15857 22703 15986 22744
rect 15857 22651 15895 22703
rect 15947 22651 15986 22703
rect 15857 22485 15986 22651
rect 15857 22433 15895 22485
rect 15947 22433 15986 22485
rect 15343 21796 15472 21837
rect 15343 21744 15381 21796
rect 15433 21744 15472 21796
rect 15343 21578 15472 21744
rect 15630 21605 15755 21606
rect 15343 21526 15381 21578
rect 15433 21526 15472 21578
rect 15343 20960 15472 21526
rect 15343 20908 15381 20960
rect 15433 20908 15472 20960
rect 15343 20867 15472 20908
rect 15628 21567 15757 21605
rect 15628 21511 15665 21567
rect 15721 21511 15757 21567
rect 15628 21349 15757 21511
rect 15628 21293 15665 21349
rect 15721 21293 15757 21349
rect 14906 19785 14944 19837
rect 14996 19785 15035 19837
rect 13305 19567 13341 19572
rect 13217 19527 13341 19567
rect 13937 19493 14556 19626
rect 14906 19619 15035 19785
rect 14906 19572 14944 19619
rect 14908 19567 14944 19572
rect 14996 19572 15035 19619
rect 15628 19626 15757 21293
rect 15857 20758 15986 22433
rect 15857 20706 15895 20758
rect 15947 20706 15986 20758
rect 15857 20665 15986 20706
rect 16118 22043 16247 27425
rect 24936 27439 25061 27478
rect 23750 27380 23875 27419
rect 23750 27324 23785 27380
rect 23841 27324 23875 27380
rect 23750 27162 23875 27324
rect 23750 27106 23785 27162
rect 23841 27106 23875 27162
rect 24936 27383 24971 27439
rect 25027 27383 25061 27439
rect 26604 27468 26733 27545
rect 24936 27221 25061 27383
rect 24936 27165 24971 27221
rect 25027 27165 25061 27221
rect 24936 27127 25061 27165
rect 25964 27394 26089 27433
rect 25964 27338 25999 27394
rect 26055 27338 26089 27394
rect 25964 27176 26089 27338
rect 23750 27068 23875 27106
rect 25964 27120 25999 27176
rect 26055 27120 26089 27176
rect 25964 27082 26089 27120
rect 26604 27416 26642 27468
rect 26694 27416 26733 27468
rect 24832 26974 25171 27015
rect 24832 26922 24869 26974
rect 24921 26922 25081 26974
rect 25133 26922 25171 26974
rect 24832 26882 25171 26922
rect 23701 26537 24036 26575
rect 23701 26481 23737 26537
rect 23793 26481 23944 26537
rect 24000 26481 24036 26537
rect 23701 26319 24036 26481
rect 23701 26263 23737 26319
rect 23793 26263 23944 26319
rect 24000 26263 24036 26319
rect 23701 26101 24036 26263
rect 23701 26045 23737 26101
rect 23793 26045 23944 26101
rect 24000 26045 24036 26101
rect 23701 25883 24036 26045
rect 23701 25827 23737 25883
rect 23793 25827 23944 25883
rect 24000 25827 24036 25883
rect 23701 25788 24036 25827
rect 24428 26537 24556 26574
rect 24428 26481 24464 26537
rect 24520 26481 24556 26537
rect 24428 26319 24556 26481
rect 24428 26263 24464 26319
rect 24520 26263 24556 26319
rect 24428 26101 24556 26263
rect 24428 26045 24464 26101
rect 24520 26045 24556 26101
rect 24428 25883 24556 26045
rect 24428 25827 24464 25883
rect 24520 25827 24556 25883
rect 24428 25789 24556 25827
rect 16887 25302 17015 25339
rect 16887 25246 16923 25302
rect 16979 25246 17015 25302
rect 16887 25084 17015 25246
rect 16887 25028 16923 25084
rect 16979 25028 17015 25084
rect 16887 24866 17015 25028
rect 16887 24810 16923 24866
rect 16979 24810 17015 24866
rect 16887 24772 17015 24810
rect 17335 25302 17463 25339
rect 17335 25246 17371 25302
rect 17427 25246 17463 25302
rect 17335 25084 17463 25246
rect 17335 25028 17371 25084
rect 17427 25028 17463 25084
rect 17335 24866 17463 25028
rect 17335 24810 17371 24866
rect 17427 24810 17463 24866
rect 17335 24772 17463 24810
rect 17783 25302 17911 25339
rect 17783 25246 17819 25302
rect 17875 25246 17911 25302
rect 17783 25084 17911 25246
rect 17783 25028 17819 25084
rect 17875 25028 17911 25084
rect 17783 24866 17911 25028
rect 17783 24810 17819 24866
rect 17875 24810 17911 24866
rect 17783 24772 17911 24810
rect 18521 25302 18649 25339
rect 18521 25246 18557 25302
rect 18613 25246 18649 25302
rect 18521 25084 18649 25246
rect 18521 25028 18557 25084
rect 18613 25028 18649 25084
rect 18521 24866 18649 25028
rect 18521 24810 18557 24866
rect 18613 24810 18649 24866
rect 18521 24772 18649 24810
rect 18969 25302 19097 25339
rect 18969 25246 19005 25302
rect 19061 25246 19097 25302
rect 18969 25084 19097 25246
rect 18969 25028 19005 25084
rect 19061 25028 19097 25084
rect 18969 24866 19097 25028
rect 18969 24810 19005 24866
rect 19061 24810 19097 24866
rect 18969 24772 19097 24810
rect 19417 25302 19545 25339
rect 19417 25246 19453 25302
rect 19509 25246 19545 25302
rect 19417 25084 19545 25246
rect 19417 25028 19453 25084
rect 19509 25028 19545 25084
rect 19417 24866 19545 25028
rect 19417 24810 19453 24866
rect 19509 24810 19545 24866
rect 19417 24772 19545 24810
rect 20154 25302 20282 25339
rect 20154 25246 20190 25302
rect 20246 25246 20282 25302
rect 20154 25084 20282 25246
rect 20154 25028 20190 25084
rect 20246 25028 20282 25084
rect 20154 24866 20282 25028
rect 20154 24810 20190 24866
rect 20246 24810 20282 24866
rect 20154 24772 20282 24810
rect 20602 25302 20730 25339
rect 20602 25246 20638 25302
rect 20694 25246 20730 25302
rect 20602 25084 20730 25246
rect 20602 25028 20638 25084
rect 20694 25028 20730 25084
rect 20602 24866 20730 25028
rect 20602 24810 20638 24866
rect 20694 24810 20730 24866
rect 20602 24772 20730 24810
rect 21050 25302 21178 25339
rect 21050 25246 21086 25302
rect 21142 25246 21178 25302
rect 21050 25084 21178 25246
rect 21050 25028 21086 25084
rect 21142 25028 21178 25084
rect 21050 24866 21178 25028
rect 21050 24810 21086 24866
rect 21142 24810 21178 24866
rect 21050 24772 21178 24810
rect 21788 25302 21916 25339
rect 21788 25246 21824 25302
rect 21880 25246 21916 25302
rect 21788 25084 21916 25246
rect 21788 25028 21824 25084
rect 21880 25028 21916 25084
rect 21788 24866 21916 25028
rect 21788 24810 21824 24866
rect 21880 24810 21916 24866
rect 21788 24772 21916 24810
rect 22236 25302 22364 25339
rect 22236 25246 22272 25302
rect 22328 25246 22364 25302
rect 22236 25084 22364 25246
rect 22236 25028 22272 25084
rect 22328 25028 22364 25084
rect 22236 24866 22364 25028
rect 22236 24810 22272 24866
rect 22328 24810 22364 24866
rect 22236 24772 22364 24810
rect 22684 25302 22812 25339
rect 22684 25246 22720 25302
rect 22776 25246 22812 25302
rect 22684 25084 22812 25246
rect 22684 25028 22720 25084
rect 22776 25028 22812 25084
rect 22684 24866 22812 25028
rect 22684 24810 22720 24866
rect 22776 24810 22812 24866
rect 22684 24772 22812 24810
rect 23701 25312 24041 25353
rect 23701 25260 23739 25312
rect 23791 25260 23951 25312
rect 24003 25260 24041 25312
rect 23701 25220 24041 25260
rect 16891 24182 17019 24219
rect 16891 24126 16927 24182
rect 16983 24126 17019 24182
rect 16891 23964 17019 24126
rect 16891 23908 16927 23964
rect 16983 23908 17019 23964
rect 16891 23747 17019 23908
rect 16891 23691 16927 23747
rect 16983 23691 17019 23747
rect 16891 23529 17019 23691
rect 16891 23473 16927 23529
rect 16983 23473 17019 23529
rect 16891 23311 17019 23473
rect 16891 23255 16927 23311
rect 16983 23255 17019 23311
rect 16891 23094 17019 23255
rect 16891 23038 16927 23094
rect 16983 23038 17019 23094
rect 16891 22876 17019 23038
rect 16891 22820 16927 22876
rect 16983 22820 17019 22876
rect 16891 22782 17019 22820
rect 17335 24182 17463 24219
rect 17335 24126 17371 24182
rect 17427 24126 17463 24182
rect 17335 23964 17463 24126
rect 17335 23908 17371 23964
rect 17427 23908 17463 23964
rect 17335 23747 17463 23908
rect 17335 23691 17371 23747
rect 17427 23691 17463 23747
rect 17335 23529 17463 23691
rect 17335 23473 17371 23529
rect 17427 23473 17463 23529
rect 17335 23311 17463 23473
rect 17335 23255 17371 23311
rect 17427 23255 17463 23311
rect 17335 23094 17463 23255
rect 17335 23038 17371 23094
rect 17427 23038 17463 23094
rect 17335 22876 17463 23038
rect 17335 22820 17371 22876
rect 17427 22820 17463 22876
rect 17335 22782 17463 22820
rect 17779 24182 17907 24219
rect 17779 24126 17815 24182
rect 17871 24126 17907 24182
rect 17779 23964 17907 24126
rect 17779 23908 17815 23964
rect 17871 23908 17907 23964
rect 17779 23747 17907 23908
rect 17779 23691 17815 23747
rect 17871 23691 17907 23747
rect 17779 23529 17907 23691
rect 17779 23473 17815 23529
rect 17871 23473 17907 23529
rect 17779 23311 17907 23473
rect 17779 23255 17815 23311
rect 17871 23255 17907 23311
rect 17779 23094 17907 23255
rect 17779 23038 17815 23094
rect 17871 23038 17907 23094
rect 17779 22876 17907 23038
rect 17779 22820 17815 22876
rect 17871 22820 17907 22876
rect 17779 22782 17907 22820
rect 18525 24182 18653 24219
rect 18525 24126 18561 24182
rect 18617 24126 18653 24182
rect 18525 23964 18653 24126
rect 18525 23908 18561 23964
rect 18617 23908 18653 23964
rect 18525 23747 18653 23908
rect 18525 23691 18561 23747
rect 18617 23691 18653 23747
rect 18525 23529 18653 23691
rect 18525 23473 18561 23529
rect 18617 23473 18653 23529
rect 18525 23311 18653 23473
rect 18525 23255 18561 23311
rect 18617 23255 18653 23311
rect 18525 23094 18653 23255
rect 18525 23038 18561 23094
rect 18617 23038 18653 23094
rect 18525 22876 18653 23038
rect 18525 22820 18561 22876
rect 18617 22820 18653 22876
rect 18525 22782 18653 22820
rect 18969 24182 19097 24219
rect 18969 24126 19005 24182
rect 19061 24126 19097 24182
rect 18969 23964 19097 24126
rect 18969 23908 19005 23964
rect 19061 23908 19097 23964
rect 18969 23747 19097 23908
rect 18969 23691 19005 23747
rect 19061 23691 19097 23747
rect 18969 23529 19097 23691
rect 18969 23473 19005 23529
rect 19061 23473 19097 23529
rect 18969 23311 19097 23473
rect 18969 23255 19005 23311
rect 19061 23255 19097 23311
rect 18969 23094 19097 23255
rect 18969 23038 19005 23094
rect 19061 23038 19097 23094
rect 18969 22876 19097 23038
rect 18969 22820 19005 22876
rect 19061 22820 19097 22876
rect 18969 22782 19097 22820
rect 19413 24182 19541 24219
rect 19413 24126 19449 24182
rect 19505 24126 19541 24182
rect 19413 23964 19541 24126
rect 19413 23908 19449 23964
rect 19505 23908 19541 23964
rect 19413 23747 19541 23908
rect 19413 23691 19449 23747
rect 19505 23691 19541 23747
rect 19413 23529 19541 23691
rect 19413 23473 19449 23529
rect 19505 23473 19541 23529
rect 19413 23311 19541 23473
rect 19413 23255 19449 23311
rect 19505 23255 19541 23311
rect 19413 23094 19541 23255
rect 19413 23038 19449 23094
rect 19505 23038 19541 23094
rect 19413 22876 19541 23038
rect 19413 22820 19449 22876
rect 19505 22820 19541 22876
rect 19413 22782 19541 22820
rect 20158 24182 20286 24219
rect 20158 24126 20194 24182
rect 20250 24126 20286 24182
rect 20158 23964 20286 24126
rect 20158 23908 20194 23964
rect 20250 23908 20286 23964
rect 20158 23747 20286 23908
rect 20158 23691 20194 23747
rect 20250 23691 20286 23747
rect 20158 23529 20286 23691
rect 20158 23473 20194 23529
rect 20250 23473 20286 23529
rect 20158 23311 20286 23473
rect 20158 23255 20194 23311
rect 20250 23255 20286 23311
rect 20158 23094 20286 23255
rect 20158 23038 20194 23094
rect 20250 23038 20286 23094
rect 20158 22876 20286 23038
rect 20158 22820 20194 22876
rect 20250 22820 20286 22876
rect 20158 22782 20286 22820
rect 20602 24182 20730 24219
rect 20602 24126 20638 24182
rect 20694 24126 20730 24182
rect 20602 23964 20730 24126
rect 20602 23908 20638 23964
rect 20694 23908 20730 23964
rect 20602 23747 20730 23908
rect 20602 23691 20638 23747
rect 20694 23691 20730 23747
rect 20602 23529 20730 23691
rect 20602 23473 20638 23529
rect 20694 23473 20730 23529
rect 20602 23311 20730 23473
rect 20602 23255 20638 23311
rect 20694 23255 20730 23311
rect 20602 23094 20730 23255
rect 20602 23038 20638 23094
rect 20694 23038 20730 23094
rect 20602 22876 20730 23038
rect 20602 22820 20638 22876
rect 20694 22820 20730 22876
rect 20602 22782 20730 22820
rect 21046 24182 21174 24219
rect 21046 24126 21082 24182
rect 21138 24126 21174 24182
rect 21046 23964 21174 24126
rect 21046 23908 21082 23964
rect 21138 23908 21174 23964
rect 21046 23747 21174 23908
rect 21046 23691 21082 23747
rect 21138 23691 21174 23747
rect 21046 23529 21174 23691
rect 21046 23473 21082 23529
rect 21138 23473 21174 23529
rect 21046 23311 21174 23473
rect 21046 23255 21082 23311
rect 21138 23255 21174 23311
rect 21046 23094 21174 23255
rect 21046 23038 21082 23094
rect 21138 23038 21174 23094
rect 21046 22876 21174 23038
rect 21046 22820 21082 22876
rect 21138 22820 21174 22876
rect 21046 22782 21174 22820
rect 21792 24182 21920 24219
rect 21792 24126 21828 24182
rect 21884 24126 21920 24182
rect 21792 23964 21920 24126
rect 21792 23908 21828 23964
rect 21884 23908 21920 23964
rect 21792 23747 21920 23908
rect 21792 23691 21828 23747
rect 21884 23691 21920 23747
rect 21792 23529 21920 23691
rect 21792 23473 21828 23529
rect 21884 23473 21920 23529
rect 21792 23311 21920 23473
rect 21792 23255 21828 23311
rect 21884 23255 21920 23311
rect 21792 23094 21920 23255
rect 21792 23038 21828 23094
rect 21884 23038 21920 23094
rect 21792 22876 21920 23038
rect 21792 22820 21828 22876
rect 21884 22820 21920 22876
rect 21792 22782 21920 22820
rect 22236 24182 22364 24219
rect 22236 24126 22272 24182
rect 22328 24126 22364 24182
rect 22236 23964 22364 24126
rect 22236 23908 22272 23964
rect 22328 23908 22364 23964
rect 22236 23747 22364 23908
rect 22236 23691 22272 23747
rect 22328 23691 22364 23747
rect 22236 23529 22364 23691
rect 22236 23473 22272 23529
rect 22328 23473 22364 23529
rect 22236 23311 22364 23473
rect 22236 23255 22272 23311
rect 22328 23255 22364 23311
rect 22236 23094 22364 23255
rect 22236 23038 22272 23094
rect 22328 23038 22364 23094
rect 22236 22876 22364 23038
rect 22236 22820 22272 22876
rect 22328 22820 22364 22876
rect 22236 22782 22364 22820
rect 22680 24182 22808 24219
rect 22680 24126 22716 24182
rect 22772 24126 22808 24182
rect 22680 23964 22808 24126
rect 22680 23908 22716 23964
rect 22772 23908 22808 23964
rect 22680 23747 22808 23908
rect 22680 23691 22716 23747
rect 22772 23691 22808 23747
rect 22680 23529 22808 23691
rect 22680 23473 22716 23529
rect 22772 23473 22808 23529
rect 22680 23311 22808 23473
rect 22680 23255 22716 23311
rect 22772 23255 22808 23311
rect 22680 23094 22808 23255
rect 22680 23038 22716 23094
rect 22772 23038 22808 23094
rect 22680 22876 22808 23038
rect 22680 22820 22716 22876
rect 22772 22820 22808 22876
rect 22680 22782 22808 22820
rect 16118 21987 16155 22043
rect 16211 21987 16247 22043
rect 16118 21825 16247 21987
rect 16118 21769 16155 21825
rect 16211 21769 16247 21825
rect 16118 19828 16247 21769
rect 16663 22230 17239 22270
rect 16663 22178 16701 22230
rect 16753 22178 17149 22230
rect 17201 22178 17239 22230
rect 16663 22012 17239 22178
rect 16663 21960 16701 22012
rect 16753 21960 17149 22012
rect 17201 21960 17239 22012
rect 16663 21919 17239 21960
rect 17559 22230 18135 22270
rect 17559 22178 17597 22230
rect 17649 22178 18045 22230
rect 18097 22178 18135 22230
rect 17559 22012 18135 22178
rect 17559 21960 17597 22012
rect 17649 21960 18045 22012
rect 18097 21960 18135 22012
rect 17559 21919 18135 21960
rect 16663 20489 16791 21919
rect 16663 20437 16701 20489
rect 16753 20437 16791 20489
rect 16663 20271 16791 20437
rect 18007 20489 18135 21919
rect 18007 20437 18045 20489
rect 18097 20437 18135 20489
rect 16663 20219 16701 20271
rect 16753 20237 16791 20271
rect 17335 20387 17463 20424
rect 17335 20331 17371 20387
rect 17427 20331 17463 20387
rect 16753 20219 16790 20237
rect 16663 20054 16790 20219
rect 16663 20002 16701 20054
rect 16753 20002 16790 20054
rect 16663 19836 16790 20002
rect 16663 19784 16701 19836
rect 16753 19784 16790 19836
rect 14996 19567 15032 19572
rect 14908 19527 15032 19567
rect 15628 19493 16247 19626
rect 16663 19618 16790 19784
rect 16663 19566 16701 19618
rect 16753 19566 16790 19618
rect 12424 19361 12461 19413
rect 12513 19361 12551 19413
rect 12424 19196 12551 19361
rect 12424 19144 12461 19196
rect 12513 19144 12551 19196
rect 12424 18978 12551 19144
rect 12424 18926 12461 18978
rect 12513 18926 12551 18978
rect 12424 18886 12551 18926
rect 16663 19400 16790 19566
rect 16663 19348 16701 19400
rect 16753 19348 16790 19400
rect 16663 19183 16790 19348
rect 16663 19131 16701 19183
rect 16753 19131 16790 19183
rect 16663 18965 16790 19131
rect 16663 18913 16701 18965
rect 16753 18913 16790 18965
rect 16663 18873 16790 18913
rect 17335 20169 17463 20331
rect 18007 20271 18135 20437
rect 18007 20237 18045 20271
rect 17335 20113 17371 20169
rect 17427 20113 17463 20169
rect 17335 19951 17463 20113
rect 17335 19895 17371 19951
rect 17427 19895 17463 19951
rect 17335 19732 17463 19895
rect 17335 19680 17373 19732
rect 17425 19680 17463 19732
rect 17335 19514 17463 19680
rect 17335 19462 17373 19514
rect 17425 19462 17463 19514
rect 17335 19297 17463 19462
rect 17335 19245 17373 19297
rect 17425 19245 17463 19297
rect 17335 19079 17463 19245
rect 17335 19027 17373 19079
rect 17425 19027 17463 19079
rect 11401 18788 11440 18840
rect 11492 18788 11723 18840
rect 11775 18788 12006 18840
rect 12058 18788 12097 18840
rect 11401 18623 12097 18788
rect 11401 18571 11440 18623
rect 11492 18571 11723 18623
rect 11775 18571 12006 18623
rect 12058 18571 12097 18623
rect 11401 18408 12097 18571
rect 11401 18352 11438 18408
rect 11494 18352 11721 18408
rect 11777 18352 12004 18408
rect 12060 18352 12097 18408
rect 11401 18190 12097 18352
rect 11401 18134 11438 18190
rect 11494 18134 11721 18190
rect 11777 18134 12004 18190
rect 12060 18134 12097 18190
rect 11401 17972 12097 18134
rect 11401 17916 11438 17972
rect 11494 17916 11721 17972
rect 11777 17916 12004 17972
rect 12060 17916 12097 17972
rect 17335 18861 17463 19027
rect 18008 20219 18045 20237
rect 18097 20219 18135 20271
rect 18008 20054 18135 20219
rect 18008 20002 18045 20054
rect 18097 20002 18135 20054
rect 18008 19836 18135 20002
rect 18008 19784 18045 19836
rect 18097 19784 18135 19836
rect 18008 19618 18135 19784
rect 18008 19566 18045 19618
rect 18097 19566 18135 19618
rect 18008 19400 18135 19566
rect 18008 19348 18045 19400
rect 18097 19348 18135 19400
rect 18008 19183 18135 19348
rect 18008 19131 18045 19183
rect 18097 19131 18135 19183
rect 18008 18965 18135 19131
rect 18008 18913 18045 18965
rect 18097 18913 18135 18965
rect 18008 18873 18135 18913
rect 18297 22230 18873 22270
rect 18297 22178 18335 22230
rect 18387 22178 18783 22230
rect 18835 22178 18873 22230
rect 18297 22012 18873 22178
rect 18297 21960 18335 22012
rect 18387 21960 18783 22012
rect 18835 21960 18873 22012
rect 18297 21919 18873 21960
rect 19193 22230 19769 22270
rect 19193 22178 19231 22230
rect 19283 22178 19679 22230
rect 19731 22178 19769 22230
rect 19193 22012 19769 22178
rect 19193 21960 19231 22012
rect 19283 21960 19679 22012
rect 19731 21960 19769 22012
rect 19193 21919 19769 21960
rect 18297 20489 18425 21919
rect 18297 20437 18335 20489
rect 18387 20437 18425 20489
rect 18297 20271 18425 20437
rect 19641 20489 19769 21919
rect 19641 20437 19679 20489
rect 19731 20437 19769 20489
rect 18297 20219 18335 20271
rect 18387 20237 18425 20271
rect 18969 20387 19097 20424
rect 18969 20331 19005 20387
rect 19061 20331 19097 20387
rect 18387 20219 18424 20237
rect 18297 20054 18424 20219
rect 18297 20002 18335 20054
rect 18387 20002 18424 20054
rect 18297 19836 18424 20002
rect 18297 19784 18335 19836
rect 18387 19784 18424 19836
rect 18297 19618 18424 19784
rect 18297 19566 18335 19618
rect 18387 19566 18424 19618
rect 18297 19400 18424 19566
rect 18297 19348 18335 19400
rect 18387 19348 18424 19400
rect 18297 19183 18424 19348
rect 18297 19131 18335 19183
rect 18387 19131 18424 19183
rect 18297 18965 18424 19131
rect 18297 18913 18335 18965
rect 18387 18913 18424 18965
rect 18297 18873 18424 18913
rect 18969 20169 19097 20331
rect 19641 20271 19769 20437
rect 19641 20237 19679 20271
rect 18969 20113 19005 20169
rect 19061 20113 19097 20169
rect 18969 19951 19097 20113
rect 18969 19895 19005 19951
rect 19061 19895 19097 19951
rect 18969 19732 19097 19895
rect 18969 19680 19007 19732
rect 19059 19680 19097 19732
rect 18969 19514 19097 19680
rect 18969 19462 19007 19514
rect 19059 19462 19097 19514
rect 18969 19297 19097 19462
rect 18969 19245 19007 19297
rect 19059 19245 19097 19297
rect 18969 19079 19097 19245
rect 18969 19027 19007 19079
rect 19059 19027 19097 19079
rect 17335 18809 17373 18861
rect 17425 18809 17463 18861
rect 17335 18644 17463 18809
rect 17335 18592 17373 18644
rect 17425 18592 17463 18644
rect 17335 18428 17463 18592
rect 17335 18372 17371 18428
rect 17427 18372 17463 18428
rect 17335 18210 17463 18372
rect 17335 18154 17371 18210
rect 17427 18154 17463 18210
rect 17335 17992 17463 18154
rect 17335 17936 17371 17992
rect 17427 17936 17463 17992
rect 11401 17754 12097 17916
rect 14220 17793 14350 17927
rect 15911 17793 16041 17927
rect 11401 17698 11438 17754
rect 11494 17698 11721 17754
rect 11777 17698 12004 17754
rect 12060 17698 12097 17754
rect 11401 17657 12097 17698
rect 17335 17774 17463 17936
rect 17335 17718 17371 17774
rect 17427 17718 17463 17774
rect 17335 17680 17463 17718
rect 18969 18861 19097 19027
rect 19642 20219 19679 20237
rect 19731 20219 19769 20271
rect 19642 20054 19769 20219
rect 19642 20002 19679 20054
rect 19731 20002 19769 20054
rect 19642 19836 19769 20002
rect 19642 19784 19679 19836
rect 19731 19784 19769 19836
rect 19642 19618 19769 19784
rect 19642 19566 19679 19618
rect 19731 19566 19769 19618
rect 19642 19400 19769 19566
rect 19642 19348 19679 19400
rect 19731 19348 19769 19400
rect 19642 19183 19769 19348
rect 19642 19131 19679 19183
rect 19731 19131 19769 19183
rect 19642 18965 19769 19131
rect 19642 18913 19679 18965
rect 19731 18913 19769 18965
rect 19642 18873 19769 18913
rect 19930 22230 20506 22270
rect 19930 22178 19968 22230
rect 20020 22178 20416 22230
rect 20468 22178 20506 22230
rect 19930 22012 20506 22178
rect 19930 21960 19968 22012
rect 20020 21960 20416 22012
rect 20468 21960 20506 22012
rect 19930 21919 20506 21960
rect 20826 22230 21402 22270
rect 20826 22178 20864 22230
rect 20916 22178 21312 22230
rect 21364 22178 21402 22230
rect 20826 22012 21402 22178
rect 20826 21960 20864 22012
rect 20916 21960 21312 22012
rect 21364 21960 21402 22012
rect 20826 21919 21402 21960
rect 19930 20489 20058 21919
rect 19930 20437 19968 20489
rect 20020 20437 20058 20489
rect 19930 20271 20058 20437
rect 21274 20489 21402 21919
rect 21274 20437 21312 20489
rect 21364 20437 21402 20489
rect 19930 20219 19968 20271
rect 20020 20237 20058 20271
rect 20602 20387 20730 20424
rect 20602 20331 20638 20387
rect 20694 20331 20730 20387
rect 20020 20219 20057 20237
rect 19930 20054 20057 20219
rect 19930 20002 19968 20054
rect 20020 20002 20057 20054
rect 19930 19836 20057 20002
rect 19930 19784 19968 19836
rect 20020 19784 20057 19836
rect 19930 19618 20057 19784
rect 19930 19566 19968 19618
rect 20020 19566 20057 19618
rect 19930 19400 20057 19566
rect 19930 19348 19968 19400
rect 20020 19348 20057 19400
rect 19930 19183 20057 19348
rect 19930 19131 19968 19183
rect 20020 19131 20057 19183
rect 19930 18965 20057 19131
rect 19930 18913 19968 18965
rect 20020 18913 20057 18965
rect 19930 18873 20057 18913
rect 20602 20169 20730 20331
rect 21274 20271 21402 20437
rect 21274 20237 21312 20271
rect 20602 20113 20638 20169
rect 20694 20113 20730 20169
rect 20602 19951 20730 20113
rect 20602 19895 20638 19951
rect 20694 19895 20730 19951
rect 20602 19732 20730 19895
rect 20602 19680 20640 19732
rect 20692 19680 20730 19732
rect 20602 19514 20730 19680
rect 20602 19462 20640 19514
rect 20692 19462 20730 19514
rect 20602 19297 20730 19462
rect 20602 19245 20640 19297
rect 20692 19245 20730 19297
rect 20602 19079 20730 19245
rect 20602 19027 20640 19079
rect 20692 19027 20730 19079
rect 18969 18809 19007 18861
rect 19059 18809 19097 18861
rect 18969 18644 19097 18809
rect 18969 18592 19007 18644
rect 19059 18592 19097 18644
rect 18969 18428 19097 18592
rect 18969 18372 19005 18428
rect 19061 18372 19097 18428
rect 18969 18210 19097 18372
rect 18969 18154 19005 18210
rect 19061 18154 19097 18210
rect 18969 17992 19097 18154
rect 18969 17936 19005 17992
rect 19061 17936 19097 17992
rect 18969 17774 19097 17936
rect 18969 17718 19005 17774
rect 19061 17718 19097 17774
rect 18969 17680 19097 17718
rect 20602 18861 20730 19027
rect 21275 20219 21312 20237
rect 21364 20219 21402 20271
rect 21275 20054 21402 20219
rect 21275 20002 21312 20054
rect 21364 20002 21402 20054
rect 21275 19836 21402 20002
rect 21275 19784 21312 19836
rect 21364 19784 21402 19836
rect 21275 19618 21402 19784
rect 21275 19566 21312 19618
rect 21364 19566 21402 19618
rect 21275 19400 21402 19566
rect 21275 19348 21312 19400
rect 21364 19348 21402 19400
rect 21275 19183 21402 19348
rect 21275 19131 21312 19183
rect 21364 19131 21402 19183
rect 21275 18965 21402 19131
rect 21275 18913 21312 18965
rect 21364 18913 21402 18965
rect 21275 18873 21402 18913
rect 21564 22230 22140 22270
rect 21564 22178 21602 22230
rect 21654 22178 22050 22230
rect 22102 22178 22140 22230
rect 21564 22012 22140 22178
rect 21564 21960 21602 22012
rect 21654 21960 22050 22012
rect 22102 21960 22140 22012
rect 21564 21919 22140 21960
rect 22460 22230 23036 22270
rect 22460 22178 22498 22230
rect 22550 22178 22946 22230
rect 22998 22178 23036 22230
rect 22460 22012 23036 22178
rect 22460 21960 22498 22012
rect 22550 21960 22946 22012
rect 22998 21960 23036 22012
rect 22460 21919 23036 21960
rect 21564 20489 21692 21919
rect 21564 20437 21602 20489
rect 21654 20437 21692 20489
rect 21564 20271 21692 20437
rect 22908 20489 23036 21919
rect 22908 20437 22946 20489
rect 22998 20437 23036 20489
rect 21564 20219 21602 20271
rect 21654 20237 21692 20271
rect 22236 20387 22364 20424
rect 22236 20331 22272 20387
rect 22328 20331 22364 20387
rect 21654 20219 21691 20237
rect 21564 20054 21691 20219
rect 21564 20002 21602 20054
rect 21654 20002 21691 20054
rect 21564 19836 21691 20002
rect 21564 19784 21602 19836
rect 21654 19784 21691 19836
rect 21564 19618 21691 19784
rect 21564 19566 21602 19618
rect 21654 19566 21691 19618
rect 21564 19400 21691 19566
rect 21564 19348 21602 19400
rect 21654 19348 21691 19400
rect 21564 19183 21691 19348
rect 21564 19131 21602 19183
rect 21654 19131 21691 19183
rect 21564 18965 21691 19131
rect 21564 18913 21602 18965
rect 21654 18913 21691 18965
rect 21564 18873 21691 18913
rect 22236 20169 22364 20331
rect 22908 20271 23036 20437
rect 22908 20237 22946 20271
rect 22236 20113 22272 20169
rect 22328 20113 22364 20169
rect 22236 19951 22364 20113
rect 22236 19895 22272 19951
rect 22328 19895 22364 19951
rect 22236 19732 22364 19895
rect 22236 19680 22274 19732
rect 22326 19680 22364 19732
rect 22236 19514 22364 19680
rect 22236 19462 22274 19514
rect 22326 19462 22364 19514
rect 22236 19297 22364 19462
rect 22236 19245 22274 19297
rect 22326 19245 22364 19297
rect 22236 19079 22364 19245
rect 22236 19027 22274 19079
rect 22326 19027 22364 19079
rect 20602 18809 20640 18861
rect 20692 18809 20730 18861
rect 20602 18644 20730 18809
rect 20602 18592 20640 18644
rect 20692 18592 20730 18644
rect 20602 18428 20730 18592
rect 20602 18372 20638 18428
rect 20694 18372 20730 18428
rect 20602 18210 20730 18372
rect 20602 18154 20638 18210
rect 20694 18154 20730 18210
rect 20602 17992 20730 18154
rect 20602 17936 20638 17992
rect 20694 17936 20730 17992
rect 20602 17774 20730 17936
rect 20602 17718 20638 17774
rect 20694 17718 20730 17774
rect 20602 17680 20730 17718
rect 22236 18861 22364 19027
rect 22909 20219 22946 20237
rect 22998 20219 23036 20271
rect 22909 20054 23036 20219
rect 22909 20002 22946 20054
rect 22998 20002 23036 20054
rect 22909 19836 23036 20002
rect 22909 19784 22946 19836
rect 22998 19784 23036 19836
rect 22909 19618 23036 19784
rect 22909 19566 22946 19618
rect 22998 19566 23036 19618
rect 23701 19837 23830 25220
rect 23921 24999 24049 25038
rect 23921 24943 23957 24999
rect 24013 24943 24049 24999
rect 23921 24782 24049 24943
rect 23921 24726 23957 24782
rect 24013 24726 24049 24782
rect 23921 24564 24049 24726
rect 23921 24508 23957 24564
rect 24013 24508 24049 24564
rect 23921 24346 24049 24508
rect 23921 24290 23957 24346
rect 24013 24290 24049 24346
rect 23921 24128 24049 24290
rect 23921 24072 23957 24128
rect 24013 24072 24049 24128
rect 23921 23911 24049 24072
rect 23921 23855 23957 23911
rect 24013 23855 24049 23911
rect 23921 23816 24049 23855
rect 24435 24999 24563 25038
rect 24435 24943 24471 24999
rect 24527 24943 24563 24999
rect 24435 24782 24563 24943
rect 24435 24726 24471 24782
rect 24527 24726 24563 24782
rect 24435 24564 24563 24726
rect 24435 24508 24471 24564
rect 24527 24508 24563 24564
rect 24435 24346 24563 24508
rect 24435 24290 24471 24346
rect 24527 24290 24563 24346
rect 24435 24128 24563 24290
rect 24435 24072 24471 24128
rect 24527 24072 24563 24128
rect 24435 23911 24563 24072
rect 24435 23855 24471 23911
rect 24527 23855 24563 23911
rect 24435 23816 24563 23855
rect 24937 23270 25066 26882
rect 25391 26537 25726 26575
rect 25391 26481 25427 26537
rect 25483 26481 25634 26537
rect 25690 26481 25726 26537
rect 25391 26319 25726 26481
rect 25391 26263 25427 26319
rect 25483 26263 25634 26319
rect 25690 26263 25726 26319
rect 25391 26101 25726 26263
rect 25391 26045 25427 26101
rect 25483 26045 25634 26101
rect 25690 26045 25726 26101
rect 25391 25883 25726 26045
rect 25391 25827 25427 25883
rect 25483 25827 25634 25883
rect 25690 25827 25726 25883
rect 25391 25788 25726 25827
rect 26118 26537 26246 26574
rect 26118 26481 26154 26537
rect 26210 26481 26246 26537
rect 26118 26319 26246 26481
rect 26118 26263 26154 26319
rect 26210 26263 26246 26319
rect 26118 26101 26246 26263
rect 26118 26045 26154 26101
rect 26210 26045 26246 26101
rect 26118 25883 26246 26045
rect 26118 25827 26154 25883
rect 26210 25827 26246 25883
rect 26118 25789 26246 25827
rect 24423 23136 25066 23270
rect 25391 25312 25731 25353
rect 25391 25260 25429 25312
rect 25481 25260 25641 25312
rect 25693 25260 25731 25312
rect 25391 25220 25731 25260
rect 24140 22200 24264 22240
rect 24140 22148 24176 22200
rect 24228 22148 24264 22200
rect 24140 21982 24264 22148
rect 24140 21930 24176 21982
rect 24228 21930 24264 21982
rect 24140 21890 24264 21930
rect 24423 21970 24552 23136
rect 24915 22446 25040 22485
rect 24915 22390 24950 22446
rect 25006 22390 25040 22446
rect 24915 22270 25040 22390
rect 24423 21914 24460 21970
rect 24516 21914 24552 21970
rect 24423 21752 24552 21914
rect 24423 21696 24460 21752
rect 24516 21696 24552 21752
rect 24423 21658 24552 21696
rect 23701 19785 23739 19837
rect 23791 19785 23830 19837
rect 23701 19619 23830 19785
rect 23701 19572 23739 19619
rect 22909 19400 23036 19566
rect 23703 19567 23739 19572
rect 23791 19572 23830 19619
rect 24424 19626 24552 21658
rect 24651 22200 24780 22240
rect 24651 22148 24690 22200
rect 24742 22148 24780 22200
rect 24651 21982 24780 22148
rect 24651 21930 24690 21982
rect 24742 21930 24780 21982
rect 24651 21162 24780 21930
rect 24651 21110 24690 21162
rect 24742 21110 24780 21162
rect 24651 21069 24780 21110
rect 24914 22228 25042 22270
rect 24914 22172 24950 22228
rect 25006 22172 25042 22228
rect 24914 19828 25042 22172
rect 25391 19837 25520 25220
rect 25611 24999 25739 25038
rect 25611 24943 25647 24999
rect 25703 24943 25739 24999
rect 25611 24782 25739 24943
rect 25611 24726 25647 24782
rect 25703 24726 25739 24782
rect 25611 24564 25739 24726
rect 25611 24508 25647 24564
rect 25703 24508 25739 24564
rect 25611 24346 25739 24508
rect 25611 24290 25647 24346
rect 25703 24290 25739 24346
rect 25611 24128 25739 24290
rect 25611 24072 25647 24128
rect 25703 24072 25739 24128
rect 25611 23911 25739 24072
rect 25611 23855 25647 23911
rect 25703 23855 25739 23911
rect 25611 23816 25739 23855
rect 26125 24999 26253 25038
rect 26125 24943 26161 24999
rect 26217 24943 26253 24999
rect 26125 24782 26253 24943
rect 26125 24726 26161 24782
rect 26217 24726 26253 24782
rect 26125 24564 26253 24726
rect 26125 24508 26161 24564
rect 26217 24508 26253 24564
rect 26125 24346 26253 24508
rect 26125 24290 26161 24346
rect 26217 24290 26253 24346
rect 26125 24128 26253 24290
rect 26125 24072 26161 24128
rect 26217 24072 26253 24128
rect 26125 23911 26253 24072
rect 26125 23855 26161 23911
rect 26217 23855 26253 23911
rect 26125 23816 26253 23855
rect 26604 22446 26733 27416
rect 27082 26537 27417 26575
rect 27082 26481 27118 26537
rect 27174 26481 27325 26537
rect 27381 26481 27417 26537
rect 27082 26319 27417 26481
rect 27082 26263 27118 26319
rect 27174 26263 27325 26319
rect 27381 26263 27417 26319
rect 27082 26101 27417 26263
rect 27082 26045 27118 26101
rect 27174 26045 27325 26101
rect 27381 26045 27417 26101
rect 27082 25883 27417 26045
rect 27082 25827 27118 25883
rect 27174 25827 27325 25883
rect 27381 25827 27417 25883
rect 27082 25788 27417 25827
rect 27809 26537 27937 26574
rect 27809 26481 27845 26537
rect 27901 26481 27937 26537
rect 27809 26319 27937 26481
rect 27809 26263 27845 26319
rect 27901 26263 27937 26319
rect 27809 26101 27937 26263
rect 27809 26045 27845 26101
rect 27901 26045 27937 26101
rect 27809 25883 27937 26045
rect 27809 25827 27845 25883
rect 27901 25827 27937 25883
rect 27809 25789 27937 25827
rect 26604 22390 26640 22446
rect 26696 22390 26733 22446
rect 25828 22200 25957 22240
rect 25828 22148 25866 22200
rect 25918 22148 25957 22200
rect 25828 21982 25957 22148
rect 26342 22200 26471 22240
rect 26342 22148 26380 22200
rect 26432 22148 26471 22200
rect 25828 21930 25866 21982
rect 25918 21930 25957 21982
rect 25828 21565 25957 21930
rect 25828 21513 25867 21565
rect 25919 21513 25957 21565
rect 25828 21472 25957 21513
rect 26114 21970 26242 22009
rect 26114 21914 26150 21970
rect 26206 21914 26242 21970
rect 26114 21752 26242 21914
rect 26114 21696 26150 21752
rect 26206 21696 26242 21752
rect 25391 19785 25429 19837
rect 25481 19785 25520 19837
rect 23791 19567 23827 19572
rect 23703 19527 23827 19567
rect 24424 19493 25042 19626
rect 25391 19619 25520 19785
rect 25391 19572 25429 19619
rect 25393 19567 25429 19572
rect 25481 19572 25520 19619
rect 26114 19626 26242 21696
rect 26342 21982 26471 22148
rect 26342 21930 26380 21982
rect 26432 21930 26471 21982
rect 26342 20960 26471 21930
rect 26342 20908 26381 20960
rect 26433 20908 26471 20960
rect 26342 20867 26471 20908
rect 26604 22228 26733 22390
rect 26604 22172 26640 22228
rect 26696 22172 26733 22228
rect 26604 22134 26733 22172
rect 27082 25312 27422 25353
rect 27082 25260 27120 25312
rect 27172 25260 27332 25312
rect 27384 25260 27422 25312
rect 27082 25220 27422 25260
rect 26604 19828 26732 22134
rect 27082 19837 27211 25220
rect 27302 24999 27430 25038
rect 27302 24943 27338 24999
rect 27394 24943 27430 24999
rect 27302 24782 27430 24943
rect 27302 24726 27338 24782
rect 27394 24726 27430 24782
rect 27302 24564 27430 24726
rect 27302 24508 27338 24564
rect 27394 24508 27430 24564
rect 27302 24346 27430 24508
rect 27302 24290 27338 24346
rect 27394 24290 27430 24346
rect 27302 24128 27430 24290
rect 27302 24072 27338 24128
rect 27394 24072 27430 24128
rect 27302 23911 27430 24072
rect 27302 23855 27338 23911
rect 27394 23855 27430 23911
rect 27302 23816 27430 23855
rect 27816 24999 27944 25038
rect 27816 24943 27852 24999
rect 27908 24943 27944 24999
rect 27816 24782 27944 24943
rect 27816 24726 27852 24782
rect 27908 24726 27944 24782
rect 27816 24564 27944 24726
rect 27816 24508 27852 24564
rect 27908 24508 27944 24564
rect 27816 24346 27944 24508
rect 27816 24290 27852 24346
rect 27908 24290 27944 24346
rect 27816 24128 27944 24290
rect 27816 24072 27852 24128
rect 27908 24072 27944 24128
rect 27816 23911 27944 24072
rect 27816 23855 27852 23911
rect 27908 23855 27944 23911
rect 27816 23816 27944 23855
rect 28296 22446 28421 22485
rect 28296 22390 28331 22446
rect 28387 22390 28421 22446
rect 28296 22270 28421 22390
rect 27519 22200 27648 22240
rect 27519 22148 27557 22200
rect 27609 22148 27648 22200
rect 27519 21982 27648 22148
rect 28035 22200 28159 22240
rect 28035 22148 28071 22200
rect 28123 22148 28159 22200
rect 28035 22009 28159 22148
rect 28295 22228 28423 22270
rect 28295 22172 28331 22228
rect 28387 22172 28423 22228
rect 27519 21930 27557 21982
rect 27609 21930 27648 21982
rect 27519 21363 27648 21930
rect 27519 21311 27558 21363
rect 27610 21311 27648 21363
rect 27519 21270 27648 21311
rect 27805 21970 27933 22009
rect 27805 21914 27841 21970
rect 27897 21914 27933 21970
rect 27805 21752 27933 21914
rect 27805 21696 27841 21752
rect 27897 21696 27933 21752
rect 27082 19785 27120 19837
rect 27172 19785 27211 19837
rect 25481 19567 25517 19572
rect 25393 19527 25517 19567
rect 26114 19493 26732 19626
rect 27082 19619 27211 19785
rect 27082 19572 27120 19619
rect 27084 19567 27120 19572
rect 27172 19572 27211 19619
rect 27805 19626 27933 21696
rect 28033 21982 28162 22009
rect 28033 21930 28071 21982
rect 28123 21930 28162 21982
rect 28033 20758 28162 21930
rect 28033 20706 28072 20758
rect 28124 20706 28162 20758
rect 28033 20665 28162 20706
rect 28295 19828 28423 22172
rect 27172 19567 27208 19572
rect 27084 19527 27208 19567
rect 27805 19493 28423 19626
rect 22909 19348 22946 19400
rect 22998 19348 23036 19400
rect 22909 19183 23036 19348
rect 22909 19131 22946 19183
rect 22998 19131 23036 19183
rect 22909 18965 23036 19131
rect 22909 18913 22946 18965
rect 22998 18913 23036 18965
rect 22909 18873 23036 18913
rect 22236 18809 22274 18861
rect 22326 18809 22364 18861
rect 22236 18644 22364 18809
rect 22236 18592 22274 18644
rect 22326 18592 22364 18644
rect 22236 18428 22364 18592
rect 22236 18372 22272 18428
rect 22328 18372 22364 18428
rect 22236 18210 22364 18372
rect 22236 18154 22272 18210
rect 22328 18154 22364 18210
rect 22236 17992 22364 18154
rect 22236 17936 22272 17992
rect 22328 17936 22364 17992
rect 22236 17774 22364 17936
rect 24706 17793 24835 17927
rect 26397 17793 26526 17927
rect 28088 17793 28217 17927
rect 22236 17718 22272 17774
rect 22328 17718 22364 17774
rect 22236 17680 22364 17718
rect 1980 16904 2056 16914
rect 1980 16848 1990 16904
rect 2046 16848 2056 16904
rect 1980 16780 2056 16848
rect 1980 16724 1990 16780
rect 2046 16724 2056 16780
rect 1980 16656 2056 16724
rect 1980 16600 1990 16656
rect 2046 16600 2056 16656
rect 1980 16532 2056 16600
rect 1980 16476 1990 16532
rect 2046 16476 2056 16532
rect 1980 16408 2056 16476
rect 1980 16352 1990 16408
rect 2046 16352 2056 16408
rect 1980 16284 2056 16352
rect 1980 16228 1990 16284
rect 2046 16228 2056 16284
rect 1980 16160 2056 16228
rect 1980 16104 1990 16160
rect 2046 16104 2056 16160
rect 1980 16036 2056 16104
rect 1980 15980 1990 16036
rect 2046 15980 2056 16036
rect 1980 15912 2056 15980
rect 1980 15856 1990 15912
rect 2046 15856 2056 15912
rect 1980 15788 2056 15856
rect 1980 15732 1990 15788
rect 2046 15732 2056 15788
rect 1980 15664 2056 15732
rect 1980 15608 1990 15664
rect 2046 15608 2056 15664
rect 1980 15540 2056 15608
rect 1980 15484 1990 15540
rect 2046 15484 2056 15540
rect 1980 15474 2056 15484
rect 2652 16904 2728 16914
rect 2652 16848 2662 16904
rect 2718 16848 2728 16904
rect 2652 16780 2728 16848
rect 2652 16724 2662 16780
rect 2718 16724 2728 16780
rect 2652 16656 2728 16724
rect 2652 16600 2662 16656
rect 2718 16600 2728 16656
rect 2652 16532 2728 16600
rect 2652 16476 2662 16532
rect 2718 16476 2728 16532
rect 2652 16408 2728 16476
rect 2652 16352 2662 16408
rect 2718 16352 2728 16408
rect 2652 16284 2728 16352
rect 2652 16228 2662 16284
rect 2718 16228 2728 16284
rect 2652 16160 2728 16228
rect 2652 16104 2662 16160
rect 2718 16104 2728 16160
rect 2652 16036 2728 16104
rect 2652 15980 2662 16036
rect 2718 15980 2728 16036
rect 2652 15912 2728 15980
rect 2652 15856 2662 15912
rect 2718 15856 2728 15912
rect 2652 15788 2728 15856
rect 2652 15732 2662 15788
rect 2718 15732 2728 15788
rect 2652 15664 2728 15732
rect 2652 15608 2662 15664
rect 2718 15608 2728 15664
rect 2652 15540 2728 15608
rect 2652 15484 2662 15540
rect 2718 15484 2728 15540
rect 2652 15474 2728 15484
rect 3100 16904 3176 16914
rect 3100 16848 3110 16904
rect 3166 16848 3176 16904
rect 3100 16780 3176 16848
rect 3100 16724 3110 16780
rect 3166 16724 3176 16780
rect 3100 16656 3176 16724
rect 3100 16600 3110 16656
rect 3166 16600 3176 16656
rect 3100 16532 3176 16600
rect 3100 16476 3110 16532
rect 3166 16476 3176 16532
rect 3100 16408 3176 16476
rect 3100 16352 3110 16408
rect 3166 16352 3176 16408
rect 3100 16284 3176 16352
rect 3100 16228 3110 16284
rect 3166 16228 3176 16284
rect 3100 16160 3176 16228
rect 3100 16104 3110 16160
rect 3166 16104 3176 16160
rect 3100 16036 3176 16104
rect 3100 15980 3110 16036
rect 3166 15980 3176 16036
rect 3100 15912 3176 15980
rect 3100 15856 3110 15912
rect 3166 15856 3176 15912
rect 3100 15788 3176 15856
rect 3100 15732 3110 15788
rect 3166 15732 3176 15788
rect 3100 15664 3176 15732
rect 3100 15608 3110 15664
rect 3166 15608 3176 15664
rect 3100 15540 3176 15608
rect 3100 15484 3110 15540
rect 3166 15484 3176 15540
rect 3100 15474 3176 15484
rect 3772 16904 3848 16914
rect 3772 16848 3782 16904
rect 3838 16848 3848 16904
rect 3772 16780 3848 16848
rect 3772 16724 3782 16780
rect 3838 16724 3848 16780
rect 3772 16656 3848 16724
rect 3772 16600 3782 16656
rect 3838 16600 3848 16656
rect 3772 16532 3848 16600
rect 3772 16476 3782 16532
rect 3838 16476 3848 16532
rect 3772 16408 3848 16476
rect 3772 16352 3782 16408
rect 3838 16352 3848 16408
rect 3772 16284 3848 16352
rect 3772 16228 3782 16284
rect 3838 16228 3848 16284
rect 3772 16160 3848 16228
rect 3772 16104 3782 16160
rect 3838 16104 3848 16160
rect 3772 16036 3848 16104
rect 3772 15980 3782 16036
rect 3838 15980 3848 16036
rect 3772 15912 3848 15980
rect 3772 15856 3782 15912
rect 3838 15856 3848 15912
rect 3772 15788 3848 15856
rect 3772 15732 3782 15788
rect 3838 15732 3848 15788
rect 3772 15664 3848 15732
rect 3772 15608 3782 15664
rect 3838 15608 3848 15664
rect 3772 15540 3848 15608
rect 3772 15484 3782 15540
rect 3838 15484 3848 15540
rect 3772 15474 3848 15484
rect 4220 16904 4296 16914
rect 4220 16848 4230 16904
rect 4286 16848 4296 16904
rect 4220 16780 4296 16848
rect 4220 16724 4230 16780
rect 4286 16724 4296 16780
rect 4220 16656 4296 16724
rect 4220 16600 4230 16656
rect 4286 16600 4296 16656
rect 4220 16532 4296 16600
rect 4220 16476 4230 16532
rect 4286 16476 4296 16532
rect 4220 16408 4296 16476
rect 4220 16352 4230 16408
rect 4286 16352 4296 16408
rect 4220 16284 4296 16352
rect 4220 16228 4230 16284
rect 4286 16228 4296 16284
rect 4220 16160 4296 16228
rect 4220 16104 4230 16160
rect 4286 16104 4296 16160
rect 4220 16036 4296 16104
rect 4220 15980 4230 16036
rect 4286 15980 4296 16036
rect 4220 15912 4296 15980
rect 4220 15856 4230 15912
rect 4286 15856 4296 15912
rect 4220 15788 4296 15856
rect 4220 15732 4230 15788
rect 4286 15732 4296 15788
rect 4220 15664 4296 15732
rect 4220 15608 4230 15664
rect 4286 15608 4296 15664
rect 4220 15540 4296 15608
rect 4220 15484 4230 15540
rect 4286 15484 4296 15540
rect 4220 15474 4296 15484
rect 4892 16904 4968 16914
rect 4892 16848 4902 16904
rect 4958 16848 4968 16904
rect 4892 16780 4968 16848
rect 4892 16724 4902 16780
rect 4958 16724 4968 16780
rect 4892 16656 4968 16724
rect 4892 16600 4902 16656
rect 4958 16600 4968 16656
rect 4892 16532 4968 16600
rect 4892 16476 4902 16532
rect 4958 16476 4968 16532
rect 4892 16408 4968 16476
rect 4892 16352 4902 16408
rect 4958 16352 4968 16408
rect 4892 16284 4968 16352
rect 4892 16228 4902 16284
rect 4958 16228 4968 16284
rect 4892 16160 4968 16228
rect 4892 16104 4902 16160
rect 4958 16104 4968 16160
rect 4892 16036 4968 16104
rect 4892 15980 4902 16036
rect 4958 15980 4968 16036
rect 4892 15912 4968 15980
rect 4892 15856 4902 15912
rect 4958 15856 4968 15912
rect 4892 15788 4968 15856
rect 4892 15732 4902 15788
rect 4958 15732 4968 15788
rect 4892 15664 4968 15732
rect 4892 15608 4902 15664
rect 4958 15608 4968 15664
rect 4892 15540 4968 15608
rect 4892 15484 4902 15540
rect 4958 15484 4968 15540
rect 4892 15474 4968 15484
rect 5340 16904 5416 16914
rect 5340 16848 5350 16904
rect 5406 16848 5416 16904
rect 5340 16780 5416 16848
rect 5340 16724 5350 16780
rect 5406 16724 5416 16780
rect 5340 16656 5416 16724
rect 5340 16600 5350 16656
rect 5406 16600 5416 16656
rect 5340 16532 5416 16600
rect 5340 16476 5350 16532
rect 5406 16476 5416 16532
rect 5340 16408 5416 16476
rect 5340 16352 5350 16408
rect 5406 16352 5416 16408
rect 5340 16284 5416 16352
rect 5340 16228 5350 16284
rect 5406 16228 5416 16284
rect 5340 16160 5416 16228
rect 5340 16104 5350 16160
rect 5406 16104 5416 16160
rect 5340 16036 5416 16104
rect 5340 15980 5350 16036
rect 5406 15980 5416 16036
rect 5340 15912 5416 15980
rect 5340 15856 5350 15912
rect 5406 15856 5416 15912
rect 5340 15788 5416 15856
rect 5340 15732 5350 15788
rect 5406 15732 5416 15788
rect 5340 15664 5416 15732
rect 5340 15608 5350 15664
rect 5406 15608 5416 15664
rect 5340 15540 5416 15608
rect 5340 15484 5350 15540
rect 5406 15484 5416 15540
rect 5340 15474 5416 15484
rect 6012 16904 6088 16914
rect 6012 16848 6022 16904
rect 6078 16848 6088 16904
rect 6012 16780 6088 16848
rect 6012 16724 6022 16780
rect 6078 16724 6088 16780
rect 6012 16656 6088 16724
rect 6012 16600 6022 16656
rect 6078 16600 6088 16656
rect 6012 16532 6088 16600
rect 6012 16476 6022 16532
rect 6078 16476 6088 16532
rect 6012 16408 6088 16476
rect 6012 16352 6022 16408
rect 6078 16352 6088 16408
rect 6012 16284 6088 16352
rect 6012 16228 6022 16284
rect 6078 16228 6088 16284
rect 6012 16160 6088 16228
rect 6012 16104 6022 16160
rect 6078 16104 6088 16160
rect 6012 16036 6088 16104
rect 6012 15980 6022 16036
rect 6078 15980 6088 16036
rect 6012 15912 6088 15980
rect 6012 15856 6022 15912
rect 6078 15856 6088 15912
rect 6012 15788 6088 15856
rect 6012 15732 6022 15788
rect 6078 15732 6088 15788
rect 6012 15664 6088 15732
rect 6012 15608 6022 15664
rect 6078 15608 6088 15664
rect 6012 15540 6088 15608
rect 6012 15484 6022 15540
rect 6078 15484 6088 15540
rect 6012 15474 6088 15484
rect 6460 16904 6536 16914
rect 6460 16848 6470 16904
rect 6526 16848 6536 16904
rect 6460 16780 6536 16848
rect 6460 16724 6470 16780
rect 6526 16724 6536 16780
rect 6460 16656 6536 16724
rect 6460 16600 6470 16656
rect 6526 16600 6536 16656
rect 6460 16532 6536 16600
rect 6460 16476 6470 16532
rect 6526 16476 6536 16532
rect 6460 16408 6536 16476
rect 6460 16352 6470 16408
rect 6526 16352 6536 16408
rect 6460 16284 6536 16352
rect 6460 16228 6470 16284
rect 6526 16228 6536 16284
rect 6460 16160 6536 16228
rect 6460 16104 6470 16160
rect 6526 16104 6536 16160
rect 6460 16036 6536 16104
rect 6460 15980 6470 16036
rect 6526 15980 6536 16036
rect 6460 15912 6536 15980
rect 6460 15856 6470 15912
rect 6526 15856 6536 15912
rect 6460 15788 6536 15856
rect 6460 15732 6470 15788
rect 6526 15732 6536 15788
rect 6460 15664 6536 15732
rect 6460 15608 6470 15664
rect 6526 15608 6536 15664
rect 6460 15540 6536 15608
rect 6460 15484 6470 15540
rect 6526 15484 6536 15540
rect 6460 15474 6536 15484
rect 7132 16904 7208 16914
rect 7132 16848 7142 16904
rect 7198 16848 7208 16904
rect 7132 16780 7208 16848
rect 7132 16724 7142 16780
rect 7198 16724 7208 16780
rect 7132 16656 7208 16724
rect 7132 16600 7142 16656
rect 7198 16600 7208 16656
rect 7132 16532 7208 16600
rect 7132 16476 7142 16532
rect 7198 16476 7208 16532
rect 7132 16408 7208 16476
rect 7132 16352 7142 16408
rect 7198 16352 7208 16408
rect 7132 16284 7208 16352
rect 7132 16228 7142 16284
rect 7198 16228 7208 16284
rect 7132 16160 7208 16228
rect 7132 16104 7142 16160
rect 7198 16104 7208 16160
rect 7132 16036 7208 16104
rect 7132 15980 7142 16036
rect 7198 15980 7208 16036
rect 7132 15912 7208 15980
rect 7132 15856 7142 15912
rect 7198 15856 7208 15912
rect 7132 15788 7208 15856
rect 7132 15732 7142 15788
rect 7198 15732 7208 15788
rect 7132 15664 7208 15732
rect 7132 15608 7142 15664
rect 7198 15608 7208 15664
rect 7132 15540 7208 15608
rect 7132 15484 7142 15540
rect 7198 15484 7208 15540
rect 7132 15474 7208 15484
rect 7580 16904 7656 16914
rect 7580 16848 7590 16904
rect 7646 16848 7656 16904
rect 7580 16780 7656 16848
rect 7580 16724 7590 16780
rect 7646 16724 7656 16780
rect 7580 16656 7656 16724
rect 7580 16600 7590 16656
rect 7646 16600 7656 16656
rect 7580 16532 7656 16600
rect 7580 16476 7590 16532
rect 7646 16476 7656 16532
rect 7580 16408 7656 16476
rect 7580 16352 7590 16408
rect 7646 16352 7656 16408
rect 7580 16284 7656 16352
rect 7580 16228 7590 16284
rect 7646 16228 7656 16284
rect 7580 16160 7656 16228
rect 7580 16104 7590 16160
rect 7646 16104 7656 16160
rect 7580 16036 7656 16104
rect 7580 15980 7590 16036
rect 7646 15980 7656 16036
rect 7580 15912 7656 15980
rect 7580 15856 7590 15912
rect 7646 15856 7656 15912
rect 7580 15788 7656 15856
rect 7580 15732 7590 15788
rect 7646 15732 7656 15788
rect 7580 15664 7656 15732
rect 7580 15608 7590 15664
rect 7646 15608 7656 15664
rect 7580 15540 7656 15608
rect 7580 15484 7590 15540
rect 7646 15484 7656 15540
rect 7580 15474 7656 15484
rect 8252 16904 8328 16914
rect 8252 16848 8262 16904
rect 8318 16848 8328 16904
rect 8252 16780 8328 16848
rect 8252 16724 8262 16780
rect 8318 16724 8328 16780
rect 8252 16656 8328 16724
rect 8252 16600 8262 16656
rect 8318 16600 8328 16656
rect 8252 16532 8328 16600
rect 8252 16476 8262 16532
rect 8318 16476 8328 16532
rect 8252 16408 8328 16476
rect 8252 16352 8262 16408
rect 8318 16352 8328 16408
rect 8252 16284 8328 16352
rect 8252 16228 8262 16284
rect 8318 16228 8328 16284
rect 8252 16160 8328 16228
rect 8252 16104 8262 16160
rect 8318 16104 8328 16160
rect 8252 16036 8328 16104
rect 8252 15980 8262 16036
rect 8318 15980 8328 16036
rect 8252 15912 8328 15980
rect 8252 15856 8262 15912
rect 8318 15856 8328 15912
rect 8252 15788 8328 15856
rect 8252 15732 8262 15788
rect 8318 15732 8328 15788
rect 8252 15664 8328 15732
rect 8252 15608 8262 15664
rect 8318 15608 8328 15664
rect 8252 15540 8328 15608
rect 8252 15484 8262 15540
rect 8318 15484 8328 15540
rect 8252 15474 8328 15484
rect 8700 16904 8776 16914
rect 8700 16848 8710 16904
rect 8766 16848 8776 16904
rect 8700 16780 8776 16848
rect 8700 16724 8710 16780
rect 8766 16724 8776 16780
rect 8700 16656 8776 16724
rect 8700 16600 8710 16656
rect 8766 16600 8776 16656
rect 8700 16532 8776 16600
rect 8700 16476 8710 16532
rect 8766 16476 8776 16532
rect 8700 16408 8776 16476
rect 8700 16352 8710 16408
rect 8766 16352 8776 16408
rect 8700 16284 8776 16352
rect 8700 16228 8710 16284
rect 8766 16228 8776 16284
rect 8700 16160 8776 16228
rect 8700 16104 8710 16160
rect 8766 16104 8776 16160
rect 8700 16036 8776 16104
rect 8700 15980 8710 16036
rect 8766 15980 8776 16036
rect 8700 15912 8776 15980
rect 8700 15856 8710 15912
rect 8766 15856 8776 15912
rect 8700 15788 8776 15856
rect 8700 15732 8710 15788
rect 8766 15732 8776 15788
rect 8700 15664 8776 15732
rect 8700 15608 8710 15664
rect 8766 15608 8776 15664
rect 8700 15540 8776 15608
rect 8700 15484 8710 15540
rect 8766 15484 8776 15540
rect 8700 15474 8776 15484
rect 9372 16904 9448 16914
rect 9372 16848 9382 16904
rect 9438 16848 9448 16904
rect 9372 16780 9448 16848
rect 9372 16724 9382 16780
rect 9438 16724 9448 16780
rect 9372 16656 9448 16724
rect 9372 16600 9382 16656
rect 9438 16600 9448 16656
rect 9372 16532 9448 16600
rect 9372 16476 9382 16532
rect 9438 16476 9448 16532
rect 9372 16408 9448 16476
rect 9372 16352 9382 16408
rect 9438 16352 9448 16408
rect 9372 16284 9448 16352
rect 9372 16228 9382 16284
rect 9438 16228 9448 16284
rect 9372 16160 9448 16228
rect 9372 16104 9382 16160
rect 9438 16104 9448 16160
rect 9372 16036 9448 16104
rect 9372 15980 9382 16036
rect 9438 15980 9448 16036
rect 9372 15912 9448 15980
rect 9372 15856 9382 15912
rect 9438 15856 9448 15912
rect 9372 15788 9448 15856
rect 9372 15732 9382 15788
rect 9438 15732 9448 15788
rect 9372 15664 9448 15732
rect 9372 15608 9382 15664
rect 9438 15608 9448 15664
rect 9372 15540 9448 15608
rect 9372 15484 9382 15540
rect 9438 15484 9448 15540
rect 9372 15474 9448 15484
rect 9820 16904 9896 16914
rect 9820 16848 9830 16904
rect 9886 16848 9896 16904
rect 9820 16780 9896 16848
rect 9820 16724 9830 16780
rect 9886 16724 9896 16780
rect 9820 16656 9896 16724
rect 9820 16600 9830 16656
rect 9886 16600 9896 16656
rect 9820 16532 9896 16600
rect 9820 16476 9830 16532
rect 9886 16476 9896 16532
rect 9820 16408 9896 16476
rect 9820 16352 9830 16408
rect 9886 16352 9896 16408
rect 9820 16284 9896 16352
rect 9820 16228 9830 16284
rect 9886 16228 9896 16284
rect 9820 16160 9896 16228
rect 9820 16104 9830 16160
rect 9886 16104 9896 16160
rect 9820 16036 9896 16104
rect 9820 15980 9830 16036
rect 9886 15980 9896 16036
rect 9820 15912 9896 15980
rect 9820 15856 9830 15912
rect 9886 15856 9896 15912
rect 9820 15788 9896 15856
rect 9820 15732 9830 15788
rect 9886 15732 9896 15788
rect 9820 15664 9896 15732
rect 9820 15608 9830 15664
rect 9886 15608 9896 15664
rect 9820 15540 9896 15608
rect 9820 15484 9830 15540
rect 9886 15484 9896 15540
rect 9820 15474 9896 15484
rect 10492 16904 10568 16914
rect 10492 16848 10502 16904
rect 10558 16848 10568 16904
rect 10492 16780 10568 16848
rect 10492 16724 10502 16780
rect 10558 16724 10568 16780
rect 10492 16656 10568 16724
rect 10492 16600 10502 16656
rect 10558 16600 10568 16656
rect 10492 16532 10568 16600
rect 10492 16476 10502 16532
rect 10558 16476 10568 16532
rect 10492 16408 10568 16476
rect 10492 16352 10502 16408
rect 10558 16352 10568 16408
rect 10492 16284 10568 16352
rect 10492 16228 10502 16284
rect 10558 16228 10568 16284
rect 10492 16160 10568 16228
rect 10492 16104 10502 16160
rect 10558 16104 10568 16160
rect 10492 16036 10568 16104
rect 10492 15980 10502 16036
rect 10558 15980 10568 16036
rect 10492 15912 10568 15980
rect 10492 15856 10502 15912
rect 10558 15856 10568 15912
rect 10492 15788 10568 15856
rect 10492 15732 10502 15788
rect 10558 15732 10568 15788
rect 10492 15664 10568 15732
rect 10492 15608 10502 15664
rect 10558 15608 10568 15664
rect 10492 15540 10568 15608
rect 10492 15484 10502 15540
rect 10558 15484 10568 15540
rect 10492 15474 10568 15484
rect 10940 16904 11016 16914
rect 10940 16848 10950 16904
rect 11006 16848 11016 16904
rect 10940 16780 11016 16848
rect 10940 16724 10950 16780
rect 11006 16724 11016 16780
rect 10940 16656 11016 16724
rect 10940 16600 10950 16656
rect 11006 16600 11016 16656
rect 10940 16532 11016 16600
rect 10940 16476 10950 16532
rect 11006 16476 11016 16532
rect 10940 16408 11016 16476
rect 10940 16352 10950 16408
rect 11006 16352 11016 16408
rect 10940 16284 11016 16352
rect 10940 16228 10950 16284
rect 11006 16228 11016 16284
rect 10940 16160 11016 16228
rect 10940 16104 10950 16160
rect 11006 16104 11016 16160
rect 10940 16036 11016 16104
rect 10940 15980 10950 16036
rect 11006 15980 11016 16036
rect 10940 15912 11016 15980
rect 10940 15856 10950 15912
rect 11006 15856 11016 15912
rect 10940 15788 11016 15856
rect 10940 15732 10950 15788
rect 11006 15732 11016 15788
rect 10940 15664 11016 15732
rect 10940 15608 10950 15664
rect 11006 15608 11016 15664
rect 10940 15540 11016 15608
rect 10940 15484 10950 15540
rect 11006 15484 11016 15540
rect 10940 15474 11016 15484
rect 11612 16904 11688 16914
rect 11612 16848 11622 16904
rect 11678 16848 11688 16904
rect 11612 16780 11688 16848
rect 11612 16724 11622 16780
rect 11678 16724 11688 16780
rect 11612 16656 11688 16724
rect 11612 16600 11622 16656
rect 11678 16600 11688 16656
rect 11612 16532 11688 16600
rect 11612 16476 11622 16532
rect 11678 16476 11688 16532
rect 11612 16408 11688 16476
rect 11612 16352 11622 16408
rect 11678 16352 11688 16408
rect 11612 16284 11688 16352
rect 11612 16228 11622 16284
rect 11678 16228 11688 16284
rect 11612 16160 11688 16228
rect 11612 16104 11622 16160
rect 11678 16104 11688 16160
rect 11612 16036 11688 16104
rect 11612 15980 11622 16036
rect 11678 15980 11688 16036
rect 11612 15912 11688 15980
rect 11612 15856 11622 15912
rect 11678 15856 11688 15912
rect 11612 15788 11688 15856
rect 11612 15732 11622 15788
rect 11678 15732 11688 15788
rect 11612 15664 11688 15732
rect 11612 15608 11622 15664
rect 11678 15608 11688 15664
rect 11612 15540 11688 15608
rect 11612 15484 11622 15540
rect 11678 15484 11688 15540
rect 11612 15474 11688 15484
rect 12060 16904 12136 16914
rect 12060 16848 12070 16904
rect 12126 16848 12136 16904
rect 12060 16780 12136 16848
rect 12060 16724 12070 16780
rect 12126 16724 12136 16780
rect 12060 16656 12136 16724
rect 12060 16600 12070 16656
rect 12126 16600 12136 16656
rect 12060 16532 12136 16600
rect 12060 16476 12070 16532
rect 12126 16476 12136 16532
rect 12060 16408 12136 16476
rect 12060 16352 12070 16408
rect 12126 16352 12136 16408
rect 12060 16284 12136 16352
rect 12060 16228 12070 16284
rect 12126 16228 12136 16284
rect 12060 16160 12136 16228
rect 12060 16104 12070 16160
rect 12126 16104 12136 16160
rect 12060 16036 12136 16104
rect 12060 15980 12070 16036
rect 12126 15980 12136 16036
rect 12060 15912 12136 15980
rect 12060 15856 12070 15912
rect 12126 15856 12136 15912
rect 12060 15788 12136 15856
rect 12060 15732 12070 15788
rect 12126 15732 12136 15788
rect 12060 15664 12136 15732
rect 12060 15608 12070 15664
rect 12126 15608 12136 15664
rect 12060 15540 12136 15608
rect 12060 15484 12070 15540
rect 12126 15484 12136 15540
rect 12060 15474 12136 15484
rect 12732 16904 12808 16914
rect 12732 16848 12742 16904
rect 12798 16848 12808 16904
rect 12732 16780 12808 16848
rect 12732 16724 12742 16780
rect 12798 16724 12808 16780
rect 12732 16656 12808 16724
rect 12732 16600 12742 16656
rect 12798 16600 12808 16656
rect 12732 16532 12808 16600
rect 12732 16476 12742 16532
rect 12798 16476 12808 16532
rect 12732 16408 12808 16476
rect 12732 16352 12742 16408
rect 12798 16352 12808 16408
rect 12732 16284 12808 16352
rect 12732 16228 12742 16284
rect 12798 16228 12808 16284
rect 12732 16160 12808 16228
rect 12732 16104 12742 16160
rect 12798 16104 12808 16160
rect 12732 16036 12808 16104
rect 12732 15980 12742 16036
rect 12798 15980 12808 16036
rect 12732 15912 12808 15980
rect 12732 15856 12742 15912
rect 12798 15856 12808 15912
rect 12732 15788 12808 15856
rect 12732 15732 12742 15788
rect 12798 15732 12808 15788
rect 12732 15664 12808 15732
rect 12732 15608 12742 15664
rect 12798 15608 12808 15664
rect 12732 15540 12808 15608
rect 12732 15484 12742 15540
rect 12798 15484 12808 15540
rect 12732 15474 12808 15484
rect 13180 16904 13256 16914
rect 13180 16848 13190 16904
rect 13246 16848 13256 16904
rect 13180 16780 13256 16848
rect 13180 16724 13190 16780
rect 13246 16724 13256 16780
rect 13180 16656 13256 16724
rect 13180 16600 13190 16656
rect 13246 16600 13256 16656
rect 13180 16532 13256 16600
rect 13180 16476 13190 16532
rect 13246 16476 13256 16532
rect 13180 16408 13256 16476
rect 13180 16352 13190 16408
rect 13246 16352 13256 16408
rect 13180 16284 13256 16352
rect 13180 16228 13190 16284
rect 13246 16228 13256 16284
rect 13180 16160 13256 16228
rect 13180 16104 13190 16160
rect 13246 16104 13256 16160
rect 13180 16036 13256 16104
rect 13180 15980 13190 16036
rect 13246 15980 13256 16036
rect 13180 15912 13256 15980
rect 13180 15856 13190 15912
rect 13246 15856 13256 15912
rect 13180 15788 13256 15856
rect 13180 15732 13190 15788
rect 13246 15732 13256 15788
rect 13180 15664 13256 15732
rect 13180 15608 13190 15664
rect 13246 15608 13256 15664
rect 13180 15540 13256 15608
rect 13180 15484 13190 15540
rect 13246 15484 13256 15540
rect 13180 15474 13256 15484
rect 13852 16904 13928 16914
rect 13852 16848 13862 16904
rect 13918 16848 13928 16904
rect 13852 16780 13928 16848
rect 13852 16724 13862 16780
rect 13918 16724 13928 16780
rect 13852 16656 13928 16724
rect 13852 16600 13862 16656
rect 13918 16600 13928 16656
rect 13852 16532 13928 16600
rect 13852 16476 13862 16532
rect 13918 16476 13928 16532
rect 13852 16408 13928 16476
rect 13852 16352 13862 16408
rect 13918 16352 13928 16408
rect 13852 16284 13928 16352
rect 13852 16228 13862 16284
rect 13918 16228 13928 16284
rect 13852 16160 13928 16228
rect 13852 16104 13862 16160
rect 13918 16104 13928 16160
rect 13852 16036 13928 16104
rect 13852 15980 13862 16036
rect 13918 15980 13928 16036
rect 13852 15912 13928 15980
rect 13852 15856 13862 15912
rect 13918 15856 13928 15912
rect 13852 15788 13928 15856
rect 13852 15732 13862 15788
rect 13918 15732 13928 15788
rect 13852 15664 13928 15732
rect 13852 15608 13862 15664
rect 13918 15608 13928 15664
rect 13852 15540 13928 15608
rect 13852 15484 13862 15540
rect 13918 15484 13928 15540
rect 13852 15474 13928 15484
rect 14300 16904 14376 16914
rect 14300 16848 14310 16904
rect 14366 16848 14376 16904
rect 14300 16780 14376 16848
rect 14300 16724 14310 16780
rect 14366 16724 14376 16780
rect 14300 16656 14376 16724
rect 14300 16600 14310 16656
rect 14366 16600 14376 16656
rect 14300 16532 14376 16600
rect 14300 16476 14310 16532
rect 14366 16476 14376 16532
rect 14300 16408 14376 16476
rect 14300 16352 14310 16408
rect 14366 16352 14376 16408
rect 14300 16284 14376 16352
rect 14300 16228 14310 16284
rect 14366 16228 14376 16284
rect 14300 16160 14376 16228
rect 14300 16104 14310 16160
rect 14366 16104 14376 16160
rect 14300 16036 14376 16104
rect 14300 15980 14310 16036
rect 14366 15980 14376 16036
rect 14300 15912 14376 15980
rect 14300 15856 14310 15912
rect 14366 15856 14376 15912
rect 14300 15788 14376 15856
rect 14300 15732 14310 15788
rect 14366 15732 14376 15788
rect 14300 15664 14376 15732
rect 14300 15608 14310 15664
rect 14366 15608 14376 15664
rect 14300 15540 14376 15608
rect 14300 15484 14310 15540
rect 14366 15484 14376 15540
rect 14300 15474 14376 15484
rect 14972 16904 15048 16914
rect 14972 16848 14982 16904
rect 15038 16848 15048 16904
rect 14972 16780 15048 16848
rect 14972 16724 14982 16780
rect 15038 16724 15048 16780
rect 14972 16656 15048 16724
rect 14972 16600 14982 16656
rect 15038 16600 15048 16656
rect 14972 16532 15048 16600
rect 14972 16476 14982 16532
rect 15038 16476 15048 16532
rect 14972 16408 15048 16476
rect 14972 16352 14982 16408
rect 15038 16352 15048 16408
rect 14972 16284 15048 16352
rect 14972 16228 14982 16284
rect 15038 16228 15048 16284
rect 14972 16160 15048 16228
rect 14972 16104 14982 16160
rect 15038 16104 15048 16160
rect 14972 16036 15048 16104
rect 14972 15980 14982 16036
rect 15038 15980 15048 16036
rect 14972 15912 15048 15980
rect 14972 15856 14982 15912
rect 15038 15856 15048 15912
rect 14972 15788 15048 15856
rect 14972 15732 14982 15788
rect 15038 15732 15048 15788
rect 14972 15664 15048 15732
rect 14972 15608 14982 15664
rect 15038 15608 15048 15664
rect 14972 15540 15048 15608
rect 14972 15484 14982 15540
rect 15038 15484 15048 15540
rect 14972 15474 15048 15484
rect 15420 16904 15496 16914
rect 15420 16848 15430 16904
rect 15486 16848 15496 16904
rect 15420 16780 15496 16848
rect 15420 16724 15430 16780
rect 15486 16724 15496 16780
rect 15420 16656 15496 16724
rect 15420 16600 15430 16656
rect 15486 16600 15496 16656
rect 15420 16532 15496 16600
rect 15420 16476 15430 16532
rect 15486 16476 15496 16532
rect 15420 16408 15496 16476
rect 15420 16352 15430 16408
rect 15486 16352 15496 16408
rect 15420 16284 15496 16352
rect 15420 16228 15430 16284
rect 15486 16228 15496 16284
rect 15420 16160 15496 16228
rect 15420 16104 15430 16160
rect 15486 16104 15496 16160
rect 15420 16036 15496 16104
rect 15420 15980 15430 16036
rect 15486 15980 15496 16036
rect 15420 15912 15496 15980
rect 15420 15856 15430 15912
rect 15486 15856 15496 15912
rect 15420 15788 15496 15856
rect 15420 15732 15430 15788
rect 15486 15732 15496 15788
rect 15420 15664 15496 15732
rect 15420 15608 15430 15664
rect 15486 15608 15496 15664
rect 15420 15540 15496 15608
rect 15420 15484 15430 15540
rect 15486 15484 15496 15540
rect 15420 15474 15496 15484
rect 16092 16904 16168 16914
rect 16092 16848 16102 16904
rect 16158 16848 16168 16904
rect 16092 16780 16168 16848
rect 16092 16724 16102 16780
rect 16158 16724 16168 16780
rect 16092 16656 16168 16724
rect 16092 16600 16102 16656
rect 16158 16600 16168 16656
rect 16092 16532 16168 16600
rect 16092 16476 16102 16532
rect 16158 16476 16168 16532
rect 16092 16408 16168 16476
rect 16092 16352 16102 16408
rect 16158 16352 16168 16408
rect 16092 16284 16168 16352
rect 16092 16228 16102 16284
rect 16158 16228 16168 16284
rect 16092 16160 16168 16228
rect 16092 16104 16102 16160
rect 16158 16104 16168 16160
rect 16092 16036 16168 16104
rect 16092 15980 16102 16036
rect 16158 15980 16168 16036
rect 16092 15912 16168 15980
rect 16092 15856 16102 15912
rect 16158 15856 16168 15912
rect 16092 15788 16168 15856
rect 16092 15732 16102 15788
rect 16158 15732 16168 15788
rect 16092 15664 16168 15732
rect 16092 15608 16102 15664
rect 16158 15608 16168 15664
rect 16092 15540 16168 15608
rect 16092 15484 16102 15540
rect 16158 15484 16168 15540
rect 16092 15474 16168 15484
rect 16540 16904 16616 16914
rect 16540 16848 16550 16904
rect 16606 16848 16616 16904
rect 16540 16780 16616 16848
rect 16540 16724 16550 16780
rect 16606 16724 16616 16780
rect 16540 16656 16616 16724
rect 16540 16600 16550 16656
rect 16606 16600 16616 16656
rect 16540 16532 16616 16600
rect 16540 16476 16550 16532
rect 16606 16476 16616 16532
rect 16540 16408 16616 16476
rect 16540 16352 16550 16408
rect 16606 16352 16616 16408
rect 16540 16284 16616 16352
rect 16540 16228 16550 16284
rect 16606 16228 16616 16284
rect 16540 16160 16616 16228
rect 16540 16104 16550 16160
rect 16606 16104 16616 16160
rect 16540 16036 16616 16104
rect 16540 15980 16550 16036
rect 16606 15980 16616 16036
rect 16540 15912 16616 15980
rect 16540 15856 16550 15912
rect 16606 15856 16616 15912
rect 16540 15788 16616 15856
rect 16540 15732 16550 15788
rect 16606 15732 16616 15788
rect 16540 15664 16616 15732
rect 16540 15608 16550 15664
rect 16606 15608 16616 15664
rect 16540 15540 16616 15608
rect 16540 15484 16550 15540
rect 16606 15484 16616 15540
rect 16540 15474 16616 15484
rect 17212 16904 17288 16914
rect 17212 16848 17222 16904
rect 17278 16848 17288 16904
rect 17212 16780 17288 16848
rect 17212 16724 17222 16780
rect 17278 16724 17288 16780
rect 17212 16656 17288 16724
rect 17212 16600 17222 16656
rect 17278 16600 17288 16656
rect 17212 16532 17288 16600
rect 17212 16476 17222 16532
rect 17278 16476 17288 16532
rect 17212 16408 17288 16476
rect 17212 16352 17222 16408
rect 17278 16352 17288 16408
rect 17212 16284 17288 16352
rect 17212 16228 17222 16284
rect 17278 16228 17288 16284
rect 17212 16160 17288 16228
rect 17212 16104 17222 16160
rect 17278 16104 17288 16160
rect 17212 16036 17288 16104
rect 17212 15980 17222 16036
rect 17278 15980 17288 16036
rect 17212 15912 17288 15980
rect 17212 15856 17222 15912
rect 17278 15856 17288 15912
rect 17212 15788 17288 15856
rect 17212 15732 17222 15788
rect 17278 15732 17288 15788
rect 17212 15664 17288 15732
rect 17212 15608 17222 15664
rect 17278 15608 17288 15664
rect 17212 15540 17288 15608
rect 17212 15484 17222 15540
rect 17278 15484 17288 15540
rect 17212 15474 17288 15484
rect 17660 16904 17736 16914
rect 17660 16848 17670 16904
rect 17726 16848 17736 16904
rect 17660 16780 17736 16848
rect 17660 16724 17670 16780
rect 17726 16724 17736 16780
rect 17660 16656 17736 16724
rect 17660 16600 17670 16656
rect 17726 16600 17736 16656
rect 17660 16532 17736 16600
rect 17660 16476 17670 16532
rect 17726 16476 17736 16532
rect 17660 16408 17736 16476
rect 17660 16352 17670 16408
rect 17726 16352 17736 16408
rect 17660 16284 17736 16352
rect 17660 16228 17670 16284
rect 17726 16228 17736 16284
rect 17660 16160 17736 16228
rect 17660 16104 17670 16160
rect 17726 16104 17736 16160
rect 17660 16036 17736 16104
rect 17660 15980 17670 16036
rect 17726 15980 17736 16036
rect 17660 15912 17736 15980
rect 17660 15856 17670 15912
rect 17726 15856 17736 15912
rect 17660 15788 17736 15856
rect 17660 15732 17670 15788
rect 17726 15732 17736 15788
rect 17660 15664 17736 15732
rect 17660 15608 17670 15664
rect 17726 15608 17736 15664
rect 17660 15540 17736 15608
rect 17660 15484 17670 15540
rect 17726 15484 17736 15540
rect 17660 15474 17736 15484
rect 18332 16904 18408 16914
rect 18332 16848 18342 16904
rect 18398 16848 18408 16904
rect 18332 16780 18408 16848
rect 18332 16724 18342 16780
rect 18398 16724 18408 16780
rect 18332 16656 18408 16724
rect 18332 16600 18342 16656
rect 18398 16600 18408 16656
rect 18332 16532 18408 16600
rect 18332 16476 18342 16532
rect 18398 16476 18408 16532
rect 18332 16408 18408 16476
rect 18332 16352 18342 16408
rect 18398 16352 18408 16408
rect 18332 16284 18408 16352
rect 18332 16228 18342 16284
rect 18398 16228 18408 16284
rect 18332 16160 18408 16228
rect 18332 16104 18342 16160
rect 18398 16104 18408 16160
rect 18332 16036 18408 16104
rect 18332 15980 18342 16036
rect 18398 15980 18408 16036
rect 18332 15912 18408 15980
rect 18332 15856 18342 15912
rect 18398 15856 18408 15912
rect 18332 15788 18408 15856
rect 18332 15732 18342 15788
rect 18398 15732 18408 15788
rect 18332 15664 18408 15732
rect 18332 15608 18342 15664
rect 18398 15608 18408 15664
rect 18332 15540 18408 15608
rect 18332 15484 18342 15540
rect 18398 15484 18408 15540
rect 18332 15474 18408 15484
rect 18780 16904 18856 16914
rect 18780 16848 18790 16904
rect 18846 16848 18856 16904
rect 18780 16780 18856 16848
rect 18780 16724 18790 16780
rect 18846 16724 18856 16780
rect 18780 16656 18856 16724
rect 18780 16600 18790 16656
rect 18846 16600 18856 16656
rect 18780 16532 18856 16600
rect 18780 16476 18790 16532
rect 18846 16476 18856 16532
rect 18780 16408 18856 16476
rect 18780 16352 18790 16408
rect 18846 16352 18856 16408
rect 18780 16284 18856 16352
rect 18780 16228 18790 16284
rect 18846 16228 18856 16284
rect 18780 16160 18856 16228
rect 18780 16104 18790 16160
rect 18846 16104 18856 16160
rect 18780 16036 18856 16104
rect 18780 15980 18790 16036
rect 18846 15980 18856 16036
rect 18780 15912 18856 15980
rect 18780 15856 18790 15912
rect 18846 15856 18856 15912
rect 18780 15788 18856 15856
rect 18780 15732 18790 15788
rect 18846 15732 18856 15788
rect 18780 15664 18856 15732
rect 18780 15608 18790 15664
rect 18846 15608 18856 15664
rect 18780 15540 18856 15608
rect 18780 15484 18790 15540
rect 18846 15484 18856 15540
rect 18780 15474 18856 15484
rect 19452 16904 19528 16914
rect 19452 16848 19462 16904
rect 19518 16848 19528 16904
rect 19452 16780 19528 16848
rect 19452 16724 19462 16780
rect 19518 16724 19528 16780
rect 19452 16656 19528 16724
rect 19452 16600 19462 16656
rect 19518 16600 19528 16656
rect 19452 16532 19528 16600
rect 19452 16476 19462 16532
rect 19518 16476 19528 16532
rect 19452 16408 19528 16476
rect 19452 16352 19462 16408
rect 19518 16352 19528 16408
rect 19452 16284 19528 16352
rect 19452 16228 19462 16284
rect 19518 16228 19528 16284
rect 19452 16160 19528 16228
rect 19452 16104 19462 16160
rect 19518 16104 19528 16160
rect 19452 16036 19528 16104
rect 19452 15980 19462 16036
rect 19518 15980 19528 16036
rect 19452 15912 19528 15980
rect 19452 15856 19462 15912
rect 19518 15856 19528 15912
rect 19452 15788 19528 15856
rect 19452 15732 19462 15788
rect 19518 15732 19528 15788
rect 19452 15664 19528 15732
rect 19452 15608 19462 15664
rect 19518 15608 19528 15664
rect 19452 15540 19528 15608
rect 19452 15484 19462 15540
rect 19518 15484 19528 15540
rect 19452 15474 19528 15484
rect 19900 16904 19976 16914
rect 19900 16848 19910 16904
rect 19966 16848 19976 16904
rect 19900 16780 19976 16848
rect 19900 16724 19910 16780
rect 19966 16724 19976 16780
rect 19900 16656 19976 16724
rect 19900 16600 19910 16656
rect 19966 16600 19976 16656
rect 19900 16532 19976 16600
rect 19900 16476 19910 16532
rect 19966 16476 19976 16532
rect 19900 16408 19976 16476
rect 19900 16352 19910 16408
rect 19966 16352 19976 16408
rect 19900 16284 19976 16352
rect 19900 16228 19910 16284
rect 19966 16228 19976 16284
rect 19900 16160 19976 16228
rect 19900 16104 19910 16160
rect 19966 16104 19976 16160
rect 19900 16036 19976 16104
rect 19900 15980 19910 16036
rect 19966 15980 19976 16036
rect 19900 15912 19976 15980
rect 19900 15856 19910 15912
rect 19966 15856 19976 15912
rect 19900 15788 19976 15856
rect 19900 15732 19910 15788
rect 19966 15732 19976 15788
rect 19900 15664 19976 15732
rect 19900 15608 19910 15664
rect 19966 15608 19976 15664
rect 19900 15540 19976 15608
rect 19900 15484 19910 15540
rect 19966 15484 19976 15540
rect 19900 15474 19976 15484
rect 2428 14996 2504 15008
rect 2428 14944 2440 14996
rect 2492 14944 2504 14996
rect 2428 14872 2504 14944
rect 2428 14820 2440 14872
rect 2492 14820 2504 14872
rect 2428 14748 2504 14820
rect 2428 14696 2440 14748
rect 2492 14696 2504 14748
rect 2428 14624 2504 14696
rect 2428 14572 2440 14624
rect 2492 14572 2504 14624
rect 2428 14500 2504 14572
rect 2428 14448 2440 14500
rect 2492 14448 2504 14500
rect 2428 14376 2504 14448
rect 2428 14324 2440 14376
rect 2492 14324 2504 14376
rect 2428 14252 2504 14324
rect 2428 14200 2440 14252
rect 2492 14200 2504 14252
rect 2428 14128 2504 14200
rect 2428 14076 2440 14128
rect 2492 14076 2504 14128
rect 2428 14004 2504 14076
rect 2428 13952 2440 14004
rect 2492 13952 2504 14004
rect 2428 13880 2504 13952
rect 2428 13828 2440 13880
rect 2492 13828 2504 13880
rect 2428 13756 2504 13828
rect 2428 13704 2440 13756
rect 2492 13704 2504 13756
rect 2428 13632 2504 13704
rect 2428 13580 2440 13632
rect 2492 13580 2504 13632
rect 2428 13508 2504 13580
rect 2428 13456 2440 13508
rect 2492 13456 2504 13508
rect 2428 13384 2504 13456
rect 2428 13332 2440 13384
rect 2492 13332 2504 13384
rect 2428 13260 2504 13332
rect 2428 13208 2440 13260
rect 2492 13208 2504 13260
rect 2428 13136 2504 13208
rect 2428 13084 2440 13136
rect 2492 13084 2504 13136
rect 2428 13012 2504 13084
rect 2428 12960 2440 13012
rect 2492 12960 2504 13012
rect 2428 12888 2504 12960
rect 2428 12836 2440 12888
rect 2492 12836 2504 12888
rect 2428 12592 2504 12836
rect 2876 14996 2952 15008
rect 2876 14944 2888 14996
rect 2940 14944 2952 14996
rect 2876 14872 2952 14944
rect 2876 14820 2888 14872
rect 2940 14820 2952 14872
rect 2876 14748 2952 14820
rect 2876 14696 2888 14748
rect 2940 14696 2952 14748
rect 2876 14624 2952 14696
rect 2876 14572 2888 14624
rect 2940 14572 2952 14624
rect 2876 14500 2952 14572
rect 2876 14448 2888 14500
rect 2940 14448 2952 14500
rect 2876 14376 2952 14448
rect 2876 14324 2888 14376
rect 2940 14324 2952 14376
rect 2876 14252 2952 14324
rect 2876 14200 2888 14252
rect 2940 14200 2952 14252
rect 2876 14128 2952 14200
rect 2876 14076 2888 14128
rect 2940 14076 2952 14128
rect 2876 14004 2952 14076
rect 2876 13952 2888 14004
rect 2940 13952 2952 14004
rect 2876 13880 2952 13952
rect 2876 13828 2888 13880
rect 2940 13828 2952 13880
rect 2876 13756 2952 13828
rect 2876 13704 2888 13756
rect 2940 13704 2952 13756
rect 2876 13632 2952 13704
rect 2876 13580 2888 13632
rect 2940 13580 2952 13632
rect 2876 13508 2952 13580
rect 2876 13456 2888 13508
rect 2940 13456 2952 13508
rect 2876 13384 2952 13456
rect 2876 13332 2888 13384
rect 2940 13332 2952 13384
rect 2876 13260 2952 13332
rect 2876 13208 2888 13260
rect 2940 13208 2952 13260
rect 2876 13136 2952 13208
rect 2876 13084 2888 13136
rect 2940 13084 2952 13136
rect 2876 13012 2952 13084
rect 2876 12960 2888 13012
rect 2940 12960 2952 13012
rect 2876 12888 2952 12960
rect 3548 14996 3624 15008
rect 3548 14944 3560 14996
rect 3612 14944 3624 14996
rect 3548 14872 3624 14944
rect 3548 14820 3560 14872
rect 3612 14820 3624 14872
rect 3548 14748 3624 14820
rect 3548 14696 3560 14748
rect 3612 14696 3624 14748
rect 3548 14624 3624 14696
rect 3548 14572 3560 14624
rect 3612 14572 3624 14624
rect 3548 14500 3624 14572
rect 3548 14448 3560 14500
rect 3612 14448 3624 14500
rect 3548 14376 3624 14448
rect 3548 14324 3560 14376
rect 3612 14324 3624 14376
rect 3548 14252 3624 14324
rect 3548 14200 3560 14252
rect 3612 14200 3624 14252
rect 3548 14128 3624 14200
rect 3548 14076 3560 14128
rect 3612 14076 3624 14128
rect 3548 14004 3624 14076
rect 3548 13952 3560 14004
rect 3612 13952 3624 14004
rect 3548 13880 3624 13952
rect 3548 13828 3560 13880
rect 3612 13828 3624 13880
rect 3548 13756 3624 13828
rect 3548 13704 3560 13756
rect 3612 13704 3624 13756
rect 3548 13632 3624 13704
rect 3548 13580 3560 13632
rect 3612 13580 3624 13632
rect 3548 13508 3624 13580
rect 3548 13456 3560 13508
rect 3612 13456 3624 13508
rect 3548 13384 3624 13456
rect 3548 13332 3560 13384
rect 3612 13332 3624 13384
rect 3548 13260 3624 13332
rect 3548 13208 3560 13260
rect 3612 13208 3624 13260
rect 3548 13136 3624 13208
rect 3548 13084 3560 13136
rect 3612 13084 3624 13136
rect 3548 13012 3624 13084
rect 3548 12960 3560 13012
rect 3612 12960 3624 13012
rect 3548 12932 3624 12960
rect 3996 14996 4072 15008
rect 3996 14944 4008 14996
rect 4060 14944 4072 14996
rect 3996 14872 4072 14944
rect 3996 14820 4008 14872
rect 4060 14820 4072 14872
rect 3996 14748 4072 14820
rect 3996 14696 4008 14748
rect 4060 14696 4072 14748
rect 3996 14624 4072 14696
rect 3996 14572 4008 14624
rect 4060 14572 4072 14624
rect 3996 14500 4072 14572
rect 3996 14448 4008 14500
rect 4060 14448 4072 14500
rect 3996 14376 4072 14448
rect 3996 14324 4008 14376
rect 4060 14324 4072 14376
rect 3996 14252 4072 14324
rect 3996 14200 4008 14252
rect 4060 14200 4072 14252
rect 3996 14128 4072 14200
rect 3996 14076 4008 14128
rect 4060 14076 4072 14128
rect 3996 14004 4072 14076
rect 3996 13952 4008 14004
rect 4060 13952 4072 14004
rect 3996 13880 4072 13952
rect 3996 13828 4008 13880
rect 4060 13828 4072 13880
rect 3996 13756 4072 13828
rect 3996 13704 4008 13756
rect 4060 13704 4072 13756
rect 3996 13632 4072 13704
rect 3996 13580 4008 13632
rect 4060 13580 4072 13632
rect 3996 13508 4072 13580
rect 3996 13456 4008 13508
rect 4060 13456 4072 13508
rect 3996 13384 4072 13456
rect 3996 13332 4008 13384
rect 4060 13332 4072 13384
rect 3996 13260 4072 13332
rect 4668 14996 4744 15008
rect 4668 14944 4680 14996
rect 4732 14944 4744 14996
rect 4668 14872 4744 14944
rect 4668 14820 4680 14872
rect 4732 14820 4744 14872
rect 4668 14748 4744 14820
rect 4668 14696 4680 14748
rect 4732 14696 4744 14748
rect 4668 14624 4744 14696
rect 4668 14572 4680 14624
rect 4732 14572 4744 14624
rect 4668 14500 4744 14572
rect 4668 14448 4680 14500
rect 4732 14448 4744 14500
rect 4668 14376 4744 14448
rect 4668 14324 4680 14376
rect 4732 14324 4744 14376
rect 4668 14252 4744 14324
rect 4668 14200 4680 14252
rect 4732 14200 4744 14252
rect 4668 14128 4744 14200
rect 4668 14076 4680 14128
rect 4732 14076 4744 14128
rect 4668 14004 4744 14076
rect 4668 13952 4680 14004
rect 4732 13952 4744 14004
rect 4668 13880 4744 13952
rect 4668 13828 4680 13880
rect 4732 13828 4744 13880
rect 4668 13756 4744 13828
rect 4668 13704 4680 13756
rect 4732 13704 4744 13756
rect 4668 13632 4744 13704
rect 4668 13580 4680 13632
rect 4732 13580 4744 13632
rect 4668 13508 4744 13580
rect 4668 13456 4680 13508
rect 4732 13456 4744 13508
rect 4668 13384 4744 13456
rect 4668 13332 4680 13384
rect 4732 13332 4744 13384
rect 4668 13272 4744 13332
rect 5116 14996 5192 15008
rect 5116 14944 5128 14996
rect 5180 14944 5192 14996
rect 5116 14872 5192 14944
rect 5116 14820 5128 14872
rect 5180 14820 5192 14872
rect 5116 14748 5192 14820
rect 5116 14696 5128 14748
rect 5180 14696 5192 14748
rect 5116 14624 5192 14696
rect 5116 14572 5128 14624
rect 5180 14572 5192 14624
rect 5116 14500 5192 14572
rect 5116 14448 5128 14500
rect 5180 14448 5192 14500
rect 5116 14376 5192 14448
rect 5116 14324 5128 14376
rect 5180 14324 5192 14376
rect 5116 14252 5192 14324
rect 5116 14200 5128 14252
rect 5180 14200 5192 14252
rect 5116 14128 5192 14200
rect 5116 14076 5128 14128
rect 5180 14076 5192 14128
rect 5116 14004 5192 14076
rect 5116 13952 5128 14004
rect 5180 13952 5192 14004
rect 5116 13880 5192 13952
rect 5116 13828 5128 13880
rect 5180 13828 5192 13880
rect 5116 13756 5192 13828
rect 5116 13704 5128 13756
rect 5180 13704 5192 13756
rect 5116 13632 5192 13704
rect 5116 13580 5128 13632
rect 5180 13580 5192 13632
rect 5788 14996 5864 15008
rect 5788 14944 5800 14996
rect 5852 14944 5864 14996
rect 5788 14872 5864 14944
rect 5788 14820 5800 14872
rect 5852 14820 5864 14872
rect 5788 14748 5864 14820
rect 5788 14696 5800 14748
rect 5852 14696 5864 14748
rect 5788 14624 5864 14696
rect 5788 14572 5800 14624
rect 5852 14572 5864 14624
rect 5788 14500 5864 14572
rect 5788 14448 5800 14500
rect 5852 14448 5864 14500
rect 5788 14376 5864 14448
rect 5788 14324 5800 14376
rect 5852 14324 5864 14376
rect 5788 14252 5864 14324
rect 5788 14200 5800 14252
rect 5852 14200 5864 14252
rect 5788 14128 5864 14200
rect 5788 14076 5800 14128
rect 5852 14076 5864 14128
rect 5788 14004 5864 14076
rect 5788 13952 5800 14004
rect 5852 13952 5864 14004
rect 5788 13880 5864 13952
rect 5788 13828 5800 13880
rect 5852 13828 5864 13880
rect 5788 13756 5864 13828
rect 5788 13704 5800 13756
rect 5852 13704 5864 13756
rect 5788 13632 5864 13704
rect 5788 13612 5800 13632
rect 5116 13508 5192 13580
rect 5116 13456 5128 13508
rect 5180 13456 5192 13508
rect 5761 13580 5800 13612
rect 5852 13612 5864 13632
rect 6236 14996 6312 15008
rect 6236 14944 6248 14996
rect 6300 14944 6312 14996
rect 6236 14872 6312 14944
rect 6236 14820 6248 14872
rect 6300 14820 6312 14872
rect 6236 14748 6312 14820
rect 6236 14696 6248 14748
rect 6300 14696 6312 14748
rect 6236 14624 6312 14696
rect 6236 14572 6248 14624
rect 6300 14572 6312 14624
rect 6236 14500 6312 14572
rect 6236 14448 6248 14500
rect 6300 14448 6312 14500
rect 6236 14376 6312 14448
rect 6236 14324 6248 14376
rect 6300 14324 6312 14376
rect 6236 14252 6312 14324
rect 6236 14200 6248 14252
rect 6300 14200 6312 14252
rect 6236 14128 6312 14200
rect 6236 14076 6248 14128
rect 6300 14076 6312 14128
rect 6236 14004 6312 14076
rect 6236 13952 6248 14004
rect 6300 13952 6312 14004
rect 6908 14996 6984 15008
rect 6908 14944 6920 14996
rect 6972 14944 6984 14996
rect 6908 14872 6984 14944
rect 6908 14820 6920 14872
rect 6972 14820 6984 14872
rect 6908 14748 6984 14820
rect 6908 14696 6920 14748
rect 6972 14696 6984 14748
rect 6908 14624 6984 14696
rect 6908 14572 6920 14624
rect 6972 14572 6984 14624
rect 6908 14500 6984 14572
rect 6908 14448 6920 14500
rect 6972 14448 6984 14500
rect 6908 14376 6984 14448
rect 6908 14324 6920 14376
rect 6972 14324 6984 14376
rect 6908 14252 6984 14324
rect 6908 14200 6920 14252
rect 6972 14200 6984 14252
rect 6908 14128 6984 14200
rect 6908 14076 6920 14128
rect 6972 14076 6984 14128
rect 6908 14004 6984 14076
rect 6908 13952 6920 14004
rect 6972 13952 6984 14004
rect 7356 14996 7432 15008
rect 7356 14944 7368 14996
rect 7420 14944 7432 14996
rect 7356 14872 7432 14944
rect 7356 14820 7368 14872
rect 7420 14820 7432 14872
rect 7356 14748 7432 14820
rect 7356 14696 7368 14748
rect 7420 14696 7432 14748
rect 7356 14624 7432 14696
rect 7356 14572 7368 14624
rect 7420 14572 7432 14624
rect 7356 14500 7432 14572
rect 7356 14448 7368 14500
rect 7420 14448 7432 14500
rect 7356 14376 7432 14448
rect 7356 14324 7368 14376
rect 7420 14324 7432 14376
rect 7356 14252 7432 14324
rect 8028 14996 8104 15008
rect 8028 14944 8040 14996
rect 8092 14944 8104 14996
rect 8028 14872 8104 14944
rect 8028 14820 8040 14872
rect 8092 14820 8104 14872
rect 8028 14748 8104 14820
rect 8028 14696 8040 14748
rect 8092 14696 8104 14748
rect 8028 14624 8104 14696
rect 8028 14572 8040 14624
rect 8092 14572 8104 14624
rect 8028 14500 8104 14572
rect 8028 14448 8040 14500
rect 8092 14448 8104 14500
rect 8028 14376 8104 14448
rect 8028 14324 8040 14376
rect 8092 14324 8104 14376
rect 8028 14292 8104 14324
rect 8476 14996 8552 15008
rect 8476 14944 8488 14996
rect 8540 14944 8552 14996
rect 8476 14872 8552 14944
rect 8476 14820 8488 14872
rect 8540 14820 8552 14872
rect 8476 14748 8552 14820
rect 8476 14696 8488 14748
rect 8540 14696 8552 14748
rect 8476 14624 8552 14696
rect 9148 14996 9224 15008
rect 9148 14944 9160 14996
rect 9212 14944 9224 14996
rect 9148 14872 9224 14944
rect 9148 14820 9160 14872
rect 9212 14820 9224 14872
rect 9148 14748 9224 14820
rect 9148 14696 9160 14748
rect 9212 14696 9224 14748
rect 9148 14633 9224 14696
rect 9596 14996 9672 15008
rect 9596 14944 9608 14996
rect 9660 14944 9672 14996
rect 10268 14996 10344 15008
rect 10268 14973 10280 14996
rect 9596 14872 9672 14944
rect 9596 14820 9608 14872
rect 9660 14820 9672 14872
rect 10240 14944 10280 14973
rect 10332 14973 10344 14996
rect 10716 14996 10792 15008
rect 10716 14973 10728 14996
rect 10332 14944 10369 14973
rect 10240 14934 10369 14944
rect 10240 14878 10277 14934
rect 10333 14878 10369 14934
rect 10240 14872 10369 14878
rect 10240 14839 10280 14872
rect 9596 14748 9672 14820
rect 9596 14696 9608 14748
rect 9660 14696 9672 14748
rect 9596 14633 9672 14696
rect 10268 14820 10280 14839
rect 10332 14839 10369 14872
rect 10688 14944 10728 14973
rect 10780 14973 10792 14996
rect 11388 14996 11464 15008
rect 10780 14944 10817 14973
rect 10688 14934 10817 14944
rect 10688 14878 10725 14934
rect 10781 14878 10817 14934
rect 10688 14872 10817 14878
rect 10688 14839 10728 14872
rect 10332 14820 10344 14839
rect 10268 14748 10344 14820
rect 10268 14696 10280 14748
rect 10332 14696 10344 14748
rect 8476 14572 8488 14624
rect 8540 14572 8552 14624
rect 8476 14500 8552 14572
rect 8476 14448 8488 14500
rect 8540 14448 8552 14500
rect 9121 14624 9250 14633
rect 9121 14594 9160 14624
rect 9212 14594 9250 14624
rect 9121 14538 9158 14594
rect 9214 14538 9250 14594
rect 9121 14500 9250 14538
rect 9121 14499 9160 14500
rect 8476 14376 8552 14448
rect 8476 14324 8488 14376
rect 8540 14324 8552 14376
rect 8476 14292 8552 14324
rect 9148 14448 9160 14499
rect 9212 14499 9250 14500
rect 9568 14624 9697 14633
rect 9568 14594 9608 14624
rect 9660 14594 9697 14624
rect 9568 14538 9605 14594
rect 9661 14538 9697 14594
rect 9568 14500 9697 14538
rect 9568 14499 9608 14500
rect 9212 14448 9224 14499
rect 9148 14376 9224 14448
rect 9148 14324 9160 14376
rect 9212 14324 9224 14376
rect 7356 14200 7368 14252
rect 7420 14200 7432 14252
rect 7356 14128 7432 14200
rect 8001 14253 8130 14292
rect 8001 14197 8038 14253
rect 8094 14197 8130 14253
rect 8001 14158 8130 14197
rect 8449 14253 8578 14292
rect 8449 14197 8486 14253
rect 8542 14197 8578 14253
rect 8449 14158 8578 14197
rect 9148 14252 9224 14324
rect 9148 14200 9160 14252
rect 9212 14200 9224 14252
rect 7356 14076 7368 14128
rect 7420 14076 7432 14128
rect 7356 14004 7432 14076
rect 7356 13952 7368 14004
rect 7420 13952 7432 14004
rect 8028 14128 8104 14158
rect 8028 14076 8040 14128
rect 8092 14076 8104 14128
rect 8028 14004 8104 14076
rect 8028 13952 8040 14004
rect 8092 13952 8104 14004
rect 6236 13880 6312 13952
rect 6236 13828 6248 13880
rect 6300 13828 6312 13880
rect 6236 13756 6312 13828
rect 6881 13913 7010 13952
rect 6881 13857 6918 13913
rect 6974 13857 7010 13913
rect 6881 13828 6920 13857
rect 6972 13828 7010 13857
rect 6881 13818 7010 13828
rect 7329 13913 7458 13952
rect 7329 13857 7366 13913
rect 7422 13857 7458 13913
rect 7329 13828 7368 13857
rect 7420 13828 7458 13857
rect 7329 13818 7458 13828
rect 8028 13880 8104 13952
rect 8028 13828 8040 13880
rect 8092 13828 8104 13880
rect 6236 13704 6248 13756
rect 6300 13704 6312 13756
rect 6236 13632 6312 13704
rect 6236 13612 6248 13632
rect 5852 13580 5890 13612
rect 5761 13573 5890 13580
rect 5761 13517 5798 13573
rect 5854 13517 5890 13573
rect 5761 13508 5890 13517
rect 5761 13478 5800 13508
rect 5116 13384 5192 13456
rect 5116 13332 5128 13384
rect 5180 13332 5192 13384
rect 5116 13272 5192 13332
rect 5788 13456 5800 13478
rect 5852 13478 5890 13508
rect 6209 13580 6248 13612
rect 6300 13612 6312 13632
rect 6908 13756 6984 13818
rect 6908 13704 6920 13756
rect 6972 13704 6984 13756
rect 6908 13632 6984 13704
rect 6300 13580 6338 13612
rect 6209 13573 6338 13580
rect 6209 13517 6246 13573
rect 6302 13517 6338 13573
rect 6209 13508 6338 13517
rect 6209 13478 6248 13508
rect 5852 13456 5864 13478
rect 5788 13384 5864 13456
rect 5788 13332 5800 13384
rect 5852 13332 5864 13384
rect 3996 13208 4008 13260
rect 4060 13208 4072 13260
rect 3996 13136 4072 13208
rect 4641 13260 4770 13272
rect 4641 13233 4680 13260
rect 4732 13233 4770 13260
rect 4641 13177 4678 13233
rect 4734 13177 4770 13233
rect 4641 13138 4770 13177
rect 5089 13260 5218 13272
rect 5089 13233 5128 13260
rect 5180 13233 5218 13260
rect 5089 13177 5126 13233
rect 5182 13177 5218 13233
rect 5089 13138 5218 13177
rect 5788 13260 5864 13332
rect 5788 13208 5800 13260
rect 5852 13208 5864 13260
rect 3996 13084 4008 13136
rect 4060 13084 4072 13136
rect 3996 13012 4072 13084
rect 3996 12960 4008 13012
rect 4060 12960 4072 13012
rect 3996 12932 4072 12960
rect 4668 13136 4744 13138
rect 4668 13084 4680 13136
rect 4732 13084 4744 13136
rect 4668 13012 4744 13084
rect 4668 12960 4680 13012
rect 4732 12960 4744 13012
rect 2876 12836 2888 12888
rect 2940 12836 2952 12888
rect 2876 12592 2952 12836
rect 3521 12893 3650 12932
rect 3521 12837 3558 12893
rect 3614 12837 3650 12893
rect 3521 12836 3560 12837
rect 3612 12836 3650 12837
rect 3521 12798 3650 12836
rect 3969 12893 4098 12932
rect 3969 12837 4006 12893
rect 4062 12837 4098 12893
rect 3969 12836 4008 12837
rect 4060 12836 4098 12837
rect 3969 12798 4098 12836
rect 4668 12888 4744 12960
rect 4668 12836 4680 12888
rect 4732 12836 4744 12888
rect 2401 12553 2530 12592
rect 2401 12497 2438 12553
rect 2494 12497 2530 12553
rect 2401 12458 2530 12497
rect 2849 12553 2978 12592
rect 2849 12497 2886 12553
rect 2942 12497 2978 12553
rect 2849 12458 2978 12497
rect 1970 12152 2095 12191
rect 1970 12096 2005 12152
rect 2061 12096 2095 12152
rect 1970 11934 2095 12096
rect 1970 11878 2005 11934
rect 2061 11878 2095 11934
rect 1970 11859 2008 11878
rect 2060 11859 2095 11878
rect 1970 11840 2095 11859
rect 2428 11758 2504 12458
rect 2428 11706 2440 11758
rect 2492 11706 2504 11758
rect 2428 11634 2504 11706
rect 2428 11582 2440 11634
rect 2492 11582 2504 11634
rect 2428 11510 2504 11582
rect 2428 11458 2440 11510
rect 2492 11458 2504 11510
rect 2428 11446 2504 11458
rect 2876 11758 2952 12458
rect 3116 11911 3192 12009
rect 3116 11889 3128 11911
rect 2876 11706 2888 11758
rect 2940 11706 2952 11758
rect 3089 11859 3128 11889
rect 3180 11889 3192 11911
rect 3180 11859 3429 11889
rect 3089 11850 3429 11859
rect 3089 11794 3125 11850
rect 3181 11794 3337 11850
rect 3393 11794 3429 11850
rect 3089 11755 3429 11794
rect 3548 11758 3624 12798
rect 2876 11634 2952 11706
rect 2876 11582 2888 11634
rect 2940 11582 2952 11634
rect 2876 11510 2952 11582
rect 2876 11458 2888 11510
rect 2940 11458 2952 11510
rect 2876 11446 2952 11458
rect 3548 11706 3560 11758
rect 3612 11706 3624 11758
rect 3548 11634 3624 11706
rect 3548 11582 3560 11634
rect 3612 11582 3624 11634
rect 3548 11510 3624 11582
rect 3548 11458 3560 11510
rect 3612 11458 3624 11510
rect 3548 11446 3624 11458
rect 3996 11758 4072 12798
rect 4236 11973 4312 12009
rect 3996 11706 4008 11758
rect 4060 11706 4072 11758
rect 3996 11634 4072 11706
rect 3996 11582 4008 11634
rect 4060 11582 4072 11634
rect 3996 11510 4072 11582
rect 4209 11911 4338 11973
rect 4209 11859 4248 11911
rect 4300 11859 4338 11911
rect 4209 11622 4338 11859
rect 4209 11568 4245 11622
rect 3996 11458 4008 11510
rect 4060 11458 4072 11510
rect 3996 11446 4072 11458
rect 4210 11566 4245 11568
rect 4301 11568 4338 11622
rect 4668 11758 4744 12836
rect 4668 11706 4680 11758
rect 4732 11706 4744 11758
rect 4668 11634 4744 11706
rect 4668 11582 4680 11634
rect 4732 11582 4744 11634
rect 4301 11566 4335 11568
rect 4210 11404 4335 11566
rect 4668 11510 4744 11582
rect 4668 11458 4680 11510
rect 4732 11458 4744 11510
rect 4668 11446 4744 11458
rect 5116 13136 5192 13138
rect 5116 13084 5128 13136
rect 5180 13084 5192 13136
rect 5116 13012 5192 13084
rect 5116 12960 5128 13012
rect 5180 12960 5192 13012
rect 5116 12888 5192 12960
rect 5116 12836 5128 12888
rect 5180 12836 5192 12888
rect 5116 11758 5192 12836
rect 5788 13136 5864 13208
rect 5788 13084 5800 13136
rect 5852 13084 5864 13136
rect 5788 13012 5864 13084
rect 5788 12960 5800 13012
rect 5852 12960 5864 13012
rect 5788 12888 5864 12960
rect 5788 12836 5800 12888
rect 5852 12836 5864 12888
rect 5356 11973 5432 12009
rect 5116 11706 5128 11758
rect 5180 11706 5192 11758
rect 5116 11634 5192 11706
rect 5116 11582 5128 11634
rect 5180 11582 5192 11634
rect 5116 11510 5192 11582
rect 5116 11458 5128 11510
rect 5180 11458 5192 11510
rect 5329 11911 5458 11973
rect 5329 11859 5368 11911
rect 5420 11859 5458 11911
rect 5329 11472 5458 11859
rect 5788 11758 5864 12836
rect 5788 11706 5800 11758
rect 5852 11706 5864 11758
rect 5788 11634 5864 11706
rect 5788 11582 5800 11634
rect 5852 11582 5864 11634
rect 5788 11510 5864 11582
rect 5116 11446 5192 11458
rect 4210 11348 4245 11404
rect 4301 11348 4335 11404
rect 4210 11310 4335 11348
rect 5328 11433 5668 11472
rect 5788 11458 5800 11510
rect 5852 11458 5864 11510
rect 5788 11446 5864 11458
rect 6236 13456 6248 13478
rect 6300 13478 6338 13508
rect 6908 13580 6920 13632
rect 6972 13580 6984 13632
rect 6908 13508 6984 13580
rect 6300 13456 6312 13478
rect 6236 13384 6312 13456
rect 6236 13332 6248 13384
rect 6300 13332 6312 13384
rect 6236 13260 6312 13332
rect 6236 13208 6248 13260
rect 6300 13208 6312 13260
rect 6236 13136 6312 13208
rect 6236 13084 6248 13136
rect 6300 13084 6312 13136
rect 6236 13012 6312 13084
rect 6236 12960 6248 13012
rect 6300 12960 6312 13012
rect 6236 12888 6312 12960
rect 6236 12836 6248 12888
rect 6300 12836 6312 12888
rect 6236 11758 6312 12836
rect 6908 13456 6920 13508
rect 6972 13456 6984 13508
rect 6908 13384 6984 13456
rect 6908 13332 6920 13384
rect 6972 13332 6984 13384
rect 6908 13260 6984 13332
rect 6908 13208 6920 13260
rect 6972 13208 6984 13260
rect 6908 13136 6984 13208
rect 6908 13084 6920 13136
rect 6972 13084 6984 13136
rect 6908 13012 6984 13084
rect 6908 12960 6920 13012
rect 6972 12960 6984 13012
rect 6908 12888 6984 12960
rect 6908 12836 6920 12888
rect 6972 12836 6984 12888
rect 6476 11973 6552 12009
rect 6236 11706 6248 11758
rect 6300 11706 6312 11758
rect 6236 11634 6312 11706
rect 6236 11582 6248 11634
rect 6300 11582 6312 11634
rect 6236 11510 6312 11582
rect 6236 11458 6248 11510
rect 6300 11458 6312 11510
rect 6236 11446 6312 11458
rect 6449 11911 6578 11973
rect 6449 11859 6488 11911
rect 6540 11859 6578 11911
rect 5328 11377 5364 11433
rect 5420 11377 5576 11433
rect 5632 11377 5668 11433
rect 5328 11338 5668 11377
rect 6449 11264 6578 11859
rect 6908 11758 6984 12836
rect 6908 11706 6920 11758
rect 6972 11706 6984 11758
rect 6908 11634 6984 11706
rect 6908 11582 6920 11634
rect 6972 11582 6984 11634
rect 6908 11510 6984 11582
rect 6908 11458 6920 11510
rect 6972 11458 6984 11510
rect 6908 11446 6984 11458
rect 7356 13756 7432 13818
rect 7356 13704 7368 13756
rect 7420 13704 7432 13756
rect 7356 13632 7432 13704
rect 7356 13580 7368 13632
rect 7420 13580 7432 13632
rect 7356 13508 7432 13580
rect 7356 13456 7368 13508
rect 7420 13456 7432 13508
rect 7356 13384 7432 13456
rect 7356 13332 7368 13384
rect 7420 13332 7432 13384
rect 7356 13260 7432 13332
rect 7356 13208 7368 13260
rect 7420 13208 7432 13260
rect 7356 13136 7432 13208
rect 7356 13084 7368 13136
rect 7420 13084 7432 13136
rect 7356 13012 7432 13084
rect 7356 12960 7368 13012
rect 7420 12960 7432 13012
rect 7356 12888 7432 12960
rect 7356 12836 7368 12888
rect 7420 12836 7432 12888
rect 7356 11758 7432 12836
rect 8028 13756 8104 13828
rect 8028 13704 8040 13756
rect 8092 13704 8104 13756
rect 8028 13632 8104 13704
rect 8028 13580 8040 13632
rect 8092 13580 8104 13632
rect 8028 13508 8104 13580
rect 8028 13456 8040 13508
rect 8092 13456 8104 13508
rect 8028 13384 8104 13456
rect 8028 13332 8040 13384
rect 8092 13332 8104 13384
rect 8028 13260 8104 13332
rect 8028 13208 8040 13260
rect 8092 13208 8104 13260
rect 8028 13136 8104 13208
rect 8028 13084 8040 13136
rect 8092 13084 8104 13136
rect 8028 13012 8104 13084
rect 8028 12960 8040 13012
rect 8092 12960 8104 13012
rect 8028 12888 8104 12960
rect 8028 12836 8040 12888
rect 8092 12836 8104 12888
rect 7596 11973 7672 12009
rect 7356 11706 7368 11758
rect 7420 11706 7432 11758
rect 7356 11634 7432 11706
rect 7356 11582 7368 11634
rect 7420 11582 7432 11634
rect 7356 11510 7432 11582
rect 7356 11458 7368 11510
rect 7420 11458 7432 11510
rect 7356 11446 7432 11458
rect 7569 11911 7698 11973
rect 7569 11859 7608 11911
rect 7660 11859 7698 11911
rect 6343 11225 6683 11264
rect 6343 11169 6379 11225
rect 6435 11169 6591 11225
rect 6647 11169 6683 11225
rect 6343 11130 6683 11169
rect 7569 11055 7698 11859
rect 8028 11758 8104 12836
rect 8028 11706 8040 11758
rect 8092 11706 8104 11758
rect 8028 11634 8104 11706
rect 8028 11582 8040 11634
rect 8092 11582 8104 11634
rect 8028 11510 8104 11582
rect 8028 11458 8040 11510
rect 8092 11458 8104 11510
rect 8028 11446 8104 11458
rect 8476 14128 8552 14158
rect 8476 14076 8488 14128
rect 8540 14076 8552 14128
rect 8476 14004 8552 14076
rect 8476 13952 8488 14004
rect 8540 13952 8552 14004
rect 8476 13880 8552 13952
rect 8476 13828 8488 13880
rect 8540 13828 8552 13880
rect 8476 13756 8552 13828
rect 8476 13704 8488 13756
rect 8540 13704 8552 13756
rect 8476 13632 8552 13704
rect 8476 13580 8488 13632
rect 8540 13580 8552 13632
rect 8476 13508 8552 13580
rect 8476 13456 8488 13508
rect 8540 13456 8552 13508
rect 8476 13384 8552 13456
rect 8476 13332 8488 13384
rect 8540 13332 8552 13384
rect 8476 13260 8552 13332
rect 8476 13208 8488 13260
rect 8540 13208 8552 13260
rect 8476 13136 8552 13208
rect 8476 13084 8488 13136
rect 8540 13084 8552 13136
rect 8476 13012 8552 13084
rect 8476 12960 8488 13012
rect 8540 12960 8552 13012
rect 8476 12888 8552 12960
rect 8476 12836 8488 12888
rect 8540 12836 8552 12888
rect 8476 11758 8552 12836
rect 9148 14128 9224 14200
rect 9148 14076 9160 14128
rect 9212 14076 9224 14128
rect 9148 14004 9224 14076
rect 9148 13952 9160 14004
rect 9212 13952 9224 14004
rect 9148 13880 9224 13952
rect 9148 13828 9160 13880
rect 9212 13828 9224 13880
rect 9148 13756 9224 13828
rect 9148 13704 9160 13756
rect 9212 13704 9224 13756
rect 9148 13632 9224 13704
rect 9148 13580 9160 13632
rect 9212 13580 9224 13632
rect 9148 13508 9224 13580
rect 9148 13456 9160 13508
rect 9212 13456 9224 13508
rect 9148 13384 9224 13456
rect 9148 13332 9160 13384
rect 9212 13332 9224 13384
rect 9148 13260 9224 13332
rect 9148 13208 9160 13260
rect 9212 13208 9224 13260
rect 9148 13136 9224 13208
rect 9148 13084 9160 13136
rect 9212 13084 9224 13136
rect 9148 13012 9224 13084
rect 9148 12960 9160 13012
rect 9212 12960 9224 13012
rect 9148 12888 9224 12960
rect 9148 12836 9160 12888
rect 9212 12836 9224 12888
rect 8716 11973 8792 12009
rect 8476 11706 8488 11758
rect 8540 11706 8552 11758
rect 8476 11634 8552 11706
rect 8476 11582 8488 11634
rect 8540 11582 8552 11634
rect 8476 11510 8552 11582
rect 8476 11458 8488 11510
rect 8540 11458 8552 11510
rect 8476 11446 8552 11458
rect 8689 11911 8818 11973
rect 8689 11859 8728 11911
rect 8780 11859 8818 11911
rect 7463 11016 7803 11055
rect 7463 10960 7499 11016
rect 7555 10960 7711 11016
rect 7767 10960 7803 11016
rect 7463 10921 7803 10960
rect 8689 10847 8818 11859
rect 9148 11758 9224 12836
rect 9148 11706 9160 11758
rect 9212 11706 9224 11758
rect 9148 11634 9224 11706
rect 9148 11582 9160 11634
rect 9212 11582 9224 11634
rect 9148 11510 9224 11582
rect 9148 11458 9160 11510
rect 9212 11458 9224 11510
rect 9148 11446 9224 11458
rect 9596 14448 9608 14499
rect 9660 14499 9697 14500
rect 10268 14624 10344 14696
rect 10268 14572 10280 14624
rect 10332 14572 10344 14624
rect 10268 14500 10344 14572
rect 9660 14448 9672 14499
rect 9596 14376 9672 14448
rect 9596 14324 9608 14376
rect 9660 14324 9672 14376
rect 9596 14252 9672 14324
rect 9596 14200 9608 14252
rect 9660 14200 9672 14252
rect 9596 14128 9672 14200
rect 9596 14076 9608 14128
rect 9660 14076 9672 14128
rect 9596 14004 9672 14076
rect 9596 13952 9608 14004
rect 9660 13952 9672 14004
rect 9596 13880 9672 13952
rect 9596 13828 9608 13880
rect 9660 13828 9672 13880
rect 9596 13756 9672 13828
rect 9596 13704 9608 13756
rect 9660 13704 9672 13756
rect 9596 13632 9672 13704
rect 9596 13580 9608 13632
rect 9660 13580 9672 13632
rect 9596 13508 9672 13580
rect 9596 13456 9608 13508
rect 9660 13456 9672 13508
rect 9596 13384 9672 13456
rect 9596 13332 9608 13384
rect 9660 13332 9672 13384
rect 9596 13260 9672 13332
rect 9596 13208 9608 13260
rect 9660 13208 9672 13260
rect 9596 13136 9672 13208
rect 9596 13084 9608 13136
rect 9660 13084 9672 13136
rect 9596 13012 9672 13084
rect 9596 12960 9608 13012
rect 9660 12960 9672 13012
rect 9596 12888 9672 12960
rect 9596 12836 9608 12888
rect 9660 12836 9672 12888
rect 9596 11758 9672 12836
rect 10268 14448 10280 14500
rect 10332 14448 10344 14500
rect 10268 14376 10344 14448
rect 10268 14324 10280 14376
rect 10332 14324 10344 14376
rect 10268 14252 10344 14324
rect 10268 14200 10280 14252
rect 10332 14200 10344 14252
rect 10268 14128 10344 14200
rect 10268 14076 10280 14128
rect 10332 14076 10344 14128
rect 10268 14004 10344 14076
rect 10268 13952 10280 14004
rect 10332 13952 10344 14004
rect 10268 13880 10344 13952
rect 10268 13828 10280 13880
rect 10332 13828 10344 13880
rect 10268 13756 10344 13828
rect 10268 13704 10280 13756
rect 10332 13704 10344 13756
rect 10268 13632 10344 13704
rect 10268 13580 10280 13632
rect 10332 13580 10344 13632
rect 10268 13508 10344 13580
rect 10268 13456 10280 13508
rect 10332 13456 10344 13508
rect 10268 13384 10344 13456
rect 10268 13332 10280 13384
rect 10332 13332 10344 13384
rect 10268 13260 10344 13332
rect 10268 13208 10280 13260
rect 10332 13208 10344 13260
rect 10268 13136 10344 13208
rect 10268 13084 10280 13136
rect 10332 13084 10344 13136
rect 10268 13012 10344 13084
rect 10268 12960 10280 13012
rect 10332 12960 10344 13012
rect 10268 12888 10344 12960
rect 10268 12836 10280 12888
rect 10332 12836 10344 12888
rect 9836 11973 9912 12009
rect 9596 11706 9608 11758
rect 9660 11706 9672 11758
rect 9596 11634 9672 11706
rect 9596 11582 9608 11634
rect 9660 11582 9672 11634
rect 9596 11510 9672 11582
rect 9596 11458 9608 11510
rect 9660 11458 9672 11510
rect 9596 11446 9672 11458
rect 9809 11911 9938 11973
rect 9809 11859 9848 11911
rect 9900 11859 9938 11911
rect 9281 11016 9621 11055
rect 9281 10960 9317 11016
rect 9373 10960 9529 11016
rect 9585 10960 9621 11016
rect 9281 10921 9621 10960
rect 8390 10846 8818 10847
rect 8302 10808 8818 10846
rect 8302 10752 8426 10808
rect 8482 10752 8638 10808
rect 8694 10752 8818 10808
rect 8302 10713 8818 10752
rect 7753 10599 8093 10638
rect 7753 10543 7789 10599
rect 7845 10543 8001 10599
rect 8057 10543 8093 10599
rect 7753 10504 8093 10543
rect 2366 9366 2701 9405
rect 2366 9310 2402 9366
rect 2458 9310 2609 9366
rect 2665 9310 2701 9366
rect 2366 9148 2701 9310
rect 2366 9092 2402 9148
rect 2458 9092 2609 9148
rect 2665 9092 2701 9148
rect 2366 8930 2701 9092
rect 2366 8874 2402 8930
rect 2458 8874 2609 8930
rect 2665 8874 2701 8930
rect 2366 8712 2701 8874
rect 2366 8656 2402 8712
rect 2458 8656 2609 8712
rect 2665 8656 2701 8712
rect 2366 8618 2701 8656
rect 3093 9366 3221 9403
rect 3093 9310 3129 9366
rect 3185 9310 3221 9366
rect 3093 9148 3221 9310
rect 3093 9092 3129 9148
rect 3185 9092 3221 9148
rect 3093 8930 3221 9092
rect 3093 8874 3129 8930
rect 3185 8874 3221 8930
rect 3093 8712 3221 8874
rect 3093 8656 3129 8712
rect 3185 8656 3221 8712
rect 3093 8618 3221 8656
rect 4057 9366 4392 9405
rect 4057 9310 4093 9366
rect 4149 9310 4300 9366
rect 4356 9310 4392 9366
rect 4057 9148 4392 9310
rect 4057 9092 4093 9148
rect 4149 9092 4300 9148
rect 4356 9092 4392 9148
rect 4057 8930 4392 9092
rect 4057 8874 4093 8930
rect 4149 8874 4300 8930
rect 4356 8874 4392 8930
rect 4057 8712 4392 8874
rect 4057 8656 4093 8712
rect 4149 8656 4300 8712
rect 4356 8656 4392 8712
rect 4057 8618 4392 8656
rect 4784 9366 4912 9403
rect 4784 9310 4820 9366
rect 4876 9310 4912 9366
rect 4784 9148 4912 9310
rect 4784 9092 4820 9148
rect 4876 9092 4912 9148
rect 4784 8930 4912 9092
rect 4784 8874 4820 8930
rect 4876 8874 4912 8930
rect 4784 8712 4912 8874
rect 4784 8656 4820 8712
rect 4876 8656 4912 8712
rect 4784 8618 4912 8656
rect 5748 9366 6083 9405
rect 5748 9310 5784 9366
rect 5840 9310 5991 9366
rect 6047 9310 6083 9366
rect 5748 9148 6083 9310
rect 5748 9092 5784 9148
rect 5840 9092 5991 9148
rect 6047 9092 6083 9148
rect 5748 8930 6083 9092
rect 5748 8874 5784 8930
rect 5840 8874 5991 8930
rect 6047 8874 6083 8930
rect 5748 8712 6083 8874
rect 5748 8656 5784 8712
rect 5840 8656 5991 8712
rect 6047 8656 6083 8712
rect 5748 8618 6083 8656
rect 6475 9366 6603 9403
rect 6475 9310 6511 9366
rect 6567 9310 6603 9366
rect 6475 9148 6603 9310
rect 6475 9092 6511 9148
rect 6567 9092 6603 9148
rect 6475 8930 6603 9092
rect 6475 8874 6511 8930
rect 6567 8874 6603 8930
rect 6475 8712 6603 8874
rect 6475 8656 6511 8712
rect 6567 8656 6603 8712
rect 6475 8618 6603 8656
rect 7633 9326 7761 9363
rect 7633 9270 7669 9326
rect 7725 9270 7761 9326
rect 7858 9287 7987 10504
rect 7633 9108 7761 9270
rect 7633 9052 7669 9108
rect 7725 9052 7761 9108
rect 7633 8890 7761 9052
rect 7633 8834 7669 8890
rect 7725 8834 7761 8890
rect 7633 8672 7761 8834
rect 7633 8616 7669 8672
rect 7725 8616 7761 8672
rect 7633 8578 7761 8616
rect 7859 8973 7987 9287
rect 7859 8921 7897 8973
rect 7949 8921 7987 8973
rect 7859 8755 7987 8921
rect 7859 8703 7897 8755
rect 7949 8703 7987 8755
rect 7859 8537 7987 8703
rect 8081 9326 8209 9363
rect 8081 9270 8117 9326
rect 8173 9270 8209 9326
rect 8302 9287 8431 10713
rect 8081 9108 8209 9270
rect 8081 9052 8117 9108
rect 8173 9052 8209 9108
rect 8081 8890 8209 9052
rect 8081 8834 8117 8890
rect 8173 8834 8209 8890
rect 8081 8672 8209 8834
rect 8081 8616 8117 8672
rect 8173 8616 8209 8672
rect 8081 8578 8209 8616
rect 8303 8973 8431 9287
rect 8303 8921 8341 8973
rect 8393 8921 8431 8973
rect 8303 8755 8431 8921
rect 8303 8703 8341 8755
rect 8393 8703 8431 8755
rect 7859 8485 7897 8537
rect 7949 8485 7987 8537
rect 7859 8445 7987 8485
rect 8303 8537 8431 8703
rect 8529 9326 8657 9363
rect 8529 9270 8565 9326
rect 8621 9270 8657 9326
rect 8529 9108 8657 9270
rect 8529 9052 8565 9108
rect 8621 9052 8657 9108
rect 8529 8890 8657 9052
rect 8529 8834 8565 8890
rect 8621 8834 8657 8890
rect 8529 8672 8657 8834
rect 8529 8616 8565 8672
rect 8621 8616 8657 8672
rect 8529 8578 8657 8616
rect 9266 9326 9394 9363
rect 9266 9270 9302 9326
rect 9358 9270 9394 9326
rect 9266 9108 9394 9270
rect 9266 9052 9302 9108
rect 9358 9052 9394 9108
rect 9266 8890 9394 9052
rect 9266 8834 9302 8890
rect 9358 8834 9394 8890
rect 9266 8672 9394 8834
rect 9266 8616 9302 8672
rect 9358 8616 9394 8672
rect 9266 8578 9394 8616
rect 9492 9287 9621 10921
rect 9809 10638 9938 11859
rect 10268 11758 10344 12836
rect 10268 11706 10280 11758
rect 10332 11706 10344 11758
rect 10268 11634 10344 11706
rect 10268 11582 10280 11634
rect 10332 11582 10344 11634
rect 10268 11510 10344 11582
rect 10268 11458 10280 11510
rect 10332 11458 10344 11510
rect 10268 11446 10344 11458
rect 10716 14820 10728 14839
rect 10780 14839 10817 14872
rect 11388 14944 11400 14996
rect 11452 14944 11464 14996
rect 11388 14872 11464 14944
rect 10780 14820 10792 14839
rect 10716 14748 10792 14820
rect 10716 14696 10728 14748
rect 10780 14696 10792 14748
rect 10716 14624 10792 14696
rect 10716 14572 10728 14624
rect 10780 14572 10792 14624
rect 10716 14500 10792 14572
rect 10716 14448 10728 14500
rect 10780 14448 10792 14500
rect 10716 14376 10792 14448
rect 10716 14324 10728 14376
rect 10780 14324 10792 14376
rect 10716 14252 10792 14324
rect 10716 14200 10728 14252
rect 10780 14200 10792 14252
rect 10716 14128 10792 14200
rect 10716 14076 10728 14128
rect 10780 14076 10792 14128
rect 10716 14004 10792 14076
rect 10716 13952 10728 14004
rect 10780 13952 10792 14004
rect 10716 13880 10792 13952
rect 10716 13828 10728 13880
rect 10780 13828 10792 13880
rect 10716 13756 10792 13828
rect 10716 13704 10728 13756
rect 10780 13704 10792 13756
rect 10716 13632 10792 13704
rect 10716 13580 10728 13632
rect 10780 13580 10792 13632
rect 10716 13508 10792 13580
rect 10716 13456 10728 13508
rect 10780 13456 10792 13508
rect 10716 13384 10792 13456
rect 10716 13332 10728 13384
rect 10780 13332 10792 13384
rect 10716 13260 10792 13332
rect 10716 13208 10728 13260
rect 10780 13208 10792 13260
rect 10716 13136 10792 13208
rect 10716 13084 10728 13136
rect 10780 13084 10792 13136
rect 10716 13012 10792 13084
rect 10716 12960 10728 13012
rect 10780 12960 10792 13012
rect 10716 12888 10792 12960
rect 10716 12836 10728 12888
rect 10780 12836 10792 12888
rect 10716 11758 10792 12836
rect 11388 14820 11400 14872
rect 11452 14820 11464 14872
rect 11388 14748 11464 14820
rect 11388 14696 11400 14748
rect 11452 14696 11464 14748
rect 11388 14624 11464 14696
rect 11388 14572 11400 14624
rect 11452 14572 11464 14624
rect 11388 14500 11464 14572
rect 11388 14448 11400 14500
rect 11452 14448 11464 14500
rect 11388 14376 11464 14448
rect 11388 14324 11400 14376
rect 11452 14324 11464 14376
rect 11388 14252 11464 14324
rect 11388 14200 11400 14252
rect 11452 14200 11464 14252
rect 11388 14128 11464 14200
rect 11388 14076 11400 14128
rect 11452 14076 11464 14128
rect 11388 14004 11464 14076
rect 11388 13952 11400 14004
rect 11452 13952 11464 14004
rect 11388 13880 11464 13952
rect 11388 13828 11400 13880
rect 11452 13828 11464 13880
rect 11388 13756 11464 13828
rect 11388 13704 11400 13756
rect 11452 13704 11464 13756
rect 11388 13632 11464 13704
rect 11388 13580 11400 13632
rect 11452 13580 11464 13632
rect 11388 13508 11464 13580
rect 11388 13456 11400 13508
rect 11452 13456 11464 13508
rect 11388 13384 11464 13456
rect 11388 13332 11400 13384
rect 11452 13332 11464 13384
rect 11388 13260 11464 13332
rect 11388 13208 11400 13260
rect 11452 13208 11464 13260
rect 11388 13136 11464 13208
rect 11388 13084 11400 13136
rect 11452 13084 11464 13136
rect 11388 13012 11464 13084
rect 11388 12960 11400 13012
rect 11452 12960 11464 13012
rect 11388 12888 11464 12960
rect 11388 12836 11400 12888
rect 11452 12836 11464 12888
rect 11388 12592 11464 12836
rect 11836 14996 11912 15008
rect 11836 14944 11848 14996
rect 11900 14944 11912 14996
rect 11836 14872 11912 14944
rect 11836 14820 11848 14872
rect 11900 14820 11912 14872
rect 11836 14748 11912 14820
rect 11836 14696 11848 14748
rect 11900 14696 11912 14748
rect 11836 14624 11912 14696
rect 11836 14572 11848 14624
rect 11900 14572 11912 14624
rect 11836 14500 11912 14572
rect 11836 14448 11848 14500
rect 11900 14448 11912 14500
rect 11836 14376 11912 14448
rect 11836 14324 11848 14376
rect 11900 14324 11912 14376
rect 11836 14252 11912 14324
rect 11836 14200 11848 14252
rect 11900 14200 11912 14252
rect 11836 14128 11912 14200
rect 11836 14076 11848 14128
rect 11900 14076 11912 14128
rect 11836 14004 11912 14076
rect 11836 13952 11848 14004
rect 11900 13952 11912 14004
rect 11836 13880 11912 13952
rect 11836 13828 11848 13880
rect 11900 13828 11912 13880
rect 11836 13756 11912 13828
rect 11836 13704 11848 13756
rect 11900 13704 11912 13756
rect 11836 13632 11912 13704
rect 11836 13580 11848 13632
rect 11900 13580 11912 13632
rect 11836 13508 11912 13580
rect 11836 13456 11848 13508
rect 11900 13456 11912 13508
rect 11836 13384 11912 13456
rect 11836 13332 11848 13384
rect 11900 13332 11912 13384
rect 11836 13260 11912 13332
rect 11836 13208 11848 13260
rect 11900 13208 11912 13260
rect 11836 13136 11912 13208
rect 11836 13084 11848 13136
rect 11900 13084 11912 13136
rect 11836 13012 11912 13084
rect 11836 12960 11848 13012
rect 11900 12960 11912 13012
rect 11836 12888 11912 12960
rect 12508 14996 12584 15008
rect 12508 14944 12520 14996
rect 12572 14944 12584 14996
rect 12508 14872 12584 14944
rect 12508 14820 12520 14872
rect 12572 14820 12584 14872
rect 12508 14748 12584 14820
rect 12508 14696 12520 14748
rect 12572 14696 12584 14748
rect 12508 14624 12584 14696
rect 12508 14572 12520 14624
rect 12572 14572 12584 14624
rect 12508 14500 12584 14572
rect 12508 14448 12520 14500
rect 12572 14448 12584 14500
rect 12508 14376 12584 14448
rect 12508 14324 12520 14376
rect 12572 14324 12584 14376
rect 12508 14252 12584 14324
rect 12508 14200 12520 14252
rect 12572 14200 12584 14252
rect 12508 14128 12584 14200
rect 12508 14076 12520 14128
rect 12572 14076 12584 14128
rect 12508 14004 12584 14076
rect 12508 13952 12520 14004
rect 12572 13952 12584 14004
rect 12508 13880 12584 13952
rect 12508 13828 12520 13880
rect 12572 13828 12584 13880
rect 12508 13756 12584 13828
rect 12508 13704 12520 13756
rect 12572 13704 12584 13756
rect 12508 13632 12584 13704
rect 12508 13580 12520 13632
rect 12572 13580 12584 13632
rect 12508 13508 12584 13580
rect 12508 13456 12520 13508
rect 12572 13456 12584 13508
rect 12508 13384 12584 13456
rect 12508 13332 12520 13384
rect 12572 13332 12584 13384
rect 12508 13260 12584 13332
rect 12508 13208 12520 13260
rect 12572 13208 12584 13260
rect 12508 13136 12584 13208
rect 12508 13084 12520 13136
rect 12572 13084 12584 13136
rect 12508 13012 12584 13084
rect 12508 12960 12520 13012
rect 12572 12960 12584 13012
rect 12508 12932 12584 12960
rect 12956 14996 13032 15008
rect 12956 14944 12968 14996
rect 13020 14944 13032 14996
rect 12956 14872 13032 14944
rect 12956 14820 12968 14872
rect 13020 14820 13032 14872
rect 12956 14748 13032 14820
rect 12956 14696 12968 14748
rect 13020 14696 13032 14748
rect 12956 14624 13032 14696
rect 12956 14572 12968 14624
rect 13020 14572 13032 14624
rect 12956 14500 13032 14572
rect 12956 14448 12968 14500
rect 13020 14448 13032 14500
rect 12956 14376 13032 14448
rect 12956 14324 12968 14376
rect 13020 14324 13032 14376
rect 12956 14252 13032 14324
rect 12956 14200 12968 14252
rect 13020 14200 13032 14252
rect 12956 14128 13032 14200
rect 12956 14076 12968 14128
rect 13020 14076 13032 14128
rect 12956 14004 13032 14076
rect 12956 13952 12968 14004
rect 13020 13952 13032 14004
rect 12956 13880 13032 13952
rect 12956 13828 12968 13880
rect 13020 13828 13032 13880
rect 12956 13756 13032 13828
rect 12956 13704 12968 13756
rect 13020 13704 13032 13756
rect 12956 13632 13032 13704
rect 12956 13580 12968 13632
rect 13020 13580 13032 13632
rect 12956 13508 13032 13580
rect 12956 13456 12968 13508
rect 13020 13456 13032 13508
rect 12956 13384 13032 13456
rect 12956 13332 12968 13384
rect 13020 13332 13032 13384
rect 12956 13260 13032 13332
rect 13628 14996 13704 15008
rect 13628 14944 13640 14996
rect 13692 14944 13704 14996
rect 13628 14872 13704 14944
rect 13628 14820 13640 14872
rect 13692 14820 13704 14872
rect 13628 14748 13704 14820
rect 13628 14696 13640 14748
rect 13692 14696 13704 14748
rect 13628 14624 13704 14696
rect 13628 14572 13640 14624
rect 13692 14572 13704 14624
rect 13628 14500 13704 14572
rect 13628 14448 13640 14500
rect 13692 14448 13704 14500
rect 13628 14376 13704 14448
rect 13628 14324 13640 14376
rect 13692 14324 13704 14376
rect 13628 14252 13704 14324
rect 13628 14200 13640 14252
rect 13692 14200 13704 14252
rect 13628 14128 13704 14200
rect 13628 14076 13640 14128
rect 13692 14076 13704 14128
rect 13628 14004 13704 14076
rect 13628 13952 13640 14004
rect 13692 13952 13704 14004
rect 13628 13880 13704 13952
rect 13628 13828 13640 13880
rect 13692 13828 13704 13880
rect 13628 13756 13704 13828
rect 13628 13704 13640 13756
rect 13692 13704 13704 13756
rect 13628 13632 13704 13704
rect 13628 13580 13640 13632
rect 13692 13580 13704 13632
rect 13628 13508 13704 13580
rect 13628 13456 13640 13508
rect 13692 13456 13704 13508
rect 13628 13384 13704 13456
rect 13628 13332 13640 13384
rect 13692 13332 13704 13384
rect 13628 13272 13704 13332
rect 14076 14996 14152 15008
rect 14076 14944 14088 14996
rect 14140 14944 14152 14996
rect 14076 14872 14152 14944
rect 14076 14820 14088 14872
rect 14140 14820 14152 14872
rect 14076 14748 14152 14820
rect 14076 14696 14088 14748
rect 14140 14696 14152 14748
rect 14076 14624 14152 14696
rect 14076 14572 14088 14624
rect 14140 14572 14152 14624
rect 14076 14500 14152 14572
rect 14076 14448 14088 14500
rect 14140 14448 14152 14500
rect 14076 14376 14152 14448
rect 14076 14324 14088 14376
rect 14140 14324 14152 14376
rect 14076 14252 14152 14324
rect 14076 14200 14088 14252
rect 14140 14200 14152 14252
rect 14076 14128 14152 14200
rect 14076 14076 14088 14128
rect 14140 14076 14152 14128
rect 14076 14004 14152 14076
rect 14076 13952 14088 14004
rect 14140 13952 14152 14004
rect 14076 13880 14152 13952
rect 14076 13828 14088 13880
rect 14140 13828 14152 13880
rect 14076 13756 14152 13828
rect 14076 13704 14088 13756
rect 14140 13704 14152 13756
rect 14076 13632 14152 13704
rect 14076 13580 14088 13632
rect 14140 13580 14152 13632
rect 14748 14996 14824 15008
rect 14748 14944 14760 14996
rect 14812 14944 14824 14996
rect 14748 14872 14824 14944
rect 14748 14820 14760 14872
rect 14812 14820 14824 14872
rect 14748 14748 14824 14820
rect 14748 14696 14760 14748
rect 14812 14696 14824 14748
rect 14748 14624 14824 14696
rect 14748 14572 14760 14624
rect 14812 14572 14824 14624
rect 14748 14500 14824 14572
rect 14748 14448 14760 14500
rect 14812 14448 14824 14500
rect 14748 14376 14824 14448
rect 14748 14324 14760 14376
rect 14812 14324 14824 14376
rect 14748 14252 14824 14324
rect 14748 14200 14760 14252
rect 14812 14200 14824 14252
rect 14748 14128 14824 14200
rect 14748 14076 14760 14128
rect 14812 14076 14824 14128
rect 14748 14004 14824 14076
rect 14748 13952 14760 14004
rect 14812 13952 14824 14004
rect 14748 13880 14824 13952
rect 14748 13828 14760 13880
rect 14812 13828 14824 13880
rect 14748 13756 14824 13828
rect 14748 13704 14760 13756
rect 14812 13704 14824 13756
rect 14748 13632 14824 13704
rect 14748 13612 14760 13632
rect 14076 13508 14152 13580
rect 14076 13456 14088 13508
rect 14140 13456 14152 13508
rect 14721 13580 14760 13612
rect 14812 13612 14824 13632
rect 15196 14996 15272 15008
rect 15196 14944 15208 14996
rect 15260 14944 15272 14996
rect 15196 14872 15272 14944
rect 15196 14820 15208 14872
rect 15260 14820 15272 14872
rect 15196 14748 15272 14820
rect 15196 14696 15208 14748
rect 15260 14696 15272 14748
rect 15196 14624 15272 14696
rect 15196 14572 15208 14624
rect 15260 14572 15272 14624
rect 15196 14500 15272 14572
rect 15196 14448 15208 14500
rect 15260 14448 15272 14500
rect 15196 14376 15272 14448
rect 15196 14324 15208 14376
rect 15260 14324 15272 14376
rect 15196 14252 15272 14324
rect 15196 14200 15208 14252
rect 15260 14200 15272 14252
rect 15196 14128 15272 14200
rect 15196 14076 15208 14128
rect 15260 14076 15272 14128
rect 15196 14004 15272 14076
rect 15196 13952 15208 14004
rect 15260 13952 15272 14004
rect 15868 14996 15944 15008
rect 15868 14944 15880 14996
rect 15932 14944 15944 14996
rect 15868 14872 15944 14944
rect 15868 14820 15880 14872
rect 15932 14820 15944 14872
rect 15868 14748 15944 14820
rect 15868 14696 15880 14748
rect 15932 14696 15944 14748
rect 15868 14624 15944 14696
rect 15868 14572 15880 14624
rect 15932 14572 15944 14624
rect 15868 14500 15944 14572
rect 15868 14448 15880 14500
rect 15932 14448 15944 14500
rect 15868 14376 15944 14448
rect 15868 14324 15880 14376
rect 15932 14324 15944 14376
rect 15868 14252 15944 14324
rect 15868 14200 15880 14252
rect 15932 14200 15944 14252
rect 15868 14128 15944 14200
rect 15868 14076 15880 14128
rect 15932 14076 15944 14128
rect 15868 14004 15944 14076
rect 15868 13952 15880 14004
rect 15932 13952 15944 14004
rect 16316 14996 16392 15008
rect 16316 14944 16328 14996
rect 16380 14944 16392 14996
rect 16316 14872 16392 14944
rect 16316 14820 16328 14872
rect 16380 14820 16392 14872
rect 16316 14748 16392 14820
rect 16316 14696 16328 14748
rect 16380 14696 16392 14748
rect 16316 14624 16392 14696
rect 16316 14572 16328 14624
rect 16380 14572 16392 14624
rect 16316 14500 16392 14572
rect 16316 14448 16328 14500
rect 16380 14448 16392 14500
rect 16316 14376 16392 14448
rect 16316 14324 16328 14376
rect 16380 14324 16392 14376
rect 16316 14252 16392 14324
rect 16988 14996 17064 15008
rect 16988 14944 17000 14996
rect 17052 14944 17064 14996
rect 16988 14872 17064 14944
rect 16988 14820 17000 14872
rect 17052 14820 17064 14872
rect 16988 14748 17064 14820
rect 16988 14696 17000 14748
rect 17052 14696 17064 14748
rect 16988 14624 17064 14696
rect 16988 14572 17000 14624
rect 17052 14572 17064 14624
rect 16988 14500 17064 14572
rect 16988 14448 17000 14500
rect 17052 14448 17064 14500
rect 16988 14376 17064 14448
rect 16988 14324 17000 14376
rect 17052 14324 17064 14376
rect 16988 14292 17064 14324
rect 17436 14996 17512 15008
rect 17436 14944 17448 14996
rect 17500 14944 17512 14996
rect 17436 14872 17512 14944
rect 17436 14820 17448 14872
rect 17500 14820 17512 14872
rect 17436 14748 17512 14820
rect 17436 14696 17448 14748
rect 17500 14696 17512 14748
rect 17436 14624 17512 14696
rect 18108 14996 18184 15008
rect 18108 14944 18120 14996
rect 18172 14944 18184 14996
rect 18108 14872 18184 14944
rect 18108 14820 18120 14872
rect 18172 14820 18184 14872
rect 18108 14748 18184 14820
rect 18108 14696 18120 14748
rect 18172 14696 18184 14748
rect 18108 14633 18184 14696
rect 18556 14996 18632 15008
rect 18556 14944 18568 14996
rect 18620 14944 18632 14996
rect 19228 14996 19304 15008
rect 19228 14973 19240 14996
rect 18556 14872 18632 14944
rect 18556 14820 18568 14872
rect 18620 14820 18632 14872
rect 19201 14944 19240 14973
rect 19292 14973 19304 14996
rect 19676 14996 19752 15008
rect 19676 14973 19688 14996
rect 19292 14944 19330 14973
rect 19201 14934 19330 14944
rect 19201 14878 19237 14934
rect 19293 14878 19330 14934
rect 19201 14872 19330 14878
rect 19201 14839 19240 14872
rect 18556 14748 18632 14820
rect 18556 14696 18568 14748
rect 18620 14696 18632 14748
rect 18556 14633 18632 14696
rect 19228 14820 19240 14839
rect 19292 14839 19330 14872
rect 19649 14944 19688 14973
rect 19740 14973 19752 14996
rect 19740 14944 19778 14973
rect 19649 14934 19778 14944
rect 19649 14878 19685 14934
rect 19741 14878 19778 14934
rect 19649 14872 19778 14878
rect 19649 14839 19688 14872
rect 19292 14820 19304 14839
rect 19228 14748 19304 14820
rect 19228 14696 19240 14748
rect 19292 14696 19304 14748
rect 17436 14572 17448 14624
rect 17500 14572 17512 14624
rect 17436 14500 17512 14572
rect 17436 14448 17448 14500
rect 17500 14448 17512 14500
rect 18081 14624 18210 14633
rect 18081 14594 18120 14624
rect 18172 14594 18210 14624
rect 18081 14538 18117 14594
rect 18173 14538 18210 14594
rect 18081 14500 18210 14538
rect 18081 14499 18120 14500
rect 17436 14376 17512 14448
rect 17436 14324 17448 14376
rect 17500 14324 17512 14376
rect 17436 14292 17512 14324
rect 18108 14448 18120 14499
rect 18172 14499 18210 14500
rect 18529 14624 18658 14633
rect 18529 14594 18568 14624
rect 18620 14594 18658 14624
rect 18529 14538 18565 14594
rect 18621 14538 18658 14594
rect 18529 14500 18658 14538
rect 18529 14499 18568 14500
rect 18172 14448 18184 14499
rect 18108 14376 18184 14448
rect 18108 14324 18120 14376
rect 18172 14324 18184 14376
rect 16316 14200 16328 14252
rect 16380 14200 16392 14252
rect 16316 14128 16392 14200
rect 16961 14253 17090 14292
rect 16961 14197 16997 14253
rect 17053 14197 17090 14253
rect 16961 14158 17090 14197
rect 17409 14253 17538 14292
rect 17409 14197 17445 14253
rect 17501 14197 17538 14253
rect 17409 14158 17538 14197
rect 18108 14252 18184 14324
rect 18108 14200 18120 14252
rect 18172 14200 18184 14252
rect 16316 14076 16328 14128
rect 16380 14076 16392 14128
rect 16316 14004 16392 14076
rect 16316 13952 16328 14004
rect 16380 13952 16392 14004
rect 16988 14128 17064 14158
rect 16988 14076 17000 14128
rect 17052 14076 17064 14128
rect 16988 14004 17064 14076
rect 16988 13952 17000 14004
rect 17052 13952 17064 14004
rect 15196 13880 15272 13952
rect 15196 13828 15208 13880
rect 15260 13828 15272 13880
rect 15196 13756 15272 13828
rect 15841 13913 15970 13952
rect 15841 13857 15877 13913
rect 15933 13857 15970 13913
rect 15841 13828 15880 13857
rect 15932 13828 15970 13857
rect 15841 13818 15970 13828
rect 16289 13913 16418 13952
rect 16289 13857 16325 13913
rect 16381 13857 16418 13913
rect 16289 13828 16328 13857
rect 16380 13828 16418 13857
rect 16289 13818 16418 13828
rect 16988 13880 17064 13952
rect 16988 13828 17000 13880
rect 17052 13828 17064 13880
rect 15196 13704 15208 13756
rect 15260 13704 15272 13756
rect 15196 13632 15272 13704
rect 15196 13612 15208 13632
rect 14812 13580 14850 13612
rect 14721 13573 14850 13580
rect 14721 13517 14757 13573
rect 14813 13517 14850 13573
rect 14721 13508 14850 13517
rect 14721 13478 14760 13508
rect 14076 13384 14152 13456
rect 14076 13332 14088 13384
rect 14140 13332 14152 13384
rect 14076 13272 14152 13332
rect 14748 13456 14760 13478
rect 14812 13478 14850 13508
rect 15169 13580 15208 13612
rect 15260 13612 15272 13632
rect 15868 13756 15944 13818
rect 15868 13704 15880 13756
rect 15932 13704 15944 13756
rect 15868 13632 15944 13704
rect 15260 13580 15298 13612
rect 15169 13573 15298 13580
rect 15169 13517 15205 13573
rect 15261 13517 15298 13573
rect 15169 13508 15298 13517
rect 15169 13478 15208 13508
rect 14812 13456 14824 13478
rect 14748 13384 14824 13456
rect 14748 13332 14760 13384
rect 14812 13332 14824 13384
rect 12956 13208 12968 13260
rect 13020 13208 13032 13260
rect 12956 13136 13032 13208
rect 13601 13260 13730 13272
rect 13601 13233 13640 13260
rect 13692 13233 13730 13260
rect 13601 13177 13637 13233
rect 13693 13177 13730 13233
rect 13601 13138 13730 13177
rect 14049 13260 14178 13272
rect 14049 13233 14088 13260
rect 14140 13233 14178 13260
rect 14049 13177 14085 13233
rect 14141 13177 14178 13233
rect 14049 13138 14178 13177
rect 14748 13260 14824 13332
rect 14748 13208 14760 13260
rect 14812 13208 14824 13260
rect 12956 13084 12968 13136
rect 13020 13084 13032 13136
rect 12956 13012 13032 13084
rect 12956 12960 12968 13012
rect 13020 12960 13032 13012
rect 12956 12932 13032 12960
rect 13628 13136 13704 13138
rect 13628 13084 13640 13136
rect 13692 13084 13704 13136
rect 13628 13012 13704 13084
rect 13628 12960 13640 13012
rect 13692 12960 13704 13012
rect 11836 12836 11848 12888
rect 11900 12836 11912 12888
rect 11836 12592 11912 12836
rect 12481 12893 12610 12932
rect 12481 12837 12517 12893
rect 12573 12837 12610 12893
rect 12481 12836 12520 12837
rect 12572 12836 12610 12837
rect 12481 12798 12610 12836
rect 12929 12893 13058 12932
rect 12929 12837 12965 12893
rect 13021 12837 13058 12893
rect 12929 12836 12968 12837
rect 13020 12836 13058 12837
rect 12929 12798 13058 12836
rect 13628 12888 13704 12960
rect 13628 12836 13640 12888
rect 13692 12836 13704 12888
rect 11361 12553 11490 12592
rect 11361 12497 11397 12553
rect 11453 12497 11490 12553
rect 11361 12458 11490 12497
rect 11809 12553 11938 12592
rect 11809 12497 11845 12553
rect 11901 12497 11938 12553
rect 11809 12458 11938 12497
rect 10928 12059 11268 12098
rect 10928 12003 10964 12059
rect 11020 12003 11176 12059
rect 11232 12003 11268 12059
rect 10928 11964 11268 12003
rect 10956 11911 11032 11964
rect 10956 11859 10968 11911
rect 11020 11859 11032 11911
rect 10956 11847 11032 11859
rect 10716 11706 10728 11758
rect 10780 11706 10792 11758
rect 10716 11634 10792 11706
rect 10716 11582 10728 11634
rect 10780 11582 10792 11634
rect 10716 11510 10792 11582
rect 10716 11458 10728 11510
rect 10780 11458 10792 11510
rect 11388 11758 11464 12458
rect 11388 11706 11400 11758
rect 11452 11706 11464 11758
rect 11388 11634 11464 11706
rect 11836 11758 11912 12458
rect 12076 11911 12152 12009
rect 12076 11889 12088 11911
rect 11836 11706 11848 11758
rect 11900 11706 11912 11758
rect 11388 11582 11400 11634
rect 11452 11582 11464 11634
rect 11388 11510 11464 11582
rect 11582 11660 11711 11681
rect 11582 11642 11712 11660
rect 11582 11586 11619 11642
rect 11675 11586 11712 11642
rect 11582 11547 11712 11586
rect 10716 11446 10792 11458
rect 10915 11433 11255 11472
rect 11388 11458 11400 11510
rect 11452 11458 11464 11510
rect 11388 11446 11464 11458
rect 10915 11377 10951 11433
rect 11007 11377 11163 11433
rect 11219 11377 11255 11433
rect 10915 11338 11255 11377
rect 10232 11225 10572 11264
rect 10232 11169 10268 11225
rect 10324 11169 10480 11225
rect 10536 11169 10572 11225
rect 10232 11130 10572 11169
rect 9808 10599 10148 10638
rect 9808 10543 9844 10599
rect 9900 10543 10056 10599
rect 10112 10543 10148 10599
rect 9808 10504 10148 10543
rect 10338 10200 10467 11130
rect 9936 10067 10467 10200
rect 9714 9326 9842 9363
rect 9492 8973 9620 9287
rect 9492 8921 9530 8973
rect 9582 8921 9620 8973
rect 9492 8755 9620 8921
rect 9492 8703 9530 8755
rect 9582 8703 9620 8755
rect 8303 8485 8341 8537
rect 8393 8485 8431 8537
rect 8303 8445 8431 8485
rect 9492 8537 9620 8703
rect 9714 9270 9750 9326
rect 9806 9270 9842 9326
rect 9714 9108 9842 9270
rect 9714 9052 9750 9108
rect 9806 9052 9842 9108
rect 9714 8890 9842 9052
rect 9714 8834 9750 8890
rect 9806 8834 9842 8890
rect 9714 8672 9842 8834
rect 9714 8616 9750 8672
rect 9806 8616 9842 8672
rect 9714 8578 9842 8616
rect 9936 9287 10065 10067
rect 10162 9326 10290 9363
rect 9936 8973 10064 9287
rect 9936 8921 9974 8973
rect 10026 8921 10064 8973
rect 9936 8755 10064 8921
rect 9936 8703 9974 8755
rect 10026 8703 10064 8755
rect 9492 8485 9530 8537
rect 9582 8485 9620 8537
rect 9492 8445 9620 8485
rect 9936 8537 10064 8703
rect 10162 9270 10198 9326
rect 10254 9270 10290 9326
rect 10162 9108 10290 9270
rect 10162 9052 10198 9108
rect 10254 9052 10290 9108
rect 10162 8890 10290 9052
rect 10162 8834 10198 8890
rect 10254 8834 10290 8890
rect 10162 8672 10290 8834
rect 10162 8616 10198 8672
rect 10254 8616 10290 8672
rect 10162 8578 10290 8616
rect 10900 9326 11028 9363
rect 10900 9270 10936 9326
rect 10992 9270 11028 9326
rect 10900 9108 11028 9270
rect 10900 9052 10936 9108
rect 10992 9052 11028 9108
rect 10900 8890 11028 9052
rect 10900 8834 10936 8890
rect 10992 8834 11028 8890
rect 10900 8672 11028 8834
rect 10900 8616 10936 8672
rect 10992 8616 11028 8672
rect 10900 8578 11028 8616
rect 11126 9287 11255 11338
rect 11583 10076 11712 11547
rect 11836 11634 11912 11706
rect 11836 11582 11848 11634
rect 11900 11582 11912 11634
rect 11836 11510 11912 11582
rect 11836 11458 11848 11510
rect 11900 11458 11912 11510
rect 11836 11446 11912 11458
rect 12048 11859 12088 11889
rect 12140 11889 12152 11911
rect 12140 11859 12388 11889
rect 12048 11850 12388 11859
rect 12048 11794 12084 11850
rect 12140 11794 12296 11850
rect 12352 11794 12388 11850
rect 12048 11755 12388 11794
rect 12508 11758 12584 12798
rect 12706 12168 12831 12207
rect 12706 12112 12741 12168
rect 12797 12112 12831 12168
rect 12706 12098 12831 12112
rect 11570 9942 11712 10076
rect 12048 10101 12177 11755
rect 12508 11706 12520 11758
rect 12572 11706 12584 11758
rect 12508 11634 12584 11706
rect 12508 11582 12520 11634
rect 12572 11582 12584 11634
rect 12508 11510 12584 11582
rect 12508 11458 12520 11510
rect 12572 11458 12584 11510
rect 12508 11446 12584 11458
rect 12705 11950 12834 12098
rect 12705 11894 12741 11950
rect 12797 11894 12834 11950
rect 12705 10465 12834 11894
rect 12956 11758 13032 12798
rect 13196 11973 13272 12009
rect 12956 11706 12968 11758
rect 13020 11706 13032 11758
rect 12956 11634 13032 11706
rect 12956 11582 12968 11634
rect 13020 11582 13032 11634
rect 12956 11510 13032 11582
rect 13168 11911 13297 11973
rect 13168 11859 13208 11911
rect 13260 11859 13297 11911
rect 13168 11688 13297 11859
rect 13628 11758 13704 12836
rect 13628 11706 13640 11758
rect 13692 11706 13704 11758
rect 13168 11687 13298 11688
rect 13168 11649 13507 11687
rect 13168 11593 13204 11649
rect 13260 11593 13416 11649
rect 13472 11593 13507 11649
rect 13168 11554 13507 11593
rect 13628 11634 13704 11706
rect 13628 11582 13640 11634
rect 13692 11582 13704 11634
rect 12956 11458 12968 11510
rect 13020 11458 13032 11510
rect 12956 11446 13032 11458
rect 13628 11510 13704 11582
rect 13628 11458 13640 11510
rect 13692 11458 13704 11510
rect 13628 11446 13704 11458
rect 14076 13136 14152 13138
rect 14076 13084 14088 13136
rect 14140 13084 14152 13136
rect 14076 13012 14152 13084
rect 14076 12960 14088 13012
rect 14140 12960 14152 13012
rect 14076 12888 14152 12960
rect 14076 12836 14088 12888
rect 14140 12836 14152 12888
rect 14076 11758 14152 12836
rect 14748 13136 14824 13208
rect 14748 13084 14760 13136
rect 14812 13084 14824 13136
rect 14748 13012 14824 13084
rect 14748 12960 14760 13012
rect 14812 12960 14824 13012
rect 14748 12888 14824 12960
rect 14748 12836 14760 12888
rect 14812 12836 14824 12888
rect 14316 11973 14392 12009
rect 14076 11706 14088 11758
rect 14140 11706 14152 11758
rect 14076 11634 14152 11706
rect 14076 11582 14088 11634
rect 14140 11582 14152 11634
rect 14076 11510 14152 11582
rect 14076 11458 14088 11510
rect 14140 11458 14152 11510
rect 14076 11446 14152 11458
rect 14288 11911 14417 11973
rect 14288 11859 14328 11911
rect 14380 11859 14417 11911
rect 14288 11672 14417 11859
rect 14288 11616 14325 11672
rect 14381 11616 14417 11672
rect 14288 11454 14417 11616
rect 14288 11398 14325 11454
rect 14381 11398 14417 11454
rect 14748 11758 14824 12836
rect 14748 11706 14760 11758
rect 14812 11706 14824 11758
rect 14748 11634 14824 11706
rect 14748 11582 14760 11634
rect 14812 11582 14824 11634
rect 14748 11510 14824 11582
rect 14748 11458 14760 11510
rect 14812 11458 14824 11510
rect 14748 11446 14824 11458
rect 15196 13456 15208 13478
rect 15260 13478 15298 13508
rect 15868 13580 15880 13632
rect 15932 13580 15944 13632
rect 15868 13508 15944 13580
rect 15260 13456 15272 13478
rect 15196 13384 15272 13456
rect 15196 13332 15208 13384
rect 15260 13332 15272 13384
rect 15196 13260 15272 13332
rect 15196 13208 15208 13260
rect 15260 13208 15272 13260
rect 15196 13136 15272 13208
rect 15196 13084 15208 13136
rect 15260 13084 15272 13136
rect 15196 13012 15272 13084
rect 15196 12960 15208 13012
rect 15260 12960 15272 13012
rect 15196 12888 15272 12960
rect 15196 12836 15208 12888
rect 15260 12836 15272 12888
rect 15196 11758 15272 12836
rect 15868 13456 15880 13508
rect 15932 13456 15944 13508
rect 15868 13384 15944 13456
rect 15868 13332 15880 13384
rect 15932 13332 15944 13384
rect 15868 13260 15944 13332
rect 15868 13208 15880 13260
rect 15932 13208 15944 13260
rect 15868 13136 15944 13208
rect 15868 13084 15880 13136
rect 15932 13084 15944 13136
rect 15868 13012 15944 13084
rect 15868 12960 15880 13012
rect 15932 12960 15944 13012
rect 15868 12888 15944 12960
rect 15868 12836 15880 12888
rect 15932 12836 15944 12888
rect 15436 11973 15512 12009
rect 15196 11706 15208 11758
rect 15260 11706 15272 11758
rect 15196 11634 15272 11706
rect 15196 11582 15208 11634
rect 15260 11582 15272 11634
rect 15196 11510 15272 11582
rect 15196 11458 15208 11510
rect 15260 11458 15272 11510
rect 15196 11446 15272 11458
rect 15408 11911 15537 11973
rect 15408 11859 15448 11911
rect 15500 11859 15537 11911
rect 15408 11463 15537 11859
rect 14288 11359 14417 11398
rect 15408 11407 15445 11463
rect 15501 11407 15537 11463
rect 15868 11758 15944 12836
rect 15868 11706 15880 11758
rect 15932 11706 15944 11758
rect 15868 11634 15944 11706
rect 15868 11582 15880 11634
rect 15932 11582 15944 11634
rect 15868 11510 15944 11582
rect 15868 11458 15880 11510
rect 15932 11458 15944 11510
rect 15868 11446 15944 11458
rect 16316 13756 16392 13818
rect 16316 13704 16328 13756
rect 16380 13704 16392 13756
rect 16316 13632 16392 13704
rect 16316 13580 16328 13632
rect 16380 13580 16392 13632
rect 16316 13508 16392 13580
rect 16316 13456 16328 13508
rect 16380 13456 16392 13508
rect 16316 13384 16392 13456
rect 16316 13332 16328 13384
rect 16380 13332 16392 13384
rect 16316 13260 16392 13332
rect 16316 13208 16328 13260
rect 16380 13208 16392 13260
rect 16316 13136 16392 13208
rect 16316 13084 16328 13136
rect 16380 13084 16392 13136
rect 16316 13012 16392 13084
rect 16316 12960 16328 13012
rect 16380 12960 16392 13012
rect 16316 12888 16392 12960
rect 16316 12836 16328 12888
rect 16380 12836 16392 12888
rect 16316 11758 16392 12836
rect 16988 13756 17064 13828
rect 16988 13704 17000 13756
rect 17052 13704 17064 13756
rect 16988 13632 17064 13704
rect 16988 13580 17000 13632
rect 17052 13580 17064 13632
rect 16988 13508 17064 13580
rect 16988 13456 17000 13508
rect 17052 13456 17064 13508
rect 16988 13384 17064 13456
rect 16988 13332 17000 13384
rect 17052 13332 17064 13384
rect 16988 13260 17064 13332
rect 16988 13208 17000 13260
rect 17052 13208 17064 13260
rect 16988 13136 17064 13208
rect 16988 13084 17000 13136
rect 17052 13084 17064 13136
rect 16988 13012 17064 13084
rect 16988 12960 17000 13012
rect 17052 12960 17064 13012
rect 16988 12888 17064 12960
rect 16988 12836 17000 12888
rect 17052 12836 17064 12888
rect 16556 11973 16632 12009
rect 16316 11706 16328 11758
rect 16380 11706 16392 11758
rect 16316 11634 16392 11706
rect 16316 11582 16328 11634
rect 16380 11582 16392 11634
rect 16316 11510 16392 11582
rect 16316 11458 16328 11510
rect 16380 11458 16392 11510
rect 16316 11446 16392 11458
rect 16528 11911 16657 11973
rect 16528 11859 16568 11911
rect 16620 11859 16657 11911
rect 15408 11245 15537 11407
rect 15408 11189 15445 11245
rect 15501 11189 15537 11245
rect 15408 11150 15537 11189
rect 16528 11254 16657 11859
rect 16988 11758 17064 12836
rect 16988 11706 17000 11758
rect 17052 11706 17064 11758
rect 16988 11634 17064 11706
rect 16988 11582 17000 11634
rect 17052 11582 17064 11634
rect 16988 11510 17064 11582
rect 16988 11458 17000 11510
rect 17052 11458 17064 11510
rect 16988 11446 17064 11458
rect 17436 14128 17512 14158
rect 17436 14076 17448 14128
rect 17500 14076 17512 14128
rect 17436 14004 17512 14076
rect 17436 13952 17448 14004
rect 17500 13952 17512 14004
rect 17436 13880 17512 13952
rect 17436 13828 17448 13880
rect 17500 13828 17512 13880
rect 17436 13756 17512 13828
rect 17436 13704 17448 13756
rect 17500 13704 17512 13756
rect 17436 13632 17512 13704
rect 17436 13580 17448 13632
rect 17500 13580 17512 13632
rect 17436 13508 17512 13580
rect 17436 13456 17448 13508
rect 17500 13456 17512 13508
rect 17436 13384 17512 13456
rect 17436 13332 17448 13384
rect 17500 13332 17512 13384
rect 17436 13260 17512 13332
rect 17436 13208 17448 13260
rect 17500 13208 17512 13260
rect 17436 13136 17512 13208
rect 17436 13084 17448 13136
rect 17500 13084 17512 13136
rect 17436 13012 17512 13084
rect 17436 12960 17448 13012
rect 17500 12960 17512 13012
rect 17436 12888 17512 12960
rect 17436 12836 17448 12888
rect 17500 12836 17512 12888
rect 17436 11758 17512 12836
rect 18108 14128 18184 14200
rect 18108 14076 18120 14128
rect 18172 14076 18184 14128
rect 18108 14004 18184 14076
rect 18108 13952 18120 14004
rect 18172 13952 18184 14004
rect 18108 13880 18184 13952
rect 18108 13828 18120 13880
rect 18172 13828 18184 13880
rect 18108 13756 18184 13828
rect 18108 13704 18120 13756
rect 18172 13704 18184 13756
rect 18108 13632 18184 13704
rect 18108 13580 18120 13632
rect 18172 13580 18184 13632
rect 18108 13508 18184 13580
rect 18108 13456 18120 13508
rect 18172 13456 18184 13508
rect 18108 13384 18184 13456
rect 18108 13332 18120 13384
rect 18172 13332 18184 13384
rect 18108 13260 18184 13332
rect 18108 13208 18120 13260
rect 18172 13208 18184 13260
rect 18108 13136 18184 13208
rect 18108 13084 18120 13136
rect 18172 13084 18184 13136
rect 18108 13012 18184 13084
rect 18108 12960 18120 13012
rect 18172 12960 18184 13012
rect 18108 12888 18184 12960
rect 18108 12836 18120 12888
rect 18172 12836 18184 12888
rect 17676 11973 17752 12009
rect 17436 11706 17448 11758
rect 17500 11706 17512 11758
rect 17436 11634 17512 11706
rect 17436 11582 17448 11634
rect 17500 11582 17512 11634
rect 17436 11510 17512 11582
rect 17436 11458 17448 11510
rect 17500 11458 17512 11510
rect 17436 11446 17512 11458
rect 17648 11911 17777 11973
rect 17648 11859 17688 11911
rect 17740 11859 17777 11911
rect 16528 11198 16565 11254
rect 16621 11198 16657 11254
rect 16528 11036 16657 11198
rect 16528 10980 16565 11036
rect 16621 10980 16657 11036
rect 16528 10942 16657 10980
rect 17648 11046 17777 11859
rect 18108 11758 18184 12836
rect 18108 11706 18120 11758
rect 18172 11706 18184 11758
rect 18108 11634 18184 11706
rect 18108 11582 18120 11634
rect 18172 11582 18184 11634
rect 18108 11510 18184 11582
rect 18108 11458 18120 11510
rect 18172 11458 18184 11510
rect 18108 11446 18184 11458
rect 18556 14448 18568 14499
rect 18620 14499 18658 14500
rect 19228 14624 19304 14696
rect 19228 14572 19240 14624
rect 19292 14572 19304 14624
rect 19228 14500 19304 14572
rect 18620 14448 18632 14499
rect 18556 14376 18632 14448
rect 18556 14324 18568 14376
rect 18620 14324 18632 14376
rect 18556 14252 18632 14324
rect 18556 14200 18568 14252
rect 18620 14200 18632 14252
rect 18556 14128 18632 14200
rect 18556 14076 18568 14128
rect 18620 14076 18632 14128
rect 18556 14004 18632 14076
rect 18556 13952 18568 14004
rect 18620 13952 18632 14004
rect 18556 13880 18632 13952
rect 18556 13828 18568 13880
rect 18620 13828 18632 13880
rect 18556 13756 18632 13828
rect 18556 13704 18568 13756
rect 18620 13704 18632 13756
rect 18556 13632 18632 13704
rect 18556 13580 18568 13632
rect 18620 13580 18632 13632
rect 18556 13508 18632 13580
rect 18556 13456 18568 13508
rect 18620 13456 18632 13508
rect 18556 13384 18632 13456
rect 18556 13332 18568 13384
rect 18620 13332 18632 13384
rect 18556 13260 18632 13332
rect 18556 13208 18568 13260
rect 18620 13208 18632 13260
rect 18556 13136 18632 13208
rect 18556 13084 18568 13136
rect 18620 13084 18632 13136
rect 18556 13012 18632 13084
rect 18556 12960 18568 13012
rect 18620 12960 18632 13012
rect 18556 12888 18632 12960
rect 18556 12836 18568 12888
rect 18620 12836 18632 12888
rect 18556 11758 18632 12836
rect 19228 14448 19240 14500
rect 19292 14448 19304 14500
rect 19228 14376 19304 14448
rect 19228 14324 19240 14376
rect 19292 14324 19304 14376
rect 19228 14252 19304 14324
rect 19228 14200 19240 14252
rect 19292 14200 19304 14252
rect 19228 14128 19304 14200
rect 19228 14076 19240 14128
rect 19292 14076 19304 14128
rect 19228 14004 19304 14076
rect 19228 13952 19240 14004
rect 19292 13952 19304 14004
rect 19228 13880 19304 13952
rect 19228 13828 19240 13880
rect 19292 13828 19304 13880
rect 19228 13756 19304 13828
rect 19228 13704 19240 13756
rect 19292 13704 19304 13756
rect 19228 13632 19304 13704
rect 19228 13580 19240 13632
rect 19292 13580 19304 13632
rect 19228 13508 19304 13580
rect 19228 13456 19240 13508
rect 19292 13456 19304 13508
rect 19228 13384 19304 13456
rect 19228 13332 19240 13384
rect 19292 13332 19304 13384
rect 19228 13260 19304 13332
rect 19228 13208 19240 13260
rect 19292 13208 19304 13260
rect 19228 13136 19304 13208
rect 19228 13084 19240 13136
rect 19292 13084 19304 13136
rect 19228 13012 19304 13084
rect 19228 12960 19240 13012
rect 19292 12960 19304 13012
rect 19228 12888 19304 12960
rect 19228 12836 19240 12888
rect 19292 12836 19304 12888
rect 18556 11706 18568 11758
rect 18620 11706 18632 11758
rect 18556 11634 18632 11706
rect 18556 11582 18568 11634
rect 18620 11582 18632 11634
rect 18556 11510 18632 11582
rect 18556 11458 18568 11510
rect 18620 11458 18632 11510
rect 18556 11446 18632 11458
rect 18768 11911 18897 12191
rect 18768 11859 18808 11911
rect 18860 11859 18897 11911
rect 17648 10990 17685 11046
rect 17741 10990 17777 11046
rect 17648 10828 17777 10990
rect 17648 10772 17685 10828
rect 17741 10772 17777 10828
rect 17648 10733 17777 10772
rect 18768 10837 18897 11859
rect 19228 11758 19304 12836
rect 19228 11706 19240 11758
rect 19292 11706 19304 11758
rect 19228 11634 19304 11706
rect 19228 11582 19240 11634
rect 19292 11582 19304 11634
rect 19228 11510 19304 11582
rect 19228 11458 19240 11510
rect 19292 11458 19304 11510
rect 19228 11446 19304 11458
rect 19676 14820 19688 14839
rect 19740 14839 19778 14872
rect 19740 14820 19752 14839
rect 19676 14748 19752 14820
rect 19676 14696 19688 14748
rect 19740 14696 19752 14748
rect 19676 14624 19752 14696
rect 19676 14572 19688 14624
rect 19740 14572 19752 14624
rect 19676 14500 19752 14572
rect 19676 14448 19688 14500
rect 19740 14448 19752 14500
rect 19676 14376 19752 14448
rect 19676 14324 19688 14376
rect 19740 14324 19752 14376
rect 19676 14252 19752 14324
rect 19676 14200 19688 14252
rect 19740 14200 19752 14252
rect 19676 14128 19752 14200
rect 19676 14076 19688 14128
rect 19740 14076 19752 14128
rect 19676 14004 19752 14076
rect 19676 13952 19688 14004
rect 19740 13952 19752 14004
rect 19676 13880 19752 13952
rect 19676 13828 19688 13880
rect 19740 13828 19752 13880
rect 19676 13756 19752 13828
rect 19676 13704 19688 13756
rect 19740 13704 19752 13756
rect 19676 13632 19752 13704
rect 19676 13580 19688 13632
rect 19740 13580 19752 13632
rect 19676 13508 19752 13580
rect 19676 13456 19688 13508
rect 19740 13456 19752 13508
rect 19676 13384 19752 13456
rect 19676 13332 19688 13384
rect 19740 13332 19752 13384
rect 19676 13260 19752 13332
rect 19676 13208 19688 13260
rect 19740 13208 19752 13260
rect 19676 13136 19752 13208
rect 19676 13084 19688 13136
rect 19740 13084 19752 13136
rect 19676 13012 19752 13084
rect 19676 12960 19688 13012
rect 19740 12960 19752 13012
rect 19676 12888 19752 12960
rect 19676 12836 19688 12888
rect 19740 12836 19752 12888
rect 19676 11758 19752 12836
rect 19676 11706 19688 11758
rect 19740 11706 19752 11758
rect 19676 11634 19752 11706
rect 19676 11582 19688 11634
rect 19740 11582 19752 11634
rect 19676 11510 19752 11582
rect 19676 11458 19688 11510
rect 19740 11458 19752 11510
rect 19676 11446 19752 11458
rect 18768 10781 18805 10837
rect 18861 10781 18897 10837
rect 18768 10619 18897 10781
rect 18768 10563 18805 10619
rect 18861 10563 18897 10619
rect 18768 10525 18897 10563
rect 12705 10332 13333 10465
rect 12048 10100 12178 10101
rect 12048 9967 12889 10100
rect 11348 9326 11476 9363
rect 11126 8973 11254 9287
rect 11126 8921 11164 8973
rect 11216 8921 11254 8973
rect 11126 8755 11254 8921
rect 11126 8703 11164 8755
rect 11216 8703 11254 8755
rect 9936 8485 9974 8537
rect 10026 8485 10064 8537
rect 9936 8445 10064 8485
rect 11126 8537 11254 8703
rect 11348 9270 11384 9326
rect 11440 9270 11476 9326
rect 11348 9108 11476 9270
rect 11348 9052 11384 9108
rect 11440 9052 11476 9108
rect 11348 8890 11476 9052
rect 11348 8834 11384 8890
rect 11440 8834 11476 8890
rect 11348 8672 11476 8834
rect 11348 8616 11384 8672
rect 11440 8616 11476 8672
rect 11348 8578 11476 8616
rect 11570 9287 11699 9942
rect 11796 9326 11924 9363
rect 11570 8973 11698 9287
rect 11570 8921 11608 8973
rect 11660 8921 11698 8973
rect 11570 8755 11698 8921
rect 11570 8703 11608 8755
rect 11660 8703 11698 8755
rect 11126 8485 11164 8537
rect 11216 8485 11254 8537
rect 11126 8445 11254 8485
rect 11570 8537 11698 8703
rect 11796 9270 11832 9326
rect 11888 9270 11924 9326
rect 11796 9108 11924 9270
rect 11796 9052 11832 9108
rect 11888 9052 11924 9108
rect 11796 8890 11924 9052
rect 11796 8834 11832 8890
rect 11888 8834 11924 8890
rect 11796 8672 11924 8834
rect 11796 8616 11832 8672
rect 11888 8616 11924 8672
rect 11796 8578 11924 8616
rect 12534 9326 12662 9363
rect 12534 9270 12570 9326
rect 12626 9270 12662 9326
rect 12534 9108 12662 9270
rect 12534 9052 12570 9108
rect 12626 9052 12662 9108
rect 12534 8890 12662 9052
rect 12534 8834 12570 8890
rect 12626 8834 12662 8890
rect 12534 8672 12662 8834
rect 12534 8616 12570 8672
rect 12626 8616 12662 8672
rect 12534 8578 12662 8616
rect 12760 9287 12889 9967
rect 12982 9326 13110 9363
rect 12760 8973 12888 9287
rect 12760 8921 12798 8973
rect 12850 8921 12888 8973
rect 12760 8755 12888 8921
rect 12760 8703 12798 8755
rect 12850 8703 12888 8755
rect 11570 8485 11608 8537
rect 11660 8485 11698 8537
rect 11570 8445 11698 8485
rect 12760 8537 12888 8703
rect 12982 9270 13018 9326
rect 13074 9270 13110 9326
rect 12982 9108 13110 9270
rect 12982 9052 13018 9108
rect 13074 9052 13110 9108
rect 12982 8890 13110 9052
rect 12982 8834 13018 8890
rect 13074 8834 13110 8890
rect 12982 8672 13110 8834
rect 12982 8616 13018 8672
rect 13074 8616 13110 8672
rect 12982 8578 13110 8616
rect 13204 9287 13333 10332
rect 28532 10044 29412 29316
rect 29525 28998 29650 29037
rect 29525 28942 29559 28998
rect 29615 28942 29650 28998
rect 29525 28780 29650 28942
rect 29525 28724 29559 28780
rect 29615 28724 29650 28780
rect 29525 28686 29650 28724
rect 28532 9988 28627 10044
rect 28683 9988 28838 10044
rect 28894 9988 29050 10044
rect 29106 9988 29261 10044
rect 29317 9988 29412 10044
rect 28532 9826 29412 9988
rect 28532 9770 28627 9826
rect 28683 9770 28838 9826
rect 28894 9770 29050 9826
rect 29106 9770 29261 9826
rect 29317 9770 29412 9826
rect 28532 9608 29412 9770
rect 28532 9552 28627 9608
rect 28683 9552 28838 9608
rect 28894 9552 29050 9608
rect 29106 9552 29261 9608
rect 29317 9552 29412 9608
rect 28532 9390 29412 9552
rect 13430 9326 13558 9363
rect 13204 8973 13332 9287
rect 13204 8921 13242 8973
rect 13294 8921 13332 8973
rect 13204 8755 13332 8921
rect 13204 8703 13242 8755
rect 13294 8703 13332 8755
rect 12760 8485 12798 8537
rect 12850 8485 12888 8537
rect 12760 8445 12888 8485
rect 13204 8537 13332 8703
rect 13430 9270 13466 9326
rect 13522 9270 13558 9326
rect 13430 9108 13558 9270
rect 13430 9052 13466 9108
rect 13522 9052 13558 9108
rect 13430 8890 13558 9052
rect 13430 8834 13466 8890
rect 13522 8834 13558 8890
rect 13430 8672 13558 8834
rect 13430 8616 13466 8672
rect 13522 8616 13558 8672
rect 13430 8578 13558 8616
rect 28532 9334 28627 9390
rect 28683 9334 28838 9390
rect 28894 9334 29050 9390
rect 29106 9334 29261 9390
rect 29317 9334 29412 9390
rect 13204 8485 13242 8537
rect 13294 8485 13332 8537
rect 13204 8445 13332 8485
rect 2366 8142 2706 8183
rect 2366 8090 2404 8142
rect 2456 8090 2616 8142
rect 2668 8090 2706 8142
rect 2366 8050 2706 8090
rect 4057 8142 4397 8183
rect 4057 8090 4095 8142
rect 4147 8090 4307 8142
rect 4359 8090 4397 8142
rect 4057 8050 4397 8090
rect 5748 8142 6088 8183
rect 5748 8090 5786 8142
rect 5838 8090 5998 8142
rect 6050 8090 6088 8142
rect 5748 8050 6088 8090
rect 2366 3211 2495 8050
rect 2586 7881 2714 7920
rect 2586 7825 2622 7881
rect 2678 7825 2714 7881
rect 2586 7664 2714 7825
rect 2586 7608 2622 7664
rect 2678 7608 2714 7664
rect 2586 7446 2714 7608
rect 2586 7390 2622 7446
rect 2678 7390 2714 7446
rect 2586 7228 2714 7390
rect 2586 7172 2622 7228
rect 2678 7172 2714 7228
rect 2586 7010 2714 7172
rect 2586 6954 2622 7010
rect 2678 6954 2714 7010
rect 2586 6793 2714 6954
rect 2586 6737 2622 6793
rect 2678 6737 2714 6793
rect 2586 6698 2714 6737
rect 3100 7881 3228 7920
rect 3100 7825 3136 7881
rect 3192 7825 3228 7881
rect 3100 7664 3228 7825
rect 3100 7608 3136 7664
rect 3192 7608 3228 7664
rect 3100 7446 3228 7608
rect 3100 7390 3136 7446
rect 3192 7390 3228 7446
rect 3100 7228 3228 7390
rect 3100 7172 3136 7228
rect 3192 7172 3228 7228
rect 3100 7010 3228 7172
rect 3100 6954 3136 7010
rect 3192 6954 3228 7010
rect 3100 6793 3228 6954
rect 3100 6737 3136 6793
rect 3192 6737 3228 6793
rect 3100 6698 3228 6737
rect 3580 5820 3705 5859
rect 3580 5764 3615 5820
rect 3671 5764 3705 5820
rect 3580 5644 3705 5764
rect 2805 5574 2929 5614
rect 2805 5522 2841 5574
rect 2893 5522 2929 5574
rect 2805 5356 2929 5522
rect 3317 5574 3446 5614
rect 3317 5522 3355 5574
rect 3407 5522 3446 5574
rect 2805 5304 2841 5356
rect 2893 5304 2929 5356
rect 2805 5264 2929 5304
rect 3089 5344 3217 5383
rect 3089 5288 3125 5344
rect 3181 5288 3217 5344
rect 2366 3159 2404 3211
rect 2456 3159 2495 3211
rect 2366 2993 2495 3159
rect 2366 2946 2404 2993
rect 2368 2941 2404 2946
rect 2456 2946 2495 2993
rect 3089 5126 3217 5288
rect 3089 5070 3125 5126
rect 3181 5070 3217 5126
rect 3089 3000 3217 5070
rect 3317 5356 3446 5522
rect 3317 5304 3355 5356
rect 3407 5304 3446 5356
rect 3317 4576 3446 5304
rect 3316 4535 3446 4576
rect 3316 4483 3355 4535
rect 3407 4483 3446 4535
rect 3316 4463 3446 4483
rect 3578 5602 3707 5644
rect 3578 5546 3615 5602
rect 3671 5546 3707 5602
rect 3316 4442 3445 4463
rect 3578 3202 3707 5546
rect 4057 3211 4186 8050
rect 4277 7881 4405 7920
rect 4277 7825 4313 7881
rect 4369 7825 4405 7881
rect 4277 7664 4405 7825
rect 4277 7608 4313 7664
rect 4369 7608 4405 7664
rect 4277 7446 4405 7608
rect 4277 7390 4313 7446
rect 4369 7390 4405 7446
rect 4277 7228 4405 7390
rect 4277 7172 4313 7228
rect 4369 7172 4405 7228
rect 4277 7010 4405 7172
rect 4277 6954 4313 7010
rect 4369 6954 4405 7010
rect 4277 6793 4405 6954
rect 4277 6737 4313 6793
rect 4369 6737 4405 6793
rect 4277 6698 4405 6737
rect 4791 7881 4919 7920
rect 4791 7825 4827 7881
rect 4883 7825 4919 7881
rect 4791 7664 4919 7825
rect 4791 7608 4827 7664
rect 4883 7608 4919 7664
rect 4791 7446 4919 7608
rect 4791 7390 4827 7446
rect 4883 7390 4919 7446
rect 4791 7228 4919 7390
rect 4791 7172 4827 7228
rect 4883 7172 4919 7228
rect 4791 7010 4919 7172
rect 4791 6954 4827 7010
rect 4883 6954 4919 7010
rect 4791 6793 4919 6954
rect 4791 6737 4827 6793
rect 4883 6737 4919 6793
rect 4791 6698 4919 6737
rect 5271 5820 5396 5859
rect 5271 5764 5306 5820
rect 5362 5764 5396 5820
rect 5271 5644 5396 5764
rect 4494 5574 4623 5614
rect 4494 5522 4532 5574
rect 4584 5522 4623 5574
rect 4494 5356 4623 5522
rect 5008 5574 5137 5614
rect 5008 5522 5046 5574
rect 5098 5522 5137 5574
rect 4494 5304 4532 5356
rect 4584 5304 4623 5356
rect 4494 4939 4623 5304
rect 4494 4887 4533 4939
rect 4585 4887 4623 4939
rect 4494 4846 4623 4887
rect 4780 5344 4908 5383
rect 4780 5288 4816 5344
rect 4872 5288 4908 5344
rect 4780 5126 4908 5288
rect 4780 5070 4816 5126
rect 4872 5070 4908 5126
rect 4057 3159 4095 3211
rect 4147 3159 4186 3211
rect 2456 2941 2492 2946
rect 2368 2901 2492 2941
rect 3089 2867 3707 3000
rect 4057 2993 4186 3159
rect 4057 2946 4095 2993
rect 4059 2941 4095 2946
rect 4147 2946 4186 2993
rect 4780 3000 4908 5070
rect 5008 5356 5137 5522
rect 5008 5304 5046 5356
rect 5098 5304 5137 5356
rect 5008 4374 5137 5304
rect 5007 4333 5137 4374
rect 5007 4281 5046 4333
rect 5098 4281 5137 4333
rect 5007 4261 5137 4281
rect 5269 5602 5398 5644
rect 5269 5546 5306 5602
rect 5362 5546 5398 5602
rect 5007 4240 5136 4261
rect 5269 3202 5398 5546
rect 5748 3211 5877 8050
rect 5968 7881 6096 7920
rect 5968 7825 6004 7881
rect 6060 7825 6096 7881
rect 5968 7664 6096 7825
rect 5968 7608 6004 7664
rect 6060 7608 6096 7664
rect 5968 7446 6096 7608
rect 5968 7390 6004 7446
rect 6060 7390 6096 7446
rect 5968 7228 6096 7390
rect 5968 7172 6004 7228
rect 6060 7172 6096 7228
rect 5968 7010 6096 7172
rect 5968 6954 6004 7010
rect 6060 6954 6096 7010
rect 5968 6793 6096 6954
rect 5968 6737 6004 6793
rect 6060 6737 6096 6793
rect 5968 6698 6096 6737
rect 6482 7881 6610 7920
rect 6482 7825 6518 7881
rect 6574 7825 6610 7881
rect 6482 7664 6610 7825
rect 6482 7608 6518 7664
rect 6574 7608 6610 7664
rect 6482 7446 6610 7608
rect 6482 7390 6518 7446
rect 6574 7390 6610 7446
rect 6482 7228 6610 7390
rect 7633 7821 7761 7858
rect 7633 7765 7669 7821
rect 7725 7765 7761 7821
rect 7633 7603 7761 7765
rect 7633 7547 7669 7603
rect 7725 7547 7761 7603
rect 7633 7385 7761 7547
rect 7633 7329 7669 7385
rect 7725 7329 7761 7385
rect 7633 7291 7761 7329
rect 8081 7821 8209 7858
rect 8081 7765 8117 7821
rect 8173 7765 8209 7821
rect 8081 7603 8209 7765
rect 8081 7547 8117 7603
rect 8173 7547 8209 7603
rect 8081 7385 8209 7547
rect 8081 7329 8117 7385
rect 8173 7329 8209 7385
rect 8081 7291 8209 7329
rect 8529 7821 8657 7858
rect 8529 7765 8565 7821
rect 8621 7765 8657 7821
rect 8529 7603 8657 7765
rect 8529 7547 8565 7603
rect 8621 7547 8657 7603
rect 8529 7385 8657 7547
rect 8529 7329 8565 7385
rect 8621 7329 8657 7385
rect 8529 7291 8657 7329
rect 9266 7821 9394 7858
rect 9266 7765 9302 7821
rect 9358 7765 9394 7821
rect 9266 7603 9394 7765
rect 9266 7547 9302 7603
rect 9358 7547 9394 7603
rect 9266 7385 9394 7547
rect 9266 7329 9302 7385
rect 9358 7329 9394 7385
rect 9266 7291 9394 7329
rect 9714 7821 9842 7858
rect 9714 7765 9750 7821
rect 9806 7765 9842 7821
rect 9714 7603 9842 7765
rect 9714 7547 9750 7603
rect 9806 7547 9842 7603
rect 9714 7385 9842 7547
rect 9714 7329 9750 7385
rect 9806 7329 9842 7385
rect 9714 7291 9842 7329
rect 10162 7821 10290 7858
rect 10162 7765 10198 7821
rect 10254 7765 10290 7821
rect 10162 7603 10290 7765
rect 10162 7547 10198 7603
rect 10254 7547 10290 7603
rect 10162 7385 10290 7547
rect 10162 7329 10198 7385
rect 10254 7329 10290 7385
rect 10162 7291 10290 7329
rect 10900 7821 11028 7858
rect 10900 7765 10936 7821
rect 10992 7765 11028 7821
rect 10900 7603 11028 7765
rect 10900 7547 10936 7603
rect 10992 7547 11028 7603
rect 10900 7385 11028 7547
rect 10900 7329 10936 7385
rect 10992 7329 11028 7385
rect 10900 7291 11028 7329
rect 11348 7821 11476 7858
rect 11348 7765 11384 7821
rect 11440 7765 11476 7821
rect 11348 7603 11476 7765
rect 11348 7547 11384 7603
rect 11440 7547 11476 7603
rect 11348 7385 11476 7547
rect 11348 7329 11384 7385
rect 11440 7329 11476 7385
rect 11348 7291 11476 7329
rect 11796 7821 11924 7858
rect 11796 7765 11832 7821
rect 11888 7765 11924 7821
rect 11796 7603 11924 7765
rect 11796 7547 11832 7603
rect 11888 7547 11924 7603
rect 11796 7385 11924 7547
rect 11796 7329 11832 7385
rect 11888 7329 11924 7385
rect 11796 7291 11924 7329
rect 12534 7821 12662 7858
rect 12534 7765 12570 7821
rect 12626 7765 12662 7821
rect 12534 7603 12662 7765
rect 12534 7547 12570 7603
rect 12626 7547 12662 7603
rect 12534 7385 12662 7547
rect 12534 7329 12570 7385
rect 12626 7329 12662 7385
rect 12534 7291 12662 7329
rect 12982 7821 13110 7858
rect 12982 7765 13018 7821
rect 13074 7765 13110 7821
rect 12982 7603 13110 7765
rect 12982 7547 13018 7603
rect 13074 7547 13110 7603
rect 12982 7385 13110 7547
rect 12982 7329 13018 7385
rect 13074 7329 13110 7385
rect 12982 7291 13110 7329
rect 13430 7821 13558 7858
rect 13430 7765 13466 7821
rect 13522 7765 13558 7821
rect 13430 7603 13558 7765
rect 13430 7547 13466 7603
rect 13522 7547 13558 7603
rect 13430 7385 13558 7547
rect 13430 7329 13466 7385
rect 13522 7329 13558 7385
rect 13430 7291 13558 7329
rect 6482 7172 6518 7228
rect 6574 7172 6610 7228
rect 6482 7010 6610 7172
rect 6482 6954 6518 7010
rect 6574 6954 6610 7010
rect 6482 6793 6610 6954
rect 6482 6737 6518 6793
rect 6574 6737 6610 6793
rect 6482 6698 6610 6737
rect 7638 6711 7765 6750
rect 7638 6655 7673 6711
rect 7729 6655 7765 6711
rect 7638 6494 7765 6655
rect 7638 6438 7673 6494
rect 7729 6438 7765 6494
rect 7638 6276 7765 6438
rect 7638 6220 7673 6276
rect 7729 6220 7765 6276
rect 7638 6058 7765 6220
rect 7638 6002 7673 6058
rect 7729 6002 7765 6058
rect 6962 5820 7087 5859
rect 6962 5764 6997 5820
rect 7053 5764 7087 5820
rect 6962 5644 7087 5764
rect 7638 5841 7765 6002
rect 7638 5785 7673 5841
rect 7729 5785 7765 5841
rect 7638 5746 7765 5785
rect 8081 6712 8209 6749
rect 8081 6656 8117 6712
rect 8173 6656 8209 6712
rect 8081 6494 8209 6656
rect 8081 6438 8117 6494
rect 8173 6438 8209 6494
rect 8081 6277 8209 6438
rect 8081 6221 8117 6277
rect 8173 6221 8209 6277
rect 8081 6059 8209 6221
rect 8081 6003 8117 6059
rect 8173 6003 8209 6059
rect 8081 5841 8209 6003
rect 8081 5785 8117 5841
rect 8173 5785 8209 5841
rect 6185 5574 6314 5614
rect 6185 5522 6223 5574
rect 6275 5522 6314 5574
rect 6185 5356 6314 5522
rect 6701 5574 6825 5614
rect 6701 5522 6737 5574
rect 6789 5522 6825 5574
rect 6701 5383 6825 5522
rect 6960 5602 7089 5644
rect 6960 5546 6997 5602
rect 7053 5546 7089 5602
rect 6185 5304 6223 5356
rect 6275 5304 6314 5356
rect 6185 4778 6314 5304
rect 6184 4737 6314 4778
rect 6184 4685 6223 4737
rect 6275 4685 6314 4737
rect 6184 4665 6314 4685
rect 6471 5344 6599 5383
rect 6471 5288 6507 5344
rect 6563 5288 6599 5344
rect 6471 5126 6599 5288
rect 6471 5070 6507 5126
rect 6563 5070 6599 5126
rect 6184 4644 6313 4665
rect 5748 3159 5786 3211
rect 5838 3159 5877 3211
rect 4147 2941 4183 2946
rect 4059 2901 4183 2941
rect 4780 2867 5398 3000
rect 5748 2993 5877 3159
rect 5748 2946 5786 2993
rect 5750 2941 5786 2946
rect 5838 2946 5877 2993
rect 6471 3000 6599 5070
rect 6699 5356 6828 5383
rect 6699 5304 6737 5356
rect 6789 5304 6828 5356
rect 6699 4173 6828 5304
rect 6698 4132 6828 4173
rect 6698 4080 6737 4132
rect 6789 4080 6828 4132
rect 6698 4059 6828 4080
rect 6698 4039 6827 4059
rect 6960 3336 7089 5546
rect 7409 5604 7985 5644
rect 7409 5552 7447 5604
rect 7499 5552 7895 5604
rect 7947 5552 7985 5604
rect 7409 5386 7985 5552
rect 7409 5334 7447 5386
rect 7499 5334 7895 5386
rect 7947 5334 7985 5386
rect 7409 5293 7985 5334
rect 8081 5624 8209 5785
rect 8525 6711 8652 6750
rect 8525 6655 8561 6711
rect 8617 6655 8652 6711
rect 8525 6494 8652 6655
rect 8525 6438 8561 6494
rect 8617 6438 8652 6494
rect 8525 6276 8652 6438
rect 8525 6220 8561 6276
rect 8617 6220 8652 6276
rect 8525 6058 8652 6220
rect 8525 6002 8561 6058
rect 8617 6002 8652 6058
rect 8525 5841 8652 6002
rect 8525 5785 8561 5841
rect 8617 5785 8652 5841
rect 8525 5746 8652 5785
rect 9271 6711 9398 6750
rect 9271 6655 9306 6711
rect 9362 6655 9398 6711
rect 9271 6494 9398 6655
rect 9271 6438 9306 6494
rect 9362 6438 9398 6494
rect 9271 6276 9398 6438
rect 9271 6220 9306 6276
rect 9362 6220 9398 6276
rect 9271 6058 9398 6220
rect 9271 6002 9306 6058
rect 9362 6002 9398 6058
rect 9271 5841 9398 6002
rect 9271 5785 9306 5841
rect 9362 5785 9398 5841
rect 9271 5746 9398 5785
rect 9714 6712 9842 6749
rect 9714 6656 9750 6712
rect 9806 6656 9842 6712
rect 9714 6494 9842 6656
rect 9714 6438 9750 6494
rect 9806 6438 9842 6494
rect 9714 6277 9842 6438
rect 9714 6221 9750 6277
rect 9806 6221 9842 6277
rect 9714 6059 9842 6221
rect 9714 6003 9750 6059
rect 9806 6003 9842 6059
rect 9714 5841 9842 6003
rect 9714 5785 9750 5841
rect 9806 5785 9842 5841
rect 8081 5568 8117 5624
rect 8173 5568 8209 5624
rect 8081 5406 8209 5568
rect 8081 5350 8117 5406
rect 8173 5350 8209 5406
rect 8081 5312 8209 5350
rect 8305 5604 8881 5644
rect 8305 5552 8343 5604
rect 8395 5552 8791 5604
rect 8843 5552 8881 5604
rect 8305 5386 8881 5552
rect 8305 5334 8343 5386
rect 8395 5334 8791 5386
rect 8843 5334 8881 5386
rect 8305 5293 8881 5334
rect 7409 5292 7538 5293
rect 8752 5292 8881 5293
rect 7409 3712 7537 5292
rect 7409 3660 7447 3712
rect 7499 3660 7537 3712
rect 7409 3611 7537 3660
rect 7410 3495 7537 3611
rect 8753 3712 8881 5292
rect 8753 3660 8791 3712
rect 8843 3660 8881 3712
rect 8753 3611 8881 3660
rect 9042 5604 9618 5644
rect 9042 5552 9080 5604
rect 9132 5552 9528 5604
rect 9580 5552 9618 5604
rect 9042 5386 9618 5552
rect 9042 5334 9080 5386
rect 9132 5334 9528 5386
rect 9580 5334 9618 5386
rect 9042 5293 9618 5334
rect 9714 5624 9842 5785
rect 10158 6711 10285 6750
rect 10158 6655 10194 6711
rect 10250 6655 10285 6711
rect 10158 6494 10285 6655
rect 10158 6438 10194 6494
rect 10250 6438 10285 6494
rect 10158 6276 10285 6438
rect 10158 6220 10194 6276
rect 10250 6220 10285 6276
rect 10158 6058 10285 6220
rect 10158 6002 10194 6058
rect 10250 6002 10285 6058
rect 10158 5841 10285 6002
rect 10158 5785 10194 5841
rect 10250 5785 10285 5841
rect 10158 5746 10285 5785
rect 10905 6711 11032 6750
rect 10905 6655 10940 6711
rect 10996 6655 11032 6711
rect 10905 6494 11032 6655
rect 10905 6438 10940 6494
rect 10996 6438 11032 6494
rect 10905 6276 11032 6438
rect 10905 6220 10940 6276
rect 10996 6220 11032 6276
rect 10905 6058 11032 6220
rect 10905 6002 10940 6058
rect 10996 6002 11032 6058
rect 10905 5841 11032 6002
rect 10905 5785 10940 5841
rect 10996 5785 11032 5841
rect 10905 5746 11032 5785
rect 11348 6712 11476 6749
rect 11348 6656 11384 6712
rect 11440 6656 11476 6712
rect 11348 6494 11476 6656
rect 11348 6438 11384 6494
rect 11440 6438 11476 6494
rect 11348 6277 11476 6438
rect 11348 6221 11384 6277
rect 11440 6221 11476 6277
rect 11348 6059 11476 6221
rect 11348 6003 11384 6059
rect 11440 6003 11476 6059
rect 11348 5841 11476 6003
rect 11348 5785 11384 5841
rect 11440 5785 11476 5841
rect 9714 5568 9750 5624
rect 9806 5568 9842 5624
rect 9714 5406 9842 5568
rect 9714 5350 9750 5406
rect 9806 5350 9842 5406
rect 9714 5312 9842 5350
rect 9938 5604 10514 5644
rect 9938 5552 9976 5604
rect 10028 5552 10424 5604
rect 10476 5552 10514 5604
rect 9938 5386 10514 5552
rect 9938 5334 9976 5386
rect 10028 5334 10424 5386
rect 10476 5334 10514 5386
rect 9938 5293 10514 5334
rect 9042 5292 9171 5293
rect 10385 5292 10514 5293
rect 9042 3712 9170 5292
rect 9042 3660 9080 3712
rect 9132 3660 9170 3712
rect 9042 3611 9170 3660
rect 7410 3443 7447 3495
rect 7499 3443 7537 3495
rect 6960 3202 7309 3336
rect 5838 2941 5874 2946
rect 5750 2901 5874 2941
rect 6471 2867 7089 3000
rect 403 1117 537 1157
rect 403 1065 444 1117
rect 496 1065 537 1117
rect 403 899 537 1065
rect 403 847 444 899
rect 496 847 537 899
rect 403 -1293 537 847
rect 645 237 1086 1382
rect 645 185 733 237
rect 785 185 945 237
rect 997 185 1086 237
rect 645 19 1086 185
rect 645 -33 733 19
rect 785 -33 945 19
rect 997 -33 1086 19
rect 645 -126 1086 -33
rect 1231 1117 1361 1158
rect 1231 1065 1270 1117
rect 1322 1065 1361 1117
rect 1231 899 1361 1065
rect 1231 847 1270 899
rect 1322 847 1361 899
rect 1231 807 1361 847
rect 1472 1117 1602 1158
rect 1472 1065 1511 1117
rect 1563 1065 1602 1117
rect 1472 899 1602 1065
rect 1472 847 1511 899
rect 1563 847 1602 899
rect 1472 807 1602 847
rect 300 -1332 640 -1293
rect 300 -1388 336 -1332
rect 392 -1388 548 -1332
rect 604 -1388 640 -1332
rect 300 -1426 640 -1388
rect 403 -1427 537 -1426
rect 1231 -1427 1360 807
rect 1473 -1427 1602 807
rect 1714 1117 1844 1158
rect 1714 1065 1753 1117
rect 1805 1065 1844 1117
rect 1714 899 1844 1065
rect 1714 847 1753 899
rect 1805 847 1844 899
rect 1714 807 1844 847
rect 1714 -1427 1843 807
rect 3370 -1427 3504 1518
rect 5061 -1427 5195 1518
rect 6754 -1427 6888 1518
rect 7180 1427 7309 3202
rect 7410 3277 7537 3443
rect 7410 3225 7447 3277
rect 7499 3225 7537 3277
rect 7410 3059 7537 3225
rect 7410 3007 7447 3059
rect 7499 3007 7537 3059
rect 7410 2842 7537 3007
rect 7410 2790 7447 2842
rect 7499 2790 7537 2842
rect 7410 2749 7537 2790
rect 8107 3586 8183 3596
rect 8107 2594 8117 3586
rect 8173 2594 8183 3586
rect 8753 3495 8880 3611
rect 8753 3443 8791 3495
rect 8843 3443 8880 3495
rect 8753 3277 8880 3443
rect 8753 3225 8791 3277
rect 8843 3225 8880 3277
rect 8753 3059 8880 3225
rect 8753 3007 8791 3059
rect 8843 3007 8880 3059
rect 8753 2842 8880 3007
rect 8753 2790 8791 2842
rect 8843 2790 8880 2842
rect 8753 2749 8880 2790
rect 9043 3495 9170 3611
rect 10386 3712 10514 5292
rect 10386 3660 10424 3712
rect 10476 3660 10514 3712
rect 10386 3611 10514 3660
rect 10676 5604 11252 5644
rect 10676 5552 10714 5604
rect 10766 5552 11162 5604
rect 11214 5552 11252 5604
rect 10676 5386 11252 5552
rect 10676 5334 10714 5386
rect 10766 5334 11162 5386
rect 11214 5334 11252 5386
rect 10676 5293 11252 5334
rect 11348 5624 11476 5785
rect 11792 6711 11919 6750
rect 11792 6655 11828 6711
rect 11884 6655 11919 6711
rect 11792 6494 11919 6655
rect 11792 6438 11828 6494
rect 11884 6438 11919 6494
rect 11792 6276 11919 6438
rect 11792 6220 11828 6276
rect 11884 6220 11919 6276
rect 11792 6058 11919 6220
rect 11792 6002 11828 6058
rect 11884 6002 11919 6058
rect 11792 5841 11919 6002
rect 11792 5785 11828 5841
rect 11884 5785 11919 5841
rect 11792 5746 11919 5785
rect 12539 6711 12666 6750
rect 12539 6655 12574 6711
rect 12630 6655 12666 6711
rect 12539 6494 12666 6655
rect 12539 6438 12574 6494
rect 12630 6438 12666 6494
rect 12539 6276 12666 6438
rect 12539 6220 12574 6276
rect 12630 6220 12666 6276
rect 12539 6058 12666 6220
rect 12539 6002 12574 6058
rect 12630 6002 12666 6058
rect 12539 5841 12666 6002
rect 12539 5785 12574 5841
rect 12630 5785 12666 5841
rect 12539 5746 12666 5785
rect 12982 6712 13110 6749
rect 12982 6656 13018 6712
rect 13074 6656 13110 6712
rect 12982 6494 13110 6656
rect 12982 6438 13018 6494
rect 13074 6438 13110 6494
rect 12982 6277 13110 6438
rect 12982 6221 13018 6277
rect 13074 6221 13110 6277
rect 12982 6059 13110 6221
rect 12982 6003 13018 6059
rect 13074 6003 13110 6059
rect 12982 5841 13110 6003
rect 12982 5785 13018 5841
rect 13074 5785 13110 5841
rect 11348 5568 11384 5624
rect 11440 5568 11476 5624
rect 11348 5406 11476 5568
rect 11348 5350 11384 5406
rect 11440 5350 11476 5406
rect 11348 5312 11476 5350
rect 11572 5604 12148 5644
rect 11572 5552 11610 5604
rect 11662 5552 12058 5604
rect 12110 5552 12148 5604
rect 11572 5386 12148 5552
rect 11572 5334 11610 5386
rect 11662 5334 12058 5386
rect 12110 5334 12148 5386
rect 11572 5293 12148 5334
rect 10676 5292 10805 5293
rect 12019 5292 12148 5293
rect 10676 3712 10804 5292
rect 10676 3660 10714 3712
rect 10766 3660 10804 3712
rect 10676 3611 10804 3660
rect 9043 3443 9080 3495
rect 9132 3443 9170 3495
rect 9043 3277 9170 3443
rect 9043 3225 9080 3277
rect 9132 3225 9170 3277
rect 9043 3059 9170 3225
rect 9043 3007 9080 3059
rect 9132 3007 9170 3059
rect 9043 2842 9170 3007
rect 9043 2790 9080 2842
rect 9132 2790 9170 2842
rect 9043 2749 9170 2790
rect 9741 3586 9817 3596
rect 8107 2584 8183 2594
rect 9741 2594 9751 3586
rect 9807 2594 9817 3586
rect 10386 3495 10513 3611
rect 10386 3443 10424 3495
rect 10476 3443 10513 3495
rect 10386 3277 10513 3443
rect 10386 3225 10424 3277
rect 10476 3225 10513 3277
rect 10386 3059 10513 3225
rect 10386 3007 10424 3059
rect 10476 3007 10513 3059
rect 10386 2842 10513 3007
rect 10386 2790 10424 2842
rect 10476 2790 10513 2842
rect 10386 2749 10513 2790
rect 10677 3495 10804 3611
rect 12020 3712 12148 5292
rect 12020 3660 12058 3712
rect 12110 3660 12148 3712
rect 12020 3611 12148 3660
rect 12310 5604 12886 5644
rect 12310 5552 12348 5604
rect 12400 5552 12796 5604
rect 12848 5552 12886 5604
rect 12310 5386 12886 5552
rect 12310 5334 12348 5386
rect 12400 5334 12796 5386
rect 12848 5334 12886 5386
rect 12310 5293 12886 5334
rect 12982 5624 13110 5785
rect 13426 6711 13553 6750
rect 13426 6655 13462 6711
rect 13518 6655 13553 6711
rect 13426 6494 13553 6655
rect 13426 6438 13462 6494
rect 13518 6438 13553 6494
rect 13426 6276 13553 6438
rect 13426 6220 13462 6276
rect 13518 6220 13553 6276
rect 13426 6058 13553 6220
rect 13426 6002 13462 6058
rect 13518 6002 13553 6058
rect 13426 5841 13553 6002
rect 13426 5785 13462 5841
rect 13518 5785 13553 5841
rect 13426 5746 13553 5785
rect 12982 5568 13018 5624
rect 13074 5568 13110 5624
rect 12982 5406 13110 5568
rect 12982 5350 13018 5406
rect 13074 5350 13110 5406
rect 12982 5312 13110 5350
rect 13206 5604 13782 5644
rect 13206 5552 13244 5604
rect 13296 5552 13692 5604
rect 13744 5552 13782 5604
rect 13206 5386 13782 5552
rect 13206 5334 13244 5386
rect 13296 5334 13692 5386
rect 13744 5334 13782 5386
rect 13206 5293 13782 5334
rect 12310 5292 12439 5293
rect 13653 5292 13782 5293
rect 12310 3712 12438 5292
rect 12310 3660 12348 3712
rect 12400 3660 12438 3712
rect 12310 3611 12438 3660
rect 10677 3443 10714 3495
rect 10766 3443 10804 3495
rect 10677 3277 10804 3443
rect 10677 3225 10714 3277
rect 10766 3225 10804 3277
rect 10677 3059 10804 3225
rect 10677 3007 10714 3059
rect 10766 3007 10804 3059
rect 10677 2842 10804 3007
rect 10677 2790 10714 2842
rect 10766 2790 10804 2842
rect 10677 2749 10804 2790
rect 11374 3586 11450 3596
rect 9741 2584 9817 2594
rect 11374 2594 11384 3586
rect 11440 2594 11450 3586
rect 12020 3495 12147 3611
rect 12020 3443 12058 3495
rect 12110 3443 12147 3495
rect 12020 3277 12147 3443
rect 12020 3225 12058 3277
rect 12110 3225 12147 3277
rect 12020 3059 12147 3225
rect 12020 3007 12058 3059
rect 12110 3007 12147 3059
rect 12020 2842 12147 3007
rect 12020 2790 12058 2842
rect 12110 2790 12147 2842
rect 12020 2749 12147 2790
rect 12311 3495 12438 3611
rect 13654 3712 13782 5292
rect 13654 3660 13692 3712
rect 13744 3660 13782 3712
rect 13654 3611 13782 3660
rect 12311 3443 12348 3495
rect 12400 3443 12438 3495
rect 12311 3277 12438 3443
rect 12311 3225 12348 3277
rect 12400 3225 12438 3277
rect 12311 3059 12438 3225
rect 12311 3007 12348 3059
rect 12400 3007 12438 3059
rect 12311 2842 12438 3007
rect 12311 2790 12348 2842
rect 12400 2790 12438 2842
rect 12311 2749 12438 2790
rect 13008 3586 13084 3596
rect 11374 2584 11450 2594
rect 13008 2594 13018 3586
rect 13074 2594 13084 3586
rect 13654 3495 13781 3611
rect 13654 3443 13692 3495
rect 13744 3443 13781 3495
rect 13654 3277 13781 3443
rect 13654 3225 13692 3277
rect 13744 3225 13781 3277
rect 13654 3059 13781 3225
rect 13654 3007 13692 3059
rect 13744 3007 13781 3059
rect 13654 2842 13781 3007
rect 13654 2790 13692 2842
rect 13744 2790 13781 2842
rect 13654 2749 13781 2790
rect 13008 2584 13084 2594
rect 9861 2010 13574 2048
rect 8963 1926 9092 1966
rect 7802 1878 7927 1917
rect 7802 1822 7836 1878
rect 7892 1822 7927 1878
rect 7802 1660 7927 1822
rect 8963 1874 9001 1926
rect 9053 1874 9092 1926
rect 8963 1749 9092 1874
rect 7802 1604 7836 1660
rect 7892 1604 7927 1660
rect 7802 1566 7927 1604
rect 8133 1708 9092 1749
rect 8133 1656 9001 1708
rect 9053 1656 9092 1708
rect 9861 1954 9898 2010
rect 9954 1954 10109 2010
rect 10165 1954 10319 2010
rect 10375 1954 10530 2010
rect 10586 1954 10741 2010
rect 10797 1954 10952 2010
rect 11008 1954 11163 2010
rect 11219 1954 11373 2010
rect 11429 1954 11584 2010
rect 11640 1954 11796 2010
rect 11852 1954 12007 2010
rect 12063 1954 12217 2010
rect 12273 1954 12428 2010
rect 12484 1954 12639 2010
rect 12695 1954 12850 2010
rect 12906 1954 13061 2010
rect 13117 1954 13271 2010
rect 13327 1954 13482 2010
rect 13538 1954 13574 2010
rect 9861 1792 13574 1954
rect 9861 1736 9898 1792
rect 9954 1736 10109 1792
rect 10165 1736 10319 1792
rect 10375 1736 10530 1792
rect 10586 1736 10741 1792
rect 10797 1736 10952 1792
rect 11008 1736 11163 1792
rect 11219 1736 11373 1792
rect 11429 1736 11584 1792
rect 11640 1736 11796 1792
rect 11852 1736 12007 1792
rect 12063 1736 12217 1792
rect 12273 1736 12428 1792
rect 12484 1736 12639 1792
rect 12695 1736 12850 1792
rect 12906 1736 13061 1792
rect 13117 1736 13271 1792
rect 13327 1736 13482 1792
rect 13538 1736 13574 1792
rect 9861 1697 13574 1736
rect 8133 1615 9092 1656
rect 7180 1375 7218 1427
rect 7270 1375 7309 1427
rect 7180 1209 7309 1375
rect 7180 1157 7218 1209
rect 7270 1157 7309 1209
rect 7180 1117 7309 1157
rect 7411 1162 7536 1201
rect 7411 1106 7445 1162
rect 7501 1106 7536 1162
rect 7411 944 7536 1106
rect 7411 888 7445 944
rect 7501 888 7536 944
rect 7411 850 7536 888
rect 8133 -1293 8262 1615
rect 16247 1595 16375 1651
rect 8630 1451 9885 1463
rect 8630 1399 8642 1451
rect 8902 1399 9613 1451
rect 9873 1399 9885 1451
rect 8630 1387 9885 1399
rect 8438 1180 8563 1219
rect 8438 1124 8472 1180
rect 8528 1124 8563 1180
rect 8438 962 8563 1124
rect 8438 906 8472 962
rect 8528 906 8563 962
rect 8438 868 8563 906
rect 8880 289 9220 1387
rect 9622 1175 13546 1214
rect 9622 1119 9658 1175
rect 9714 1119 9869 1175
rect 9925 1119 10080 1175
rect 10136 1119 10291 1175
rect 10347 1119 10502 1175
rect 10558 1119 10712 1175
rect 10768 1119 10923 1175
rect 10979 1119 11134 1175
rect 11190 1119 11345 1175
rect 11401 1119 11556 1175
rect 11612 1119 11767 1175
rect 11823 1119 11978 1175
rect 12034 1119 12189 1175
rect 12245 1119 12400 1175
rect 12456 1119 12610 1175
rect 12666 1119 12821 1175
rect 12877 1119 13032 1175
rect 13088 1119 13243 1175
rect 13299 1119 13454 1175
rect 13510 1119 13546 1175
rect 9622 957 13546 1119
rect 9622 901 9658 957
rect 9714 901 9869 957
rect 9925 901 10080 957
rect 10136 901 10291 957
rect 10347 901 10502 957
rect 10558 901 10712 957
rect 10768 901 10923 957
rect 10979 901 11134 957
rect 11190 901 11345 957
rect 11401 901 11556 957
rect 11612 901 11767 957
rect 11823 901 11978 957
rect 12034 901 12189 957
rect 12245 901 12400 957
rect 12456 901 12610 957
rect 12666 901 12821 957
rect 12877 901 13032 957
rect 13088 901 13243 957
rect 13299 901 13454 957
rect 13510 901 13546 957
rect 9622 863 13546 901
rect 8880 237 8918 289
rect 8970 237 9130 289
rect 9182 237 9220 289
rect 8880 71 9220 237
rect 8880 19 8918 71
rect 8970 19 9130 71
rect 9182 19 9220 71
rect 8880 -21 9220 19
rect 8028 -1332 8368 -1293
rect 8028 -1388 8064 -1332
rect 8120 -1388 8276 -1332
rect 8332 -1388 8368 -1332
rect 8028 -1426 8368 -1388
rect 8133 -1427 8262 -1426
rect 16319 -1833 16375 1595
rect 21612 879 21965 3456
rect 28532 1382 29412 9334
rect 21612 615 21660 879
rect 21924 615 21965 879
rect 28007 1130 28136 1171
rect 28007 1078 28045 1130
rect 28097 1078 28136 1130
rect 28007 912 28136 1078
rect 28007 860 28045 912
rect 28097 860 28136 912
rect 28007 694 28136 860
rect 28007 642 28045 694
rect 28097 642 28136 694
rect 21612 -189 21965 615
rect 21612 -453 21660 -189
rect 21924 -453 21965 -189
rect 21612 -548 21965 -453
rect 22855 -1427 22989 618
rect 28007 -1427 28136 642
rect 28248 1130 28378 1171
rect 28248 1078 28287 1130
rect 28339 1078 28378 1130
rect 28248 912 28378 1078
rect 28248 860 28287 912
rect 28339 860 28378 912
rect 28248 694 28378 860
rect 28248 642 28287 694
rect 28339 642 28378 694
rect 28248 -1427 28378 642
rect 28490 1130 28619 1171
rect 28490 1078 28529 1130
rect 28581 1078 28619 1130
rect 28490 912 28619 1078
rect 28490 860 28529 912
rect 28581 860 28619 912
rect 28490 694 28619 860
rect 28490 642 28529 694
rect 28581 642 28619 694
rect 28490 -1427 28619 642
rect 28731 1130 28861 1171
rect 28731 1078 28770 1130
rect 28822 1078 28861 1130
rect 28731 912 28861 1078
rect 28731 860 28770 912
rect 28822 860 28861 912
rect 28731 694 28861 860
rect 28731 642 28770 694
rect 28822 642 28861 694
rect 28731 -1427 28861 642
rect 28971 237 29412 1382
rect 28971 185 29059 237
rect 29111 185 29271 237
rect 29323 185 29412 237
rect 28971 19 29412 185
rect 28971 -33 29059 19
rect 29111 -33 29271 19
rect 29323 -33 29412 19
rect 28971 -126 29412 -33
rect 29520 1117 29654 1157
rect 29520 1065 29561 1117
rect 29613 1065 29654 1117
rect 29520 899 29654 1065
rect 29520 847 29561 899
rect 29613 847 29654 899
rect 29520 -1293 29654 847
rect 29417 -1332 29757 -1293
rect 29417 -1388 29453 -1332
rect 29509 -1388 29665 -1332
rect 29721 -1388 29757 -1332
rect 29417 -1426 29757 -1388
rect 29520 -1427 29654 -1426
<< via2 >>
rect 740 29970 796 30026
rect 951 29970 1007 30026
rect 1163 29970 1219 30026
rect 1374 29970 1430 30026
rect 740 29752 796 29808
rect 951 29752 1007 29808
rect 1163 29752 1219 29808
rect 1374 29752 1430 29808
rect 740 29534 796 29590
rect 951 29534 1007 29590
rect 1163 29534 1219 29590
rect 1374 29534 1430 29590
rect 740 29316 796 29372
rect 951 29316 1007 29372
rect 1163 29316 1219 29372
rect 1374 29316 1430 29372
rect 442 28996 498 28998
rect 442 28944 444 28996
rect 444 28944 496 28996
rect 496 28944 498 28996
rect 442 28942 498 28944
rect 442 28778 498 28780
rect 442 28726 444 28778
rect 444 28726 496 28778
rect 496 28726 498 28778
rect 442 28724 498 28726
rect 5479 29970 5535 30026
rect 5691 29970 5747 30026
rect 5479 29752 5535 29808
rect 5691 29752 5747 29808
rect 5479 29534 5535 29590
rect 5691 29534 5747 29590
rect 5479 29316 5535 29372
rect 5691 29316 5747 29372
rect 1654 28500 1710 28502
rect 1654 28448 1656 28500
rect 1656 28448 1708 28500
rect 1708 28448 1710 28500
rect 1654 28446 1710 28448
rect 1654 28282 1710 28284
rect 1654 28230 1656 28282
rect 1656 28230 1708 28282
rect 1708 28230 1710 28282
rect 1654 28228 1710 28230
rect 1654 28064 1710 28066
rect 1654 28012 1656 28064
rect 1656 28012 1708 28064
rect 1708 28012 1710 28064
rect 1654 28010 1710 28012
rect 1654 27846 1710 27848
rect 1654 27794 1656 27846
rect 1656 27794 1708 27846
rect 1708 27794 1710 27846
rect 1654 27792 1710 27794
rect 2094 28500 2150 28502
rect 2094 28448 2096 28500
rect 2096 28448 2148 28500
rect 2148 28448 2150 28500
rect 2094 28446 2150 28448
rect 2094 28282 2150 28284
rect 2094 28230 2096 28282
rect 2096 28230 2148 28282
rect 2148 28230 2150 28282
rect 2094 28228 2150 28230
rect 2094 28064 2150 28066
rect 2094 28012 2096 28064
rect 2096 28012 2148 28064
rect 2148 28012 2150 28064
rect 2094 28010 2150 28012
rect 2094 27846 2150 27848
rect 2094 27794 2096 27846
rect 2096 27794 2148 27846
rect 2148 27794 2150 27846
rect 2094 27792 2150 27794
rect 3006 28500 3062 28502
rect 3006 28448 3008 28500
rect 3008 28448 3060 28500
rect 3060 28448 3062 28500
rect 3006 28446 3062 28448
rect 3006 28282 3062 28284
rect 3006 28230 3008 28282
rect 3008 28230 3060 28282
rect 3060 28230 3062 28282
rect 3006 28228 3062 28230
rect 3006 28064 3062 28066
rect 3006 28012 3008 28064
rect 3008 28012 3060 28064
rect 3060 28012 3062 28064
rect 3006 28010 3062 28012
rect 3006 27846 3062 27848
rect 3006 27794 3008 27846
rect 3008 27794 3060 27846
rect 3060 27794 3062 27846
rect 3006 27792 3062 27794
rect 3446 28500 3502 28502
rect 3446 28448 3448 28500
rect 3448 28448 3500 28500
rect 3500 28448 3502 28500
rect 3446 28446 3502 28448
rect 3446 28282 3502 28284
rect 3446 28230 3448 28282
rect 3448 28230 3500 28282
rect 3500 28230 3502 28282
rect 3446 28228 3502 28230
rect 3446 28064 3502 28066
rect 3446 28012 3448 28064
rect 3448 28012 3500 28064
rect 3500 28012 3502 28064
rect 3446 28010 3502 28012
rect 3446 27846 3502 27848
rect 3446 27794 3448 27846
rect 3448 27794 3500 27846
rect 3500 27794 3502 27846
rect 3446 27792 3502 27794
rect 3886 28500 3942 28502
rect 3886 28448 3888 28500
rect 3888 28448 3940 28500
rect 3940 28448 3942 28500
rect 3886 28446 3942 28448
rect 3886 28282 3942 28284
rect 3886 28230 3888 28282
rect 3888 28230 3940 28282
rect 3940 28230 3942 28282
rect 3886 28228 3942 28230
rect 3886 28064 3942 28066
rect 3886 28012 3888 28064
rect 3888 28012 3940 28064
rect 3940 28012 3942 28064
rect 3886 28010 3942 28012
rect 3886 27846 3942 27848
rect 3886 27794 3888 27846
rect 3888 27794 3940 27846
rect 3940 27794 3942 27846
rect 3886 27792 3942 27794
rect 4798 28500 4854 28502
rect 4798 28448 4800 28500
rect 4800 28448 4852 28500
rect 4852 28448 4854 28500
rect 4798 28446 4854 28448
rect 4798 28282 4854 28284
rect 4798 28230 4800 28282
rect 4800 28230 4852 28282
rect 4852 28230 4854 28282
rect 4798 28228 4854 28230
rect 4798 28064 4854 28066
rect 4798 28012 4800 28064
rect 4800 28012 4852 28064
rect 4852 28012 4854 28064
rect 4798 28010 4854 28012
rect 4798 27846 4854 27848
rect 4798 27794 4800 27846
rect 4800 27794 4852 27846
rect 4852 27794 4854 27846
rect 4798 27792 4854 27794
rect 5238 28500 5294 28502
rect 5238 28448 5240 28500
rect 5240 28448 5292 28500
rect 5292 28448 5294 28500
rect 5238 28446 5294 28448
rect 5238 28282 5294 28284
rect 5238 28230 5240 28282
rect 5240 28230 5292 28282
rect 5292 28230 5294 28282
rect 5238 28228 5294 28230
rect 5238 28064 5294 28066
rect 5238 28012 5240 28064
rect 5240 28012 5292 28064
rect 5292 28012 5294 28064
rect 5238 28010 5294 28012
rect 5238 27846 5294 27848
rect 5238 27794 5240 27846
rect 5240 27794 5292 27846
rect 5292 27794 5294 27846
rect 5238 27792 5294 27794
rect 16395 29970 16451 30026
rect 16607 29970 16663 30026
rect 16395 29752 16451 29808
rect 16607 29752 16663 29808
rect 16395 29534 16451 29590
rect 16607 29534 16663 29590
rect 16395 29316 16451 29372
rect 16607 29316 16663 29372
rect 6580 28943 6636 28999
rect 6580 28725 6636 28781
rect 13958 28943 14014 28999
rect 23343 29970 23399 30026
rect 23555 29970 23611 30026
rect 23343 29752 23399 29808
rect 23555 29752 23611 29808
rect 23343 29534 23399 29590
rect 23555 29534 23611 29590
rect 23343 29316 23399 29372
rect 23555 29316 23611 29372
rect 5921 28401 5977 28403
rect 5921 28349 5923 28401
rect 5923 28349 5975 28401
rect 5975 28349 5977 28401
rect 5921 28347 5977 28349
rect 5921 28183 5977 28185
rect 5921 28131 5923 28183
rect 5923 28131 5975 28183
rect 5975 28131 5977 28183
rect 5921 28129 5977 28131
rect 5921 27965 5977 27967
rect 5921 27913 5923 27965
rect 5923 27913 5975 27965
rect 5975 27913 5977 27965
rect 5921 27911 5977 27913
rect 6360 28401 6416 28403
rect 6360 28349 6362 28401
rect 6362 28349 6414 28401
rect 6414 28349 6416 28401
rect 6360 28347 6416 28349
rect 6360 28183 6416 28185
rect 6360 28131 6362 28183
rect 6362 28131 6414 28183
rect 6414 28131 6416 28183
rect 6360 28129 6416 28131
rect 6360 27965 6416 27967
rect 6360 27913 6362 27965
rect 6362 27913 6414 27965
rect 6414 27913 6416 27965
rect 6360 27911 6416 27913
rect 9033 28500 9089 28502
rect 9033 28448 9035 28500
rect 9035 28448 9087 28500
rect 9087 28448 9089 28500
rect 9033 28446 9089 28448
rect 7744 28344 7800 28346
rect 7744 28292 7746 28344
rect 7746 28292 7798 28344
rect 7798 28292 7800 28344
rect 7744 28290 7800 28292
rect 7744 28126 7800 28128
rect 7744 28074 7746 28126
rect 7746 28074 7798 28126
rect 7798 28074 7800 28126
rect 7744 28072 7800 28074
rect 7744 27908 7800 27910
rect 7744 27856 7746 27908
rect 7746 27856 7798 27908
rect 7798 27856 7800 27908
rect 7744 27854 7800 27856
rect 9033 28282 9089 28284
rect 9033 28230 9035 28282
rect 9035 28230 9087 28282
rect 9087 28230 9089 28282
rect 9033 28228 9089 28230
rect 9033 28064 9089 28066
rect 9033 28012 9035 28064
rect 9035 28012 9087 28064
rect 9087 28012 9089 28064
rect 9033 28010 9089 28012
rect 9033 27846 9089 27848
rect 9033 27794 9035 27846
rect 9035 27794 9087 27846
rect 9087 27794 9089 27846
rect 9033 27792 9089 27794
rect 9473 28500 9529 28502
rect 9473 28448 9475 28500
rect 9475 28448 9527 28500
rect 9527 28448 9529 28500
rect 9473 28446 9529 28448
rect 9473 28282 9529 28284
rect 9473 28230 9475 28282
rect 9475 28230 9527 28282
rect 9527 28230 9529 28282
rect 9473 28228 9529 28230
rect 9473 28064 9529 28066
rect 9473 28012 9475 28064
rect 9475 28012 9527 28064
rect 9527 28012 9529 28064
rect 9473 28010 9529 28012
rect 9473 27846 9529 27848
rect 9473 27794 9475 27846
rect 9475 27794 9527 27846
rect 9527 27794 9529 27846
rect 9473 27792 9529 27794
rect 10385 28500 10441 28502
rect 10385 28448 10387 28500
rect 10387 28448 10439 28500
rect 10439 28448 10441 28500
rect 10385 28446 10441 28448
rect 10385 28282 10441 28284
rect 10385 28230 10387 28282
rect 10387 28230 10439 28282
rect 10439 28230 10441 28282
rect 10385 28228 10441 28230
rect 10385 28064 10441 28066
rect 10385 28012 10387 28064
rect 10387 28012 10439 28064
rect 10439 28012 10441 28064
rect 10385 28010 10441 28012
rect 10385 27846 10441 27848
rect 10385 27794 10387 27846
rect 10387 27794 10439 27846
rect 10439 27794 10441 27846
rect 10385 27792 10441 27794
rect 10825 28500 10881 28502
rect 10825 28448 10827 28500
rect 10827 28448 10879 28500
rect 10879 28448 10881 28500
rect 10825 28446 10881 28448
rect 10825 28282 10881 28284
rect 10825 28230 10827 28282
rect 10827 28230 10879 28282
rect 10879 28230 10881 28282
rect 10825 28228 10881 28230
rect 10825 28064 10881 28066
rect 10825 28012 10827 28064
rect 10827 28012 10879 28064
rect 10879 28012 10881 28064
rect 10825 28010 10881 28012
rect 10825 27846 10881 27848
rect 10825 27794 10827 27846
rect 10827 27794 10879 27846
rect 10879 27794 10881 27846
rect 10825 27792 10881 27794
rect 11265 28500 11321 28502
rect 11265 28448 11267 28500
rect 11267 28448 11319 28500
rect 11319 28448 11321 28500
rect 11265 28446 11321 28448
rect 11265 28282 11321 28284
rect 11265 28230 11267 28282
rect 11267 28230 11319 28282
rect 11319 28230 11321 28282
rect 11265 28228 11321 28230
rect 11265 28064 11321 28066
rect 11265 28012 11267 28064
rect 11267 28012 11319 28064
rect 11319 28012 11321 28064
rect 11265 28010 11321 28012
rect 11265 27846 11321 27848
rect 11265 27794 11267 27846
rect 11267 27794 11319 27846
rect 11319 27794 11321 27846
rect 11265 27792 11321 27794
rect 13958 28725 14014 28781
rect 12177 28500 12233 28502
rect 12177 28448 12179 28500
rect 12179 28448 12231 28500
rect 12231 28448 12233 28500
rect 12177 28446 12233 28448
rect 12177 28282 12233 28284
rect 12177 28230 12179 28282
rect 12179 28230 12231 28282
rect 12231 28230 12233 28282
rect 12177 28228 12233 28230
rect 12177 28064 12233 28066
rect 12177 28012 12179 28064
rect 12179 28012 12231 28064
rect 12231 28012 12233 28064
rect 12177 28010 12233 28012
rect 12177 27846 12233 27848
rect 12177 27794 12179 27846
rect 12179 27794 12231 27846
rect 12231 27794 12233 27846
rect 12177 27792 12233 27794
rect 12617 28500 12673 28502
rect 12617 28448 12619 28500
rect 12619 28448 12671 28500
rect 12671 28448 12673 28500
rect 12617 28446 12673 28448
rect 12617 28282 12673 28284
rect 12617 28230 12619 28282
rect 12619 28230 12671 28282
rect 12671 28230 12673 28282
rect 12617 28228 12673 28230
rect 12617 28064 12673 28066
rect 12617 28012 12619 28064
rect 12619 28012 12671 28064
rect 12671 28012 12673 28064
rect 12617 28010 12673 28012
rect 13300 28401 13356 28403
rect 13300 28349 13302 28401
rect 13302 28349 13354 28401
rect 13354 28349 13356 28401
rect 13300 28347 13356 28349
rect 13300 28183 13356 28185
rect 13300 28131 13302 28183
rect 13302 28131 13354 28183
rect 13354 28131 13356 28183
rect 13300 28129 13356 28131
rect 13300 27965 13356 27967
rect 13300 27913 13302 27965
rect 13302 27913 13354 27965
rect 13354 27913 13356 27965
rect 13300 27911 13356 27913
rect 13739 28401 13795 28403
rect 13739 28349 13741 28401
rect 13741 28349 13793 28401
rect 13793 28349 13795 28401
rect 13739 28347 13795 28349
rect 13739 28183 13795 28185
rect 13739 28131 13741 28183
rect 13741 28131 13793 28183
rect 13793 28131 13795 28183
rect 13739 28129 13795 28131
rect 13739 27965 13795 27967
rect 13739 27913 13741 27965
rect 13741 27913 13793 27965
rect 13793 27913 13795 27965
rect 13739 27911 13795 27913
rect 12617 27846 12673 27848
rect 12617 27794 12619 27846
rect 12619 27794 12671 27846
rect 12671 27794 12673 27846
rect 12617 27792 12673 27794
rect 15123 28344 15179 28346
rect 15123 28292 15125 28344
rect 15125 28292 15177 28344
rect 15177 28292 15179 28344
rect 15123 28290 15179 28292
rect 15123 28126 15179 28128
rect 15123 28074 15125 28126
rect 15125 28074 15177 28126
rect 15177 28074 15179 28126
rect 15123 28072 15179 28074
rect 15123 27908 15179 27910
rect 15123 27856 15125 27908
rect 15125 27856 15177 27908
rect 15177 27856 15179 27908
rect 15123 27854 15179 27856
rect 16916 28392 16972 28394
rect 16916 28340 16918 28392
rect 16918 28340 16970 28392
rect 16970 28340 16972 28392
rect 16916 28338 16972 28340
rect 16916 28174 16972 28176
rect 16916 28122 16918 28174
rect 16918 28122 16970 28174
rect 16970 28122 16972 28174
rect 16916 28120 16972 28122
rect 16916 27956 16972 27958
rect 16916 27904 16918 27956
rect 16918 27904 16970 27956
rect 16970 27904 16972 27956
rect 16916 27902 16972 27904
rect 16916 27738 16972 27740
rect 16916 27686 16918 27738
rect 16918 27686 16970 27738
rect 16970 27686 16972 27738
rect 16916 27684 16972 27686
rect 1654 27353 1710 27355
rect 1654 27301 1656 27353
rect 1656 27301 1708 27353
rect 1708 27301 1710 27353
rect 1654 27299 1710 27301
rect 1654 27135 1710 27137
rect 1654 27083 1656 27135
rect 1656 27083 1708 27135
rect 1708 27083 1710 27135
rect 1654 27081 1710 27083
rect 1654 26917 1710 26919
rect 1654 26865 1656 26917
rect 1656 26865 1708 26917
rect 1708 26865 1710 26917
rect 1654 26863 1710 26865
rect 2102 27353 2158 27355
rect 2102 27301 2104 27353
rect 2104 27301 2156 27353
rect 2156 27301 2158 27353
rect 2102 27299 2158 27301
rect 2102 27135 2158 27137
rect 2102 27083 2104 27135
rect 2104 27083 2156 27135
rect 2156 27083 2158 27135
rect 2102 27081 2158 27083
rect 2102 26917 2158 26919
rect 2102 26865 2104 26917
rect 2104 26865 2156 26917
rect 2156 26865 2158 26917
rect 2102 26863 2158 26865
rect 2550 27353 2606 27355
rect 2550 27301 2552 27353
rect 2552 27301 2604 27353
rect 2604 27301 2606 27353
rect 2550 27299 2606 27301
rect 2550 27135 2606 27137
rect 2550 27083 2552 27135
rect 2552 27083 2604 27135
rect 2604 27083 2606 27135
rect 2550 27081 2606 27083
rect 2550 26917 2606 26919
rect 2550 26865 2552 26917
rect 2552 26865 2604 26917
rect 2604 26865 2606 26917
rect 2550 26863 2606 26865
rect 2998 27353 3054 27355
rect 2998 27301 3000 27353
rect 3000 27301 3052 27353
rect 3052 27301 3054 27353
rect 2998 27299 3054 27301
rect 2998 27135 3054 27137
rect 2998 27083 3000 27135
rect 3000 27083 3052 27135
rect 3052 27083 3054 27135
rect 2998 27081 3054 27083
rect 2998 26917 3054 26919
rect 2998 26865 3000 26917
rect 3000 26865 3052 26917
rect 3052 26865 3054 26917
rect 2998 26863 3054 26865
rect 3446 27353 3502 27355
rect 3446 27301 3448 27353
rect 3448 27301 3500 27353
rect 3500 27301 3502 27353
rect 3446 27299 3502 27301
rect 3446 27135 3502 27137
rect 3446 27083 3448 27135
rect 3448 27083 3500 27135
rect 3500 27083 3502 27135
rect 3446 27081 3502 27083
rect 3446 26917 3502 26919
rect 3446 26865 3448 26917
rect 3448 26865 3500 26917
rect 3500 26865 3502 26917
rect 3446 26863 3502 26865
rect 3894 27353 3950 27355
rect 3894 27301 3896 27353
rect 3896 27301 3948 27353
rect 3948 27301 3950 27353
rect 3894 27299 3950 27301
rect 3894 27135 3950 27137
rect 3894 27083 3896 27135
rect 3896 27083 3948 27135
rect 3948 27083 3950 27135
rect 3894 27081 3950 27083
rect 3894 26917 3950 26919
rect 3894 26865 3896 26917
rect 3896 26865 3948 26917
rect 3948 26865 3950 26917
rect 3894 26863 3950 26865
rect 4342 27353 4398 27355
rect 4342 27301 4344 27353
rect 4344 27301 4396 27353
rect 4396 27301 4398 27353
rect 4342 27299 4398 27301
rect 4342 27135 4398 27137
rect 4342 27083 4344 27135
rect 4344 27083 4396 27135
rect 4396 27083 4398 27135
rect 4342 27081 4398 27083
rect 4342 26917 4398 26919
rect 4342 26865 4344 26917
rect 4344 26865 4396 26917
rect 4396 26865 4398 26917
rect 4342 26863 4398 26865
rect 4790 27353 4846 27355
rect 4790 27301 4792 27353
rect 4792 27301 4844 27353
rect 4844 27301 4846 27353
rect 4790 27299 4846 27301
rect 4790 27135 4846 27137
rect 4790 27083 4792 27135
rect 4792 27083 4844 27135
rect 4844 27083 4846 27135
rect 4790 27081 4846 27083
rect 4790 26917 4846 26919
rect 4790 26865 4792 26917
rect 4792 26865 4844 26917
rect 4844 26865 4846 26917
rect 4790 26863 4846 26865
rect 5238 27353 5294 27355
rect 5238 27301 5240 27353
rect 5240 27301 5292 27353
rect 5292 27301 5294 27353
rect 5238 27299 5294 27301
rect 5238 27135 5294 27137
rect 5238 27083 5240 27135
rect 5240 27083 5292 27135
rect 5292 27083 5294 27135
rect 5238 27081 5294 27083
rect 5238 26917 5294 26919
rect 5238 26865 5240 26917
rect 5240 26865 5292 26917
rect 5292 26865 5294 26917
rect 5238 26863 5294 26865
rect 5645 27378 5701 27380
rect 5645 27326 5647 27378
rect 5647 27326 5699 27378
rect 5699 27326 5701 27378
rect 5645 27324 5701 27326
rect 5645 27160 5701 27162
rect 5645 27108 5647 27160
rect 5647 27108 5699 27160
rect 5699 27108 5701 27160
rect 5645 27106 5701 27108
rect 5645 26888 5701 26944
rect 5921 27378 5977 27380
rect 5921 27326 5923 27378
rect 5923 27326 5975 27378
rect 5975 27326 5977 27378
rect 5921 27324 5977 27326
rect 8134 27392 8190 27394
rect 8134 27340 8136 27392
rect 8136 27340 8188 27392
rect 8188 27340 8190 27392
rect 8134 27338 8190 27340
rect 5921 27160 5977 27162
rect 5921 27108 5923 27160
rect 5923 27108 5975 27160
rect 5975 27108 5977 27160
rect 5921 27106 5977 27108
rect 7005 27210 7061 27212
rect 7005 27158 7007 27210
rect 7007 27158 7059 27210
rect 7059 27158 7061 27210
rect 7005 27156 7061 27158
rect 7217 27210 7273 27212
rect 7217 27158 7219 27210
rect 7219 27158 7271 27210
rect 7271 27158 7273 27210
rect 7217 27156 7273 27158
rect 8134 27174 8190 27176
rect 8134 27122 8136 27174
rect 8136 27122 8188 27174
rect 8188 27122 8190 27174
rect 8134 27120 8190 27122
rect 5921 26888 5977 26944
rect 8134 26902 8190 26958
rect 5872 26514 5928 26516
rect 5872 26462 5874 26514
rect 5874 26462 5926 26514
rect 5926 26462 5928 26514
rect 5872 26460 5928 26462
rect 6079 26514 6135 26516
rect 6079 26462 6081 26514
rect 6081 26462 6133 26514
rect 6133 26462 6135 26514
rect 6079 26460 6135 26462
rect 5872 26296 5928 26298
rect 5872 26244 5874 26296
rect 5874 26244 5926 26296
rect 5926 26244 5928 26296
rect 5872 26242 5928 26244
rect 6079 26296 6135 26298
rect 6079 26244 6081 26296
rect 6081 26244 6133 26296
rect 6133 26244 6135 26296
rect 6079 26242 6135 26244
rect 5872 26078 5928 26080
rect 5872 26026 5874 26078
rect 5874 26026 5926 26078
rect 5926 26026 5928 26078
rect 5872 26024 5928 26026
rect 6079 26078 6135 26080
rect 6079 26026 6081 26078
rect 6081 26026 6133 26078
rect 6133 26026 6135 26078
rect 6079 26024 6135 26026
rect 5872 25860 5928 25862
rect 5872 25808 5874 25860
rect 5874 25808 5926 25860
rect 5926 25808 5928 25860
rect 5872 25806 5928 25808
rect 6079 25860 6135 25862
rect 6079 25808 6081 25860
rect 6081 25808 6133 25860
rect 6133 25808 6135 25860
rect 6079 25806 6135 25808
rect 6599 26491 6655 26493
rect 6599 26439 6601 26491
rect 6601 26439 6653 26491
rect 6653 26439 6655 26491
rect 6599 26437 6655 26439
rect 6599 26273 6655 26275
rect 6599 26221 6601 26273
rect 6601 26221 6653 26273
rect 6653 26221 6655 26273
rect 6599 26219 6655 26221
rect 6599 26055 6655 26057
rect 6599 26003 6601 26055
rect 6601 26003 6653 26055
rect 6653 26003 6655 26055
rect 6599 26001 6655 26003
rect 6599 25837 6655 25839
rect 6599 25785 6601 25837
rect 6601 25785 6653 25837
rect 6653 25785 6655 25837
rect 6599 25783 6655 25785
rect 1815 24773 1871 24775
rect 1815 24721 1817 24773
rect 1817 24721 1869 24773
rect 1869 24721 1871 24773
rect 1815 24719 1871 24721
rect 1815 24556 1871 24558
rect 1815 24504 1817 24556
rect 1817 24504 1869 24556
rect 1869 24504 1871 24556
rect 1815 24502 1871 24504
rect 1815 24338 1871 24340
rect 1815 24286 1817 24338
rect 1817 24286 1869 24338
rect 1869 24286 1871 24338
rect 1815 24284 1871 24286
rect 1815 24121 1871 24123
rect 1815 24069 1817 24121
rect 1817 24069 1869 24121
rect 1869 24069 1871 24121
rect 1815 24067 1871 24069
rect 1815 23903 1871 23905
rect 1815 23851 1817 23903
rect 1817 23851 1869 23903
rect 1869 23851 1871 23903
rect 1815 23849 1871 23851
rect 1815 23685 1871 23687
rect 1815 23633 1817 23685
rect 1817 23633 1869 23685
rect 1869 23633 1871 23685
rect 1815 23631 1871 23633
rect 1815 23467 1871 23469
rect 1815 23415 1817 23467
rect 1817 23415 1869 23467
rect 1869 23415 1871 23467
rect 1815 23413 1871 23415
rect 1815 23250 1871 23252
rect 1815 23198 1817 23250
rect 1817 23198 1869 23250
rect 1869 23198 1871 23250
rect 1815 23196 1871 23198
rect 1815 23032 1871 23034
rect 1815 22980 1817 23032
rect 1817 22980 1869 23032
rect 1869 22980 1871 23032
rect 1815 22978 1871 22980
rect 1815 22815 1871 22817
rect 1815 22763 1817 22815
rect 1817 22763 1869 22815
rect 1869 22763 1871 22815
rect 1815 22761 1871 22763
rect 2267 24773 2323 24775
rect 2267 24721 2269 24773
rect 2269 24721 2321 24773
rect 2321 24721 2323 24773
rect 2267 24719 2323 24721
rect 2550 24773 2606 24775
rect 2550 24721 2552 24773
rect 2552 24721 2604 24773
rect 2604 24721 2606 24773
rect 2550 24719 2606 24721
rect 2833 24773 2889 24775
rect 2833 24721 2835 24773
rect 2835 24721 2887 24773
rect 2887 24721 2889 24773
rect 2833 24719 2889 24721
rect 2267 24556 2323 24558
rect 2267 24504 2269 24556
rect 2269 24504 2321 24556
rect 2321 24504 2323 24556
rect 2267 24502 2323 24504
rect 2550 24556 2606 24558
rect 2550 24504 2552 24556
rect 2552 24504 2604 24556
rect 2604 24504 2606 24556
rect 2550 24502 2606 24504
rect 2833 24556 2889 24558
rect 2833 24504 2835 24556
rect 2835 24504 2887 24556
rect 2887 24504 2889 24556
rect 2833 24502 2889 24504
rect 2267 24338 2323 24340
rect 2267 24286 2269 24338
rect 2269 24286 2321 24338
rect 2321 24286 2323 24338
rect 2267 24284 2323 24286
rect 2550 24338 2606 24340
rect 2550 24286 2552 24338
rect 2552 24286 2604 24338
rect 2604 24286 2606 24338
rect 2550 24284 2606 24286
rect 2833 24338 2889 24340
rect 2833 24286 2835 24338
rect 2835 24286 2887 24338
rect 2887 24286 2889 24338
rect 2833 24284 2889 24286
rect 2267 24121 2323 24123
rect 2267 24069 2269 24121
rect 2269 24069 2321 24121
rect 2321 24069 2323 24121
rect 2267 24067 2323 24069
rect 2550 24121 2606 24123
rect 2550 24069 2552 24121
rect 2552 24069 2604 24121
rect 2604 24069 2606 24121
rect 2550 24067 2606 24069
rect 2833 24121 2889 24123
rect 2833 24069 2835 24121
rect 2835 24069 2887 24121
rect 2887 24069 2889 24121
rect 2833 24067 2889 24069
rect 2267 23903 2323 23905
rect 2267 23851 2269 23903
rect 2269 23851 2321 23903
rect 2321 23851 2323 23903
rect 2267 23849 2323 23851
rect 2550 23903 2606 23905
rect 2550 23851 2552 23903
rect 2552 23851 2604 23903
rect 2604 23851 2606 23903
rect 2550 23849 2606 23851
rect 2833 23903 2889 23905
rect 2833 23851 2835 23903
rect 2835 23851 2887 23903
rect 2887 23851 2889 23903
rect 2833 23849 2889 23851
rect 2267 23685 2323 23687
rect 2267 23633 2269 23685
rect 2269 23633 2321 23685
rect 2321 23633 2323 23685
rect 2267 23631 2323 23633
rect 2550 23685 2606 23687
rect 2550 23633 2552 23685
rect 2552 23633 2604 23685
rect 2604 23633 2606 23685
rect 2550 23631 2606 23633
rect 2833 23685 2889 23687
rect 2833 23633 2835 23685
rect 2835 23633 2887 23685
rect 2887 23633 2889 23685
rect 2833 23631 2889 23633
rect 2267 23467 2323 23469
rect 2267 23415 2269 23467
rect 2269 23415 2321 23467
rect 2321 23415 2323 23467
rect 2267 23413 2323 23415
rect 2550 23467 2606 23469
rect 2550 23415 2552 23467
rect 2552 23415 2604 23467
rect 2604 23415 2606 23467
rect 2550 23413 2606 23415
rect 2833 23467 2889 23469
rect 2833 23415 2835 23467
rect 2835 23415 2887 23467
rect 2887 23415 2889 23467
rect 2833 23413 2889 23415
rect 2267 23250 2323 23252
rect 2267 23198 2269 23250
rect 2269 23198 2321 23250
rect 2321 23198 2323 23250
rect 2267 23196 2323 23198
rect 2550 23250 2606 23252
rect 2550 23198 2552 23250
rect 2552 23198 2604 23250
rect 2604 23198 2606 23250
rect 2550 23196 2606 23198
rect 2833 23250 2889 23252
rect 2833 23198 2835 23250
rect 2835 23198 2887 23250
rect 2887 23198 2889 23250
rect 2833 23196 2889 23198
rect 2267 23032 2323 23034
rect 2267 22980 2269 23032
rect 2269 22980 2321 23032
rect 2321 22980 2323 23032
rect 2267 22978 2323 22980
rect 2550 23032 2606 23034
rect 2550 22980 2552 23032
rect 2552 22980 2604 23032
rect 2604 22980 2606 23032
rect 2550 22978 2606 22980
rect 2833 23032 2889 23034
rect 2833 22980 2835 23032
rect 2835 22980 2887 23032
rect 2887 22980 2889 23032
rect 2833 22978 2889 22980
rect 2267 22815 2323 22817
rect 2267 22763 2269 22815
rect 2269 22763 2321 22815
rect 2321 22763 2323 22815
rect 2267 22761 2323 22763
rect 2550 22815 2606 22817
rect 2550 22763 2552 22815
rect 2552 22763 2604 22815
rect 2604 22763 2606 22815
rect 2550 22761 2606 22763
rect 2833 22815 2889 22817
rect 2833 22763 2835 22815
rect 2835 22763 2887 22815
rect 2887 22763 2889 22815
rect 2833 22761 2889 22763
rect 3285 24773 3341 24775
rect 3285 24721 3287 24773
rect 3287 24721 3339 24773
rect 3339 24721 3341 24773
rect 3285 24719 3341 24721
rect 3285 24556 3341 24558
rect 3285 24504 3287 24556
rect 3287 24504 3339 24556
rect 3339 24504 3341 24556
rect 3285 24502 3341 24504
rect 3285 24338 3341 24340
rect 3285 24286 3287 24338
rect 3287 24286 3339 24338
rect 3339 24286 3341 24338
rect 3285 24284 3341 24286
rect 3285 24121 3341 24123
rect 3285 24069 3287 24121
rect 3287 24069 3339 24121
rect 3339 24069 3341 24121
rect 3285 24067 3341 24069
rect 3285 23903 3341 23905
rect 3285 23851 3287 23903
rect 3287 23851 3339 23903
rect 3339 23851 3341 23903
rect 3285 23849 3341 23851
rect 3285 23685 3341 23687
rect 3285 23633 3287 23685
rect 3287 23633 3339 23685
rect 3339 23633 3341 23685
rect 3285 23631 3341 23633
rect 3285 23467 3341 23469
rect 3285 23415 3287 23467
rect 3287 23415 3339 23467
rect 3339 23415 3341 23467
rect 3285 23413 3341 23415
rect 3285 23250 3341 23252
rect 3285 23198 3287 23250
rect 3287 23198 3339 23250
rect 3339 23198 3341 23250
rect 3285 23196 3341 23198
rect 3285 23032 3341 23034
rect 3285 22980 3287 23032
rect 3287 22980 3339 23032
rect 3339 22980 3341 23032
rect 3285 22978 3341 22980
rect 3285 22815 3341 22817
rect 3285 22763 3287 22815
rect 3287 22763 3339 22815
rect 3339 22763 3341 22815
rect 3285 22761 3341 22763
rect 3607 24773 3663 24775
rect 3607 24721 3609 24773
rect 3609 24721 3661 24773
rect 3661 24721 3663 24773
rect 3607 24719 3663 24721
rect 3607 24556 3663 24558
rect 3607 24504 3609 24556
rect 3609 24504 3661 24556
rect 3661 24504 3663 24556
rect 3607 24502 3663 24504
rect 3607 24338 3663 24340
rect 3607 24286 3609 24338
rect 3609 24286 3661 24338
rect 3661 24286 3663 24338
rect 3607 24284 3663 24286
rect 3607 24121 3663 24123
rect 3607 24069 3609 24121
rect 3609 24069 3661 24121
rect 3661 24069 3663 24121
rect 3607 24067 3663 24069
rect 3607 23903 3663 23905
rect 3607 23851 3609 23903
rect 3609 23851 3661 23903
rect 3661 23851 3663 23903
rect 3607 23849 3663 23851
rect 3607 23685 3663 23687
rect 3607 23633 3609 23685
rect 3609 23633 3661 23685
rect 3661 23633 3663 23685
rect 3607 23631 3663 23633
rect 3607 23467 3663 23469
rect 3607 23415 3609 23467
rect 3609 23415 3661 23467
rect 3661 23415 3663 23467
rect 3607 23413 3663 23415
rect 3607 23250 3663 23252
rect 3607 23198 3609 23250
rect 3609 23198 3661 23250
rect 3661 23198 3663 23250
rect 3607 23196 3663 23198
rect 3607 23032 3663 23034
rect 3607 22980 3609 23032
rect 3609 22980 3661 23032
rect 3661 22980 3663 23032
rect 3607 22978 3663 22980
rect 3607 22815 3663 22817
rect 3607 22763 3609 22815
rect 3609 22763 3661 22815
rect 3661 22763 3663 22815
rect 3607 22761 3663 22763
rect 4059 24773 4115 24775
rect 4059 24721 4061 24773
rect 4061 24721 4113 24773
rect 4113 24721 4115 24773
rect 4059 24719 4115 24721
rect 4342 24773 4398 24775
rect 4342 24721 4344 24773
rect 4344 24721 4396 24773
rect 4396 24721 4398 24773
rect 4342 24719 4398 24721
rect 4625 24773 4681 24775
rect 4625 24721 4627 24773
rect 4627 24721 4679 24773
rect 4679 24721 4681 24773
rect 4625 24719 4681 24721
rect 4059 24556 4115 24558
rect 4059 24504 4061 24556
rect 4061 24504 4113 24556
rect 4113 24504 4115 24556
rect 4059 24502 4115 24504
rect 4342 24556 4398 24558
rect 4342 24504 4344 24556
rect 4344 24504 4396 24556
rect 4396 24504 4398 24556
rect 4342 24502 4398 24504
rect 4625 24556 4681 24558
rect 4625 24504 4627 24556
rect 4627 24504 4679 24556
rect 4679 24504 4681 24556
rect 4625 24502 4681 24504
rect 4059 24338 4115 24340
rect 4059 24286 4061 24338
rect 4061 24286 4113 24338
rect 4113 24286 4115 24338
rect 4059 24284 4115 24286
rect 4342 24338 4398 24340
rect 4342 24286 4344 24338
rect 4344 24286 4396 24338
rect 4396 24286 4398 24338
rect 4342 24284 4398 24286
rect 4625 24338 4681 24340
rect 4625 24286 4627 24338
rect 4627 24286 4679 24338
rect 4679 24286 4681 24338
rect 4625 24284 4681 24286
rect 4059 24121 4115 24123
rect 4059 24069 4061 24121
rect 4061 24069 4113 24121
rect 4113 24069 4115 24121
rect 4059 24067 4115 24069
rect 4342 24121 4398 24123
rect 4342 24069 4344 24121
rect 4344 24069 4396 24121
rect 4396 24069 4398 24121
rect 4342 24067 4398 24069
rect 4625 24121 4681 24123
rect 4625 24069 4627 24121
rect 4627 24069 4679 24121
rect 4679 24069 4681 24121
rect 4625 24067 4681 24069
rect 4059 23903 4115 23905
rect 4059 23851 4061 23903
rect 4061 23851 4113 23903
rect 4113 23851 4115 23903
rect 4059 23849 4115 23851
rect 4342 23903 4398 23905
rect 4342 23851 4344 23903
rect 4344 23851 4396 23903
rect 4396 23851 4398 23903
rect 4342 23849 4398 23851
rect 4625 23903 4681 23905
rect 4625 23851 4627 23903
rect 4627 23851 4679 23903
rect 4679 23851 4681 23903
rect 4625 23849 4681 23851
rect 4059 23685 4115 23687
rect 4059 23633 4061 23685
rect 4061 23633 4113 23685
rect 4113 23633 4115 23685
rect 4059 23631 4115 23633
rect 4342 23685 4398 23687
rect 4342 23633 4344 23685
rect 4344 23633 4396 23685
rect 4396 23633 4398 23685
rect 4342 23631 4398 23633
rect 4625 23685 4681 23687
rect 4625 23633 4627 23685
rect 4627 23633 4679 23685
rect 4679 23633 4681 23685
rect 4625 23631 4681 23633
rect 4059 23467 4115 23469
rect 4059 23415 4061 23467
rect 4061 23415 4113 23467
rect 4113 23415 4115 23467
rect 4059 23413 4115 23415
rect 4342 23467 4398 23469
rect 4342 23415 4344 23467
rect 4344 23415 4396 23467
rect 4396 23415 4398 23467
rect 4342 23413 4398 23415
rect 4625 23467 4681 23469
rect 4625 23415 4627 23467
rect 4627 23415 4679 23467
rect 4679 23415 4681 23467
rect 4625 23413 4681 23415
rect 4059 23250 4115 23252
rect 4059 23198 4061 23250
rect 4061 23198 4113 23250
rect 4113 23198 4115 23250
rect 4059 23196 4115 23198
rect 4342 23250 4398 23252
rect 4342 23198 4344 23250
rect 4344 23198 4396 23250
rect 4396 23198 4398 23250
rect 4342 23196 4398 23198
rect 4625 23250 4681 23252
rect 4625 23198 4627 23250
rect 4627 23198 4679 23250
rect 4679 23198 4681 23250
rect 4625 23196 4681 23198
rect 4059 23032 4115 23034
rect 4059 22980 4061 23032
rect 4061 22980 4113 23032
rect 4113 22980 4115 23032
rect 4059 22978 4115 22980
rect 4342 23032 4398 23034
rect 4342 22980 4344 23032
rect 4344 22980 4396 23032
rect 4396 22980 4398 23032
rect 4342 22978 4398 22980
rect 4625 23032 4681 23034
rect 4625 22980 4627 23032
rect 4627 22980 4679 23032
rect 4679 22980 4681 23032
rect 4625 22978 4681 22980
rect 4059 22815 4115 22817
rect 4059 22763 4061 22815
rect 4061 22763 4113 22815
rect 4113 22763 4115 22815
rect 4059 22761 4115 22763
rect 4342 22815 4398 22817
rect 4342 22763 4344 22815
rect 4344 22763 4396 22815
rect 4396 22763 4398 22815
rect 4342 22761 4398 22763
rect 4625 22815 4681 22817
rect 4625 22763 4627 22815
rect 4627 22763 4679 22815
rect 4679 22763 4681 22815
rect 4625 22761 4681 22763
rect 5077 24773 5133 24775
rect 5077 24721 5079 24773
rect 5079 24721 5131 24773
rect 5131 24721 5133 24773
rect 5077 24719 5133 24721
rect 5077 24556 5133 24558
rect 5077 24504 5079 24556
rect 5079 24504 5131 24556
rect 5131 24504 5133 24556
rect 5077 24502 5133 24504
rect 5077 24338 5133 24340
rect 5077 24286 5079 24338
rect 5079 24286 5131 24338
rect 5131 24286 5133 24338
rect 5077 24284 5133 24286
rect 5077 24121 5133 24123
rect 5077 24069 5079 24121
rect 5079 24069 5131 24121
rect 5131 24069 5133 24121
rect 5077 24067 5133 24069
rect 5077 23903 5133 23905
rect 5077 23851 5079 23903
rect 5079 23851 5131 23903
rect 5131 23851 5133 23903
rect 5077 23849 5133 23851
rect 5077 23685 5133 23687
rect 5077 23633 5079 23685
rect 5079 23633 5131 23685
rect 5131 23633 5133 23685
rect 5077 23631 5133 23633
rect 5077 23467 5133 23469
rect 5077 23415 5079 23467
rect 5079 23415 5131 23467
rect 5131 23415 5133 23467
rect 5077 23413 5133 23415
rect 5077 23250 5133 23252
rect 5077 23198 5079 23250
rect 5079 23198 5131 23250
rect 5131 23198 5133 23250
rect 5077 23196 5133 23198
rect 5077 23032 5133 23034
rect 5077 22980 5079 23032
rect 5079 22980 5131 23032
rect 5131 22980 5133 23032
rect 5077 22978 5133 22980
rect 5077 22815 5133 22817
rect 5077 22763 5079 22815
rect 5079 22763 5131 22815
rect 5131 22763 5133 22815
rect 5077 22761 5133 22763
rect 2267 20364 2323 20366
rect 2267 20312 2269 20364
rect 2269 20312 2321 20364
rect 2321 20312 2323 20364
rect 2267 20310 2323 20312
rect 2550 20364 2606 20366
rect 2550 20312 2552 20364
rect 2552 20312 2604 20364
rect 2604 20312 2606 20364
rect 2550 20310 2606 20312
rect 2833 20364 2889 20366
rect 2833 20312 2835 20364
rect 2835 20312 2887 20364
rect 2887 20312 2889 20364
rect 2833 20310 2889 20312
rect 2267 20146 2323 20148
rect 2267 20094 2269 20146
rect 2269 20094 2321 20146
rect 2321 20094 2323 20146
rect 2267 20092 2323 20094
rect 2550 20146 2606 20148
rect 2550 20094 2552 20146
rect 2552 20094 2604 20146
rect 2604 20094 2606 20146
rect 2550 20092 2606 20094
rect 2833 20146 2889 20148
rect 2833 20094 2835 20146
rect 2835 20094 2887 20146
rect 2887 20094 2889 20146
rect 2833 20092 2889 20094
rect 2267 19929 2323 19930
rect 2267 19877 2269 19929
rect 2269 19877 2321 19929
rect 2321 19877 2323 19929
rect 2267 19874 2323 19877
rect 2550 19929 2606 19930
rect 2550 19877 2552 19929
rect 2552 19877 2604 19929
rect 2604 19877 2606 19929
rect 2550 19874 2606 19877
rect 2833 19929 2889 19930
rect 2833 19877 2835 19929
rect 2835 19877 2887 19929
rect 2887 19877 2889 19929
rect 2833 19874 2889 19877
rect 4059 20364 4115 20366
rect 4059 20312 4061 20364
rect 4061 20312 4113 20364
rect 4113 20312 4115 20364
rect 4059 20310 4115 20312
rect 4342 20364 4398 20366
rect 4342 20312 4344 20364
rect 4344 20312 4396 20364
rect 4396 20312 4398 20364
rect 4342 20310 4398 20312
rect 4625 20364 4681 20366
rect 4625 20312 4627 20364
rect 4627 20312 4679 20364
rect 4679 20312 4681 20364
rect 4625 20310 4681 20312
rect 4059 20146 4115 20148
rect 4059 20094 4061 20146
rect 4061 20094 4113 20146
rect 4113 20094 4115 20146
rect 4059 20092 4115 20094
rect 4342 20146 4398 20148
rect 4342 20094 4344 20146
rect 4344 20094 4396 20146
rect 4396 20094 4398 20146
rect 4342 20092 4398 20094
rect 4625 20146 4681 20148
rect 4625 20094 4627 20146
rect 4627 20094 4679 20146
rect 4679 20094 4681 20146
rect 4625 20092 4681 20094
rect 4059 19929 4115 19930
rect 4059 19877 4061 19929
rect 4061 19877 4113 19929
rect 4113 19877 4115 19929
rect 4059 19874 4115 19877
rect 4342 19929 4398 19930
rect 4342 19877 4344 19929
rect 4344 19877 4396 19929
rect 4396 19877 4398 19929
rect 4342 19874 4398 19877
rect 4625 19929 4681 19930
rect 4625 19877 4627 19929
rect 4627 19877 4679 19929
rect 4679 19877 4681 19929
rect 4625 19874 4681 19877
rect 2267 18405 2323 18408
rect 2267 18353 2269 18405
rect 2269 18353 2321 18405
rect 2321 18353 2323 18405
rect 2267 18352 2323 18353
rect 2550 18405 2606 18408
rect 2550 18353 2552 18405
rect 2552 18353 2604 18405
rect 2604 18353 2606 18405
rect 2550 18352 2606 18353
rect 2833 18405 2889 18408
rect 2833 18353 2835 18405
rect 2835 18353 2887 18405
rect 2887 18353 2889 18405
rect 2833 18352 2889 18353
rect 2267 18188 2323 18190
rect 2267 18136 2269 18188
rect 2269 18136 2321 18188
rect 2321 18136 2323 18188
rect 2267 18134 2323 18136
rect 2550 18188 2606 18190
rect 2550 18136 2552 18188
rect 2552 18136 2604 18188
rect 2604 18136 2606 18188
rect 2550 18134 2606 18136
rect 2833 18188 2889 18190
rect 2833 18136 2835 18188
rect 2835 18136 2887 18188
rect 2887 18136 2889 18188
rect 2833 18134 2889 18136
rect 2267 17970 2323 17972
rect 2267 17918 2269 17970
rect 2269 17918 2321 17970
rect 2321 17918 2323 17970
rect 2267 17916 2323 17918
rect 2550 17970 2606 17972
rect 2550 17918 2552 17970
rect 2552 17918 2604 17970
rect 2604 17918 2606 17970
rect 2550 17916 2606 17918
rect 2833 17970 2889 17972
rect 2833 17918 2835 17970
rect 2835 17918 2887 17970
rect 2887 17918 2889 17970
rect 2833 17916 2889 17918
rect 2267 17698 2323 17754
rect 2550 17698 2606 17754
rect 2833 17698 2889 17754
rect 6092 24802 6148 24804
rect 6092 24750 6094 24802
rect 6094 24750 6146 24802
rect 6146 24750 6148 24802
rect 6092 24748 6148 24750
rect 6092 24585 6148 24587
rect 6092 24533 6094 24585
rect 6094 24533 6146 24585
rect 6146 24533 6148 24585
rect 6092 24531 6148 24533
rect 6092 24367 6148 24369
rect 6092 24315 6094 24367
rect 6094 24315 6146 24367
rect 6146 24315 6148 24367
rect 6092 24313 6148 24315
rect 6092 24150 6148 24152
rect 6092 24098 6094 24150
rect 6094 24098 6146 24150
rect 6146 24098 6148 24150
rect 6092 24096 6148 24098
rect 6092 23932 6148 23934
rect 6092 23880 6094 23932
rect 6094 23880 6146 23932
rect 6146 23880 6148 23932
rect 6092 23878 6148 23880
rect 6092 23714 6148 23716
rect 6092 23662 6094 23714
rect 6094 23662 6146 23714
rect 6146 23662 6148 23714
rect 6092 23660 6148 23662
rect 6092 23496 6148 23498
rect 6092 23444 6094 23496
rect 6094 23444 6146 23496
rect 6146 23444 6148 23496
rect 6092 23442 6148 23444
rect 6092 23279 6148 23281
rect 6092 23227 6094 23279
rect 6094 23227 6146 23279
rect 6146 23227 6148 23279
rect 6092 23225 6148 23227
rect 6606 24811 6662 24813
rect 6606 24759 6608 24811
rect 6608 24759 6660 24811
rect 6660 24759 6662 24811
rect 6606 24757 6662 24759
rect 6606 24593 6662 24595
rect 6606 24541 6608 24593
rect 6608 24541 6660 24593
rect 6660 24541 6662 24593
rect 6606 24539 6662 24541
rect 6606 24376 6662 24378
rect 6606 24324 6608 24376
rect 6608 24324 6660 24376
rect 6660 24324 6662 24376
rect 6606 24322 6662 24324
rect 6606 24158 6662 24160
rect 6606 24106 6608 24158
rect 6608 24106 6660 24158
rect 6660 24106 6662 24158
rect 6606 24104 6662 24106
rect 6606 23940 6662 23942
rect 6606 23888 6608 23940
rect 6608 23888 6660 23940
rect 6660 23888 6662 23940
rect 6606 23886 6662 23888
rect 6606 23722 6662 23724
rect 6606 23670 6608 23722
rect 6608 23670 6660 23722
rect 6660 23670 6662 23722
rect 6606 23668 6662 23670
rect 6606 23505 6662 23507
rect 6606 23453 6608 23505
rect 6608 23453 6660 23505
rect 6660 23453 6662 23505
rect 6606 23451 6662 23453
rect 6606 23287 6662 23289
rect 6606 23235 6608 23287
rect 6608 23235 6660 23287
rect 6660 23235 6662 23287
rect 6606 23233 6662 23235
rect 6092 23061 6148 23063
rect 6092 23009 6094 23061
rect 6094 23009 6146 23061
rect 6146 23009 6148 23061
rect 6092 23007 6148 23009
rect 17826 28392 17882 28394
rect 17826 28340 17828 28392
rect 17828 28340 17880 28392
rect 17880 28340 17882 28392
rect 17826 28338 17882 28340
rect 17826 28174 17882 28176
rect 17826 28122 17828 28174
rect 17828 28122 17880 28174
rect 17880 28122 17882 28174
rect 17826 28120 17882 28122
rect 17826 27956 17882 27958
rect 17826 27904 17828 27956
rect 17828 27904 17880 27956
rect 17880 27904 17882 27956
rect 17826 27902 17882 27904
rect 17826 27738 17882 27740
rect 17826 27686 17828 27738
rect 17828 27686 17880 27738
rect 17880 27686 17882 27738
rect 17826 27684 17882 27686
rect 18550 28392 18606 28394
rect 18550 28340 18552 28392
rect 18552 28340 18604 28392
rect 18604 28340 18606 28392
rect 18550 28338 18606 28340
rect 18550 28174 18606 28176
rect 18550 28122 18552 28174
rect 18552 28122 18604 28174
rect 18604 28122 18606 28174
rect 18550 28120 18606 28122
rect 18550 27956 18606 27958
rect 18550 27904 18552 27956
rect 18552 27904 18604 27956
rect 18604 27904 18606 27956
rect 18550 27902 18606 27904
rect 18550 27738 18606 27740
rect 18550 27686 18552 27738
rect 18552 27686 18604 27738
rect 18604 27686 18606 27738
rect 18550 27684 18606 27686
rect 19460 28392 19516 28394
rect 19460 28340 19462 28392
rect 19462 28340 19514 28392
rect 19514 28340 19516 28392
rect 19460 28338 19516 28340
rect 19460 28174 19516 28176
rect 19460 28122 19462 28174
rect 19462 28122 19514 28174
rect 19514 28122 19516 28174
rect 19460 28120 19516 28122
rect 19460 27956 19516 27958
rect 19460 27904 19462 27956
rect 19462 27904 19514 27956
rect 19514 27904 19516 27956
rect 19460 27902 19516 27904
rect 19460 27738 19516 27740
rect 19460 27686 19462 27738
rect 19462 27686 19514 27738
rect 19514 27686 19516 27738
rect 19460 27684 19516 27686
rect 20183 28392 20239 28394
rect 20183 28340 20185 28392
rect 20185 28340 20237 28392
rect 20237 28340 20239 28392
rect 20183 28338 20239 28340
rect 20183 28174 20239 28176
rect 20183 28122 20185 28174
rect 20185 28122 20237 28174
rect 20237 28122 20239 28174
rect 20183 28120 20239 28122
rect 20183 27956 20239 27958
rect 20183 27904 20185 27956
rect 20185 27904 20237 27956
rect 20237 27904 20239 27956
rect 20183 27902 20239 27904
rect 20183 27738 20239 27740
rect 20183 27686 20185 27738
rect 20185 27686 20237 27738
rect 20237 27686 20239 27738
rect 20183 27684 20239 27686
rect 21093 28392 21149 28394
rect 21093 28340 21095 28392
rect 21095 28340 21147 28392
rect 21147 28340 21149 28392
rect 21093 28338 21149 28340
rect 21093 28174 21149 28176
rect 21093 28122 21095 28174
rect 21095 28122 21147 28174
rect 21147 28122 21149 28174
rect 21093 28120 21149 28122
rect 21093 27956 21149 27958
rect 21093 27904 21095 27956
rect 21095 27904 21147 27956
rect 21147 27904 21149 27956
rect 21093 27902 21149 27904
rect 21093 27738 21149 27740
rect 21093 27686 21095 27738
rect 21095 27686 21147 27738
rect 21147 27686 21149 27738
rect 21093 27684 21149 27686
rect 21817 28392 21873 28394
rect 21817 28340 21819 28392
rect 21819 28340 21871 28392
rect 21871 28340 21873 28392
rect 21817 28338 21873 28340
rect 21817 28174 21873 28176
rect 21817 28122 21819 28174
rect 21819 28122 21871 28174
rect 21871 28122 21873 28174
rect 21817 28120 21873 28122
rect 21817 27956 21873 27958
rect 21817 27904 21819 27956
rect 21819 27904 21871 27956
rect 21871 27904 21873 27956
rect 21817 27902 21873 27904
rect 21817 27738 21873 27740
rect 21817 27686 21819 27738
rect 21819 27686 21871 27738
rect 21871 27686 21873 27738
rect 21817 27684 21873 27686
rect 22727 28392 22783 28394
rect 22727 28340 22729 28392
rect 22729 28340 22781 28392
rect 22781 28340 22783 28392
rect 22727 28338 22783 28340
rect 22727 28174 22783 28176
rect 22727 28122 22729 28174
rect 22729 28122 22781 28174
rect 22781 28122 22783 28174
rect 22727 28120 22783 28122
rect 22727 27956 22783 27958
rect 22727 27904 22729 27956
rect 22729 27904 22781 27956
rect 22781 27904 22783 27956
rect 22727 27902 22783 27904
rect 22727 27738 22783 27740
rect 22727 27686 22729 27738
rect 22729 27686 22781 27738
rect 22781 27686 22783 27738
rect 22727 27684 22783 27686
rect 28627 29970 28683 30026
rect 28838 29970 28894 30026
rect 29050 29970 29106 30026
rect 29261 29970 29317 30026
rect 28627 29752 28683 29808
rect 28838 29752 28894 29808
rect 29050 29752 29106 29808
rect 29261 29752 29317 29808
rect 28627 29534 28683 29590
rect 28838 29534 28894 29590
rect 29050 29534 29106 29590
rect 29261 29534 29317 29590
rect 28627 29316 28683 29372
rect 28838 29316 28894 29372
rect 29050 29316 29106 29372
rect 29261 29316 29317 29372
rect 24444 28943 24500 28999
rect 24444 28725 24500 28781
rect 23785 28401 23841 28403
rect 23785 28349 23787 28401
rect 23787 28349 23839 28401
rect 23839 28349 23841 28401
rect 23785 28347 23841 28349
rect 23785 28183 23841 28185
rect 23785 28131 23787 28183
rect 23787 28131 23839 28183
rect 23839 28131 23841 28183
rect 23785 28129 23841 28131
rect 23785 27965 23841 27967
rect 23785 27913 23787 27965
rect 23787 27913 23839 27965
rect 23839 27913 23841 27965
rect 23785 27911 23841 27913
rect 24224 28401 24280 28403
rect 24224 28349 24226 28401
rect 24226 28349 24278 28401
rect 24278 28349 24280 28401
rect 24224 28347 24280 28349
rect 24224 28183 24280 28185
rect 24224 28131 24226 28183
rect 24226 28131 24278 28183
rect 24278 28131 24280 28183
rect 24224 28129 24280 28131
rect 24224 27965 24280 27967
rect 24224 27913 24226 27965
rect 24226 27913 24278 27965
rect 24278 27913 24280 27965
rect 24224 27911 24280 27913
rect 25608 28344 25664 28346
rect 25608 28292 25610 28344
rect 25610 28292 25662 28344
rect 25662 28292 25664 28344
rect 25608 28290 25664 28292
rect 25608 28126 25664 28128
rect 25608 28074 25610 28126
rect 25610 28074 25662 28126
rect 25662 28074 25664 28126
rect 25608 28072 25664 28074
rect 25608 27908 25664 27910
rect 25608 27856 25610 27908
rect 25610 27856 25662 27908
rect 25662 27856 25664 27908
rect 25608 27854 25664 27856
rect 7563 26514 7619 26516
rect 7563 26462 7565 26514
rect 7565 26462 7617 26514
rect 7617 26462 7619 26514
rect 7563 26460 7619 26462
rect 7770 26514 7826 26516
rect 7770 26462 7772 26514
rect 7772 26462 7824 26514
rect 7824 26462 7826 26514
rect 7770 26460 7826 26462
rect 7563 26296 7619 26298
rect 7563 26244 7565 26296
rect 7565 26244 7617 26296
rect 7617 26244 7619 26296
rect 7563 26242 7619 26244
rect 7770 26296 7826 26298
rect 7770 26244 7772 26296
rect 7772 26244 7824 26296
rect 7824 26244 7826 26296
rect 7770 26242 7826 26244
rect 7563 26078 7619 26080
rect 7563 26026 7565 26078
rect 7565 26026 7617 26078
rect 7617 26026 7619 26078
rect 7563 26024 7619 26026
rect 7770 26078 7826 26080
rect 7770 26026 7772 26078
rect 7772 26026 7824 26078
rect 7824 26026 7826 26078
rect 7770 26024 7826 26026
rect 7563 25860 7619 25862
rect 7563 25808 7565 25860
rect 7565 25808 7617 25860
rect 7617 25808 7619 25860
rect 7563 25806 7619 25808
rect 7770 25860 7826 25862
rect 7770 25808 7772 25860
rect 7772 25808 7824 25860
rect 7824 25808 7826 25860
rect 7770 25806 7826 25808
rect 8290 26491 8346 26493
rect 8290 26439 8292 26491
rect 8292 26439 8344 26491
rect 8344 26439 8346 26491
rect 8290 26437 8346 26439
rect 8290 26273 8346 26275
rect 8290 26221 8292 26273
rect 8292 26221 8344 26273
rect 8344 26221 8346 26273
rect 8290 26219 8346 26221
rect 8290 26055 8346 26057
rect 8290 26003 8292 26055
rect 8292 26003 8344 26055
rect 8344 26003 8346 26055
rect 8290 26001 8346 26003
rect 8290 25837 8346 25839
rect 8290 25785 8292 25837
rect 8292 25785 8344 25837
rect 8344 25785 8346 25837
rect 8290 25783 8346 25785
rect 6092 22844 6148 22846
rect 6092 22792 6094 22844
rect 6094 22792 6146 22844
rect 6146 22792 6148 22844
rect 6092 22790 6148 22792
rect 6595 21511 6651 21567
rect 6595 21293 6651 21349
rect 7085 21987 7141 22043
rect 7085 21769 7141 21825
rect 7783 24802 7839 24804
rect 7783 24750 7785 24802
rect 7785 24750 7837 24802
rect 7837 24750 7839 24802
rect 7783 24748 7839 24750
rect 7783 24585 7839 24587
rect 7783 24533 7785 24585
rect 7785 24533 7837 24585
rect 7837 24533 7839 24585
rect 7783 24531 7839 24533
rect 7783 24367 7839 24369
rect 7783 24315 7785 24367
rect 7785 24315 7837 24367
rect 7837 24315 7839 24367
rect 7783 24313 7839 24315
rect 7783 24150 7839 24152
rect 7783 24098 7785 24150
rect 7785 24098 7837 24150
rect 7837 24098 7839 24150
rect 7783 24096 7839 24098
rect 7783 23932 7839 23934
rect 7783 23880 7785 23932
rect 7785 23880 7837 23932
rect 7837 23880 7839 23932
rect 7783 23878 7839 23880
rect 7783 23714 7839 23716
rect 7783 23662 7785 23714
rect 7785 23662 7837 23714
rect 7837 23662 7839 23714
rect 7783 23660 7839 23662
rect 7783 23496 7839 23498
rect 7783 23444 7785 23496
rect 7785 23444 7837 23496
rect 7837 23444 7839 23496
rect 7783 23442 7839 23444
rect 7783 23279 7839 23281
rect 7783 23227 7785 23279
rect 7785 23227 7837 23279
rect 7837 23227 7839 23279
rect 7783 23225 7839 23227
rect 8297 24811 8353 24813
rect 8297 24759 8299 24811
rect 8299 24759 8351 24811
rect 8351 24759 8353 24811
rect 8297 24757 8353 24759
rect 8297 24593 8353 24595
rect 8297 24541 8299 24593
rect 8299 24541 8351 24593
rect 8351 24541 8353 24593
rect 8297 24539 8353 24541
rect 8297 24376 8353 24378
rect 8297 24324 8299 24376
rect 8299 24324 8351 24376
rect 8351 24324 8353 24376
rect 8297 24322 8353 24324
rect 8297 24158 8353 24160
rect 8297 24106 8299 24158
rect 8299 24106 8351 24158
rect 8351 24106 8353 24158
rect 8297 24104 8353 24106
rect 8297 23940 8353 23942
rect 8297 23888 8299 23940
rect 8299 23888 8351 23940
rect 8351 23888 8353 23940
rect 8297 23886 8353 23888
rect 8297 23722 8353 23724
rect 8297 23670 8299 23722
rect 8299 23670 8351 23722
rect 8351 23670 8353 23722
rect 8297 23668 8353 23670
rect 8297 23505 8353 23507
rect 8297 23453 8299 23505
rect 8299 23453 8351 23505
rect 8351 23453 8353 23505
rect 8297 23451 8353 23453
rect 8297 23287 8353 23289
rect 8297 23235 8299 23287
rect 8299 23235 8351 23287
rect 8351 23235 8353 23287
rect 8297 23233 8353 23235
rect 7783 23061 7839 23063
rect 7783 23009 7785 23061
rect 7785 23009 7837 23061
rect 7837 23009 7839 23061
rect 7783 23007 7839 23009
rect 7783 22844 7839 22846
rect 7783 22792 7785 22844
rect 7785 22792 7837 22844
rect 7837 22792 7839 22844
rect 7783 22790 7839 22792
rect 8286 21511 8342 21567
rect 8286 21293 8342 21349
rect 9033 27353 9089 27355
rect 9033 27301 9035 27353
rect 9035 27301 9087 27353
rect 9087 27301 9089 27353
rect 9033 27299 9089 27301
rect 9033 27135 9089 27137
rect 9033 27083 9035 27135
rect 9035 27083 9087 27135
rect 9087 27083 9089 27135
rect 9033 27081 9089 27083
rect 9033 26917 9089 26919
rect 9033 26865 9035 26917
rect 9035 26865 9087 26917
rect 9087 26865 9089 26917
rect 9033 26863 9089 26865
rect 9481 27353 9537 27355
rect 9481 27301 9483 27353
rect 9483 27301 9535 27353
rect 9535 27301 9537 27353
rect 9481 27299 9537 27301
rect 9481 27135 9537 27137
rect 9481 27083 9483 27135
rect 9483 27083 9535 27135
rect 9535 27083 9537 27135
rect 9481 27081 9537 27083
rect 9481 26917 9537 26919
rect 9481 26865 9483 26917
rect 9483 26865 9535 26917
rect 9535 26865 9537 26917
rect 9481 26863 9537 26865
rect 9929 27353 9985 27355
rect 9929 27301 9931 27353
rect 9931 27301 9983 27353
rect 9983 27301 9985 27353
rect 9929 27299 9985 27301
rect 9929 27135 9985 27137
rect 9929 27083 9931 27135
rect 9931 27083 9983 27135
rect 9983 27083 9985 27135
rect 9929 27081 9985 27083
rect 9929 26917 9985 26919
rect 9929 26865 9931 26917
rect 9931 26865 9983 26917
rect 9983 26865 9985 26917
rect 9929 26863 9985 26865
rect 10377 27353 10433 27355
rect 10377 27301 10379 27353
rect 10379 27301 10431 27353
rect 10431 27301 10433 27353
rect 10377 27299 10433 27301
rect 10377 27135 10433 27137
rect 10377 27083 10379 27135
rect 10379 27083 10431 27135
rect 10431 27083 10433 27135
rect 10377 27081 10433 27083
rect 10377 26917 10433 26919
rect 10377 26865 10379 26917
rect 10379 26865 10431 26917
rect 10431 26865 10433 26917
rect 10377 26863 10433 26865
rect 10825 27353 10881 27355
rect 10825 27301 10827 27353
rect 10827 27301 10879 27353
rect 10879 27301 10881 27353
rect 10825 27299 10881 27301
rect 10825 27135 10881 27137
rect 10825 27083 10827 27135
rect 10827 27083 10879 27135
rect 10879 27083 10881 27135
rect 10825 27081 10881 27083
rect 10825 26917 10881 26919
rect 10825 26865 10827 26917
rect 10827 26865 10879 26917
rect 10879 26865 10881 26917
rect 10825 26863 10881 26865
rect 11273 27353 11329 27355
rect 11273 27301 11275 27353
rect 11275 27301 11327 27353
rect 11327 27301 11329 27353
rect 11273 27299 11329 27301
rect 11273 27135 11329 27137
rect 11273 27083 11275 27135
rect 11275 27083 11327 27135
rect 11327 27083 11329 27135
rect 11273 27081 11329 27083
rect 11273 26917 11329 26919
rect 11273 26865 11275 26917
rect 11275 26865 11327 26917
rect 11327 26865 11329 26917
rect 11273 26863 11329 26865
rect 11721 27353 11777 27355
rect 11721 27301 11723 27353
rect 11723 27301 11775 27353
rect 11775 27301 11777 27353
rect 11721 27299 11777 27301
rect 11721 27135 11777 27137
rect 11721 27083 11723 27135
rect 11723 27083 11775 27135
rect 11775 27083 11777 27135
rect 11721 27081 11777 27083
rect 11721 26917 11777 26919
rect 11721 26865 11723 26917
rect 11723 26865 11775 26917
rect 11775 26865 11777 26917
rect 11721 26863 11777 26865
rect 12169 27353 12225 27355
rect 12169 27301 12171 27353
rect 12171 27301 12223 27353
rect 12223 27301 12225 27353
rect 12169 27299 12225 27301
rect 12169 27135 12225 27137
rect 12169 27083 12171 27135
rect 12171 27083 12223 27135
rect 12223 27083 12225 27135
rect 12169 27081 12225 27083
rect 12169 26917 12225 26919
rect 12169 26865 12171 26917
rect 12171 26865 12223 26917
rect 12223 26865 12225 26917
rect 12169 26863 12225 26865
rect 12617 27353 12673 27355
rect 12617 27301 12619 27353
rect 12619 27301 12671 27353
rect 12671 27301 12673 27353
rect 12617 27299 12673 27301
rect 12617 27135 12673 27137
rect 12617 27083 12619 27135
rect 12619 27083 12671 27135
rect 12671 27083 12673 27135
rect 12617 27081 12673 27083
rect 12617 26917 12673 26919
rect 12617 26865 12619 26917
rect 12619 26865 12671 26917
rect 12671 26865 12673 26917
rect 12617 26863 12673 26865
rect 13024 27378 13080 27380
rect 13024 27326 13026 27378
rect 13026 27326 13078 27378
rect 13078 27326 13080 27378
rect 13024 27324 13080 27326
rect 13024 27160 13080 27162
rect 13024 27108 13026 27160
rect 13026 27108 13078 27160
rect 13078 27108 13080 27160
rect 13024 27106 13080 27108
rect 13024 26888 13080 26944
rect 13300 27378 13356 27380
rect 13300 27326 13302 27378
rect 13302 27326 13354 27378
rect 13354 27326 13356 27378
rect 13300 27324 13356 27326
rect 15513 27392 15569 27394
rect 15513 27340 15515 27392
rect 15515 27340 15567 27392
rect 15567 27340 15569 27392
rect 15513 27338 15569 27340
rect 13300 27160 13356 27162
rect 13300 27108 13302 27160
rect 13302 27108 13354 27160
rect 13354 27108 13356 27160
rect 13300 27106 13356 27108
rect 14384 27210 14440 27212
rect 14384 27158 14386 27210
rect 14386 27158 14438 27210
rect 14438 27158 14440 27210
rect 14384 27156 14440 27158
rect 14596 27210 14652 27212
rect 14596 27158 14598 27210
rect 14598 27158 14650 27210
rect 14650 27158 14652 27210
rect 14596 27156 14652 27158
rect 15513 27174 15569 27176
rect 15513 27122 15515 27174
rect 15515 27122 15567 27174
rect 15567 27122 15569 27174
rect 15513 27120 15569 27122
rect 13300 26888 13356 26944
rect 15513 26902 15569 26958
rect 13251 26514 13307 26516
rect 13251 26462 13253 26514
rect 13253 26462 13305 26514
rect 13305 26462 13307 26514
rect 13251 26460 13307 26462
rect 13458 26514 13514 26516
rect 13458 26462 13460 26514
rect 13460 26462 13512 26514
rect 13512 26462 13514 26514
rect 13458 26460 13514 26462
rect 13251 26296 13307 26298
rect 13251 26244 13253 26296
rect 13253 26244 13305 26296
rect 13305 26244 13307 26296
rect 13251 26242 13307 26244
rect 13458 26296 13514 26298
rect 13458 26244 13460 26296
rect 13460 26244 13512 26296
rect 13512 26244 13514 26296
rect 13458 26242 13514 26244
rect 13251 26078 13307 26080
rect 13251 26026 13253 26078
rect 13253 26026 13305 26078
rect 13305 26026 13307 26078
rect 13251 26024 13307 26026
rect 13458 26078 13514 26080
rect 13458 26026 13460 26078
rect 13460 26026 13512 26078
rect 13512 26026 13514 26078
rect 13458 26024 13514 26026
rect 13251 25860 13307 25862
rect 13251 25808 13253 25860
rect 13253 25808 13305 25860
rect 13305 25808 13307 25860
rect 13251 25806 13307 25808
rect 13458 25860 13514 25862
rect 13458 25808 13460 25860
rect 13460 25808 13512 25860
rect 13512 25808 13514 25860
rect 13458 25806 13514 25808
rect 13978 26491 14034 26493
rect 13978 26439 13980 26491
rect 13980 26439 14032 26491
rect 14032 26439 14034 26491
rect 13978 26437 14034 26439
rect 13978 26273 14034 26275
rect 13978 26221 13980 26273
rect 13980 26221 14032 26273
rect 14032 26221 14034 26273
rect 13978 26219 14034 26221
rect 13978 26055 14034 26057
rect 13978 26003 13980 26055
rect 13980 26003 14032 26055
rect 14032 26003 14034 26055
rect 13978 26001 14034 26003
rect 13978 25837 14034 25839
rect 13978 25785 13980 25837
rect 13980 25785 14032 25837
rect 14032 25785 14034 25837
rect 13978 25783 14034 25785
rect 9194 24773 9250 24775
rect 9194 24721 9196 24773
rect 9196 24721 9248 24773
rect 9248 24721 9250 24773
rect 9194 24719 9250 24721
rect 9194 24556 9250 24558
rect 9194 24504 9196 24556
rect 9196 24504 9248 24556
rect 9248 24504 9250 24556
rect 9194 24502 9250 24504
rect 9194 24338 9250 24340
rect 9194 24286 9196 24338
rect 9196 24286 9248 24338
rect 9248 24286 9250 24338
rect 9194 24284 9250 24286
rect 9194 24121 9250 24123
rect 9194 24069 9196 24121
rect 9196 24069 9248 24121
rect 9248 24069 9250 24121
rect 9194 24067 9250 24069
rect 9194 23903 9250 23905
rect 9194 23851 9196 23903
rect 9196 23851 9248 23903
rect 9248 23851 9250 23903
rect 9194 23849 9250 23851
rect 9194 23685 9250 23687
rect 9194 23633 9196 23685
rect 9196 23633 9248 23685
rect 9248 23633 9250 23685
rect 9194 23631 9250 23633
rect 9194 23467 9250 23469
rect 9194 23415 9196 23467
rect 9196 23415 9248 23467
rect 9248 23415 9250 23467
rect 9194 23413 9250 23415
rect 9194 23250 9250 23252
rect 9194 23198 9196 23250
rect 9196 23198 9248 23250
rect 9248 23198 9250 23250
rect 9194 23196 9250 23198
rect 9194 23032 9250 23034
rect 9194 22980 9196 23032
rect 9196 22980 9248 23032
rect 9248 22980 9250 23032
rect 9194 22978 9250 22980
rect 9194 22815 9250 22817
rect 9194 22763 9196 22815
rect 9196 22763 9248 22815
rect 9248 22763 9250 22815
rect 9194 22761 9250 22763
rect 9646 24773 9702 24775
rect 9646 24721 9648 24773
rect 9648 24721 9700 24773
rect 9700 24721 9702 24773
rect 9646 24719 9702 24721
rect 9929 24773 9985 24775
rect 9929 24721 9931 24773
rect 9931 24721 9983 24773
rect 9983 24721 9985 24773
rect 9929 24719 9985 24721
rect 10212 24773 10268 24775
rect 10212 24721 10214 24773
rect 10214 24721 10266 24773
rect 10266 24721 10268 24773
rect 10212 24719 10268 24721
rect 9646 24556 9702 24558
rect 9646 24504 9648 24556
rect 9648 24504 9700 24556
rect 9700 24504 9702 24556
rect 9646 24502 9702 24504
rect 9929 24556 9985 24558
rect 9929 24504 9931 24556
rect 9931 24504 9983 24556
rect 9983 24504 9985 24556
rect 9929 24502 9985 24504
rect 10212 24556 10268 24558
rect 10212 24504 10214 24556
rect 10214 24504 10266 24556
rect 10266 24504 10268 24556
rect 10212 24502 10268 24504
rect 9646 24338 9702 24340
rect 9646 24286 9648 24338
rect 9648 24286 9700 24338
rect 9700 24286 9702 24338
rect 9646 24284 9702 24286
rect 9929 24338 9985 24340
rect 9929 24286 9931 24338
rect 9931 24286 9983 24338
rect 9983 24286 9985 24338
rect 9929 24284 9985 24286
rect 10212 24338 10268 24340
rect 10212 24286 10214 24338
rect 10214 24286 10266 24338
rect 10266 24286 10268 24338
rect 10212 24284 10268 24286
rect 9646 24121 9702 24123
rect 9646 24069 9648 24121
rect 9648 24069 9700 24121
rect 9700 24069 9702 24121
rect 9646 24067 9702 24069
rect 9929 24121 9985 24123
rect 9929 24069 9931 24121
rect 9931 24069 9983 24121
rect 9983 24069 9985 24121
rect 9929 24067 9985 24069
rect 10212 24121 10268 24123
rect 10212 24069 10214 24121
rect 10214 24069 10266 24121
rect 10266 24069 10268 24121
rect 10212 24067 10268 24069
rect 9646 23903 9702 23905
rect 9646 23851 9648 23903
rect 9648 23851 9700 23903
rect 9700 23851 9702 23903
rect 9646 23849 9702 23851
rect 9929 23903 9985 23905
rect 9929 23851 9931 23903
rect 9931 23851 9983 23903
rect 9983 23851 9985 23903
rect 9929 23849 9985 23851
rect 10212 23903 10268 23905
rect 10212 23851 10214 23903
rect 10214 23851 10266 23903
rect 10266 23851 10268 23903
rect 10212 23849 10268 23851
rect 9646 23685 9702 23687
rect 9646 23633 9648 23685
rect 9648 23633 9700 23685
rect 9700 23633 9702 23685
rect 9646 23631 9702 23633
rect 9929 23685 9985 23687
rect 9929 23633 9931 23685
rect 9931 23633 9983 23685
rect 9983 23633 9985 23685
rect 9929 23631 9985 23633
rect 10212 23685 10268 23687
rect 10212 23633 10214 23685
rect 10214 23633 10266 23685
rect 10266 23633 10268 23685
rect 10212 23631 10268 23633
rect 9646 23467 9702 23469
rect 9646 23415 9648 23467
rect 9648 23415 9700 23467
rect 9700 23415 9702 23467
rect 9646 23413 9702 23415
rect 9929 23467 9985 23469
rect 9929 23415 9931 23467
rect 9931 23415 9983 23467
rect 9983 23415 9985 23467
rect 9929 23413 9985 23415
rect 10212 23467 10268 23469
rect 10212 23415 10214 23467
rect 10214 23415 10266 23467
rect 10266 23415 10268 23467
rect 10212 23413 10268 23415
rect 9646 23250 9702 23252
rect 9646 23198 9648 23250
rect 9648 23198 9700 23250
rect 9700 23198 9702 23250
rect 9646 23196 9702 23198
rect 9929 23250 9985 23252
rect 9929 23198 9931 23250
rect 9931 23198 9983 23250
rect 9983 23198 9985 23250
rect 9929 23196 9985 23198
rect 10212 23250 10268 23252
rect 10212 23198 10214 23250
rect 10214 23198 10266 23250
rect 10266 23198 10268 23250
rect 10212 23196 10268 23198
rect 9646 23032 9702 23034
rect 9646 22980 9648 23032
rect 9648 22980 9700 23032
rect 9700 22980 9702 23032
rect 9646 22978 9702 22980
rect 9929 23032 9985 23034
rect 9929 22980 9931 23032
rect 9931 22980 9983 23032
rect 9983 22980 9985 23032
rect 9929 22978 9985 22980
rect 10212 23032 10268 23034
rect 10212 22980 10214 23032
rect 10214 22980 10266 23032
rect 10266 22980 10268 23032
rect 10212 22978 10268 22980
rect 9646 22815 9702 22817
rect 9646 22763 9648 22815
rect 9648 22763 9700 22815
rect 9700 22763 9702 22815
rect 9646 22761 9702 22763
rect 9929 22815 9985 22817
rect 9929 22763 9931 22815
rect 9931 22763 9983 22815
rect 9983 22763 9985 22815
rect 9929 22761 9985 22763
rect 10212 22815 10268 22817
rect 10212 22763 10214 22815
rect 10214 22763 10266 22815
rect 10266 22763 10268 22815
rect 10212 22761 10268 22763
rect 10664 24773 10720 24775
rect 10664 24721 10666 24773
rect 10666 24721 10718 24773
rect 10718 24721 10720 24773
rect 10664 24719 10720 24721
rect 10664 24556 10720 24558
rect 10664 24504 10666 24556
rect 10666 24504 10718 24556
rect 10718 24504 10720 24556
rect 10664 24502 10720 24504
rect 10664 24338 10720 24340
rect 10664 24286 10666 24338
rect 10666 24286 10718 24338
rect 10718 24286 10720 24338
rect 10664 24284 10720 24286
rect 10664 24121 10720 24123
rect 10664 24069 10666 24121
rect 10666 24069 10718 24121
rect 10718 24069 10720 24121
rect 10664 24067 10720 24069
rect 10664 23903 10720 23905
rect 10664 23851 10666 23903
rect 10666 23851 10718 23903
rect 10718 23851 10720 23903
rect 10664 23849 10720 23851
rect 10664 23685 10720 23687
rect 10664 23633 10666 23685
rect 10666 23633 10718 23685
rect 10718 23633 10720 23685
rect 10664 23631 10720 23633
rect 10664 23467 10720 23469
rect 10664 23415 10666 23467
rect 10666 23415 10718 23467
rect 10718 23415 10720 23467
rect 10664 23413 10720 23415
rect 10664 23250 10720 23252
rect 10664 23198 10666 23250
rect 10666 23198 10718 23250
rect 10718 23198 10720 23250
rect 10664 23196 10720 23198
rect 10664 23032 10720 23034
rect 10664 22980 10666 23032
rect 10666 22980 10718 23032
rect 10718 22980 10720 23032
rect 10664 22978 10720 22980
rect 10664 22815 10720 22817
rect 10664 22763 10666 22815
rect 10666 22763 10718 22815
rect 10718 22763 10720 22815
rect 10664 22761 10720 22763
rect 10986 24773 11042 24775
rect 10986 24721 10988 24773
rect 10988 24721 11040 24773
rect 11040 24721 11042 24773
rect 10986 24719 11042 24721
rect 10986 24556 11042 24558
rect 10986 24504 10988 24556
rect 10988 24504 11040 24556
rect 11040 24504 11042 24556
rect 10986 24502 11042 24504
rect 10986 24338 11042 24340
rect 10986 24286 10988 24338
rect 10988 24286 11040 24338
rect 11040 24286 11042 24338
rect 10986 24284 11042 24286
rect 10986 24121 11042 24123
rect 10986 24069 10988 24121
rect 10988 24069 11040 24121
rect 11040 24069 11042 24121
rect 10986 24067 11042 24069
rect 10986 23903 11042 23905
rect 10986 23851 10988 23903
rect 10988 23851 11040 23903
rect 11040 23851 11042 23903
rect 10986 23849 11042 23851
rect 10986 23685 11042 23687
rect 10986 23633 10988 23685
rect 10988 23633 11040 23685
rect 11040 23633 11042 23685
rect 10986 23631 11042 23633
rect 10986 23467 11042 23469
rect 10986 23415 10988 23467
rect 10988 23415 11040 23467
rect 11040 23415 11042 23467
rect 10986 23413 11042 23415
rect 10986 23250 11042 23252
rect 10986 23198 10988 23250
rect 10988 23198 11040 23250
rect 11040 23198 11042 23250
rect 10986 23196 11042 23198
rect 10986 23032 11042 23034
rect 10986 22980 10988 23032
rect 10988 22980 11040 23032
rect 11040 22980 11042 23032
rect 10986 22978 11042 22980
rect 10986 22815 11042 22817
rect 10986 22763 10988 22815
rect 10988 22763 11040 22815
rect 11040 22763 11042 22815
rect 10986 22761 11042 22763
rect 11438 24773 11494 24775
rect 11438 24721 11440 24773
rect 11440 24721 11492 24773
rect 11492 24721 11494 24773
rect 11438 24719 11494 24721
rect 11721 24773 11777 24775
rect 11721 24721 11723 24773
rect 11723 24721 11775 24773
rect 11775 24721 11777 24773
rect 11721 24719 11777 24721
rect 12004 24773 12060 24775
rect 12004 24721 12006 24773
rect 12006 24721 12058 24773
rect 12058 24721 12060 24773
rect 12004 24719 12060 24721
rect 11438 24556 11494 24558
rect 11438 24504 11440 24556
rect 11440 24504 11492 24556
rect 11492 24504 11494 24556
rect 11438 24502 11494 24504
rect 11721 24556 11777 24558
rect 11721 24504 11723 24556
rect 11723 24504 11775 24556
rect 11775 24504 11777 24556
rect 11721 24502 11777 24504
rect 12004 24556 12060 24558
rect 12004 24504 12006 24556
rect 12006 24504 12058 24556
rect 12058 24504 12060 24556
rect 12004 24502 12060 24504
rect 11438 24338 11494 24340
rect 11438 24286 11440 24338
rect 11440 24286 11492 24338
rect 11492 24286 11494 24338
rect 11438 24284 11494 24286
rect 11721 24338 11777 24340
rect 11721 24286 11723 24338
rect 11723 24286 11775 24338
rect 11775 24286 11777 24338
rect 11721 24284 11777 24286
rect 12004 24338 12060 24340
rect 12004 24286 12006 24338
rect 12006 24286 12058 24338
rect 12058 24286 12060 24338
rect 12004 24284 12060 24286
rect 11438 24121 11494 24123
rect 11438 24069 11440 24121
rect 11440 24069 11492 24121
rect 11492 24069 11494 24121
rect 11438 24067 11494 24069
rect 11721 24121 11777 24123
rect 11721 24069 11723 24121
rect 11723 24069 11775 24121
rect 11775 24069 11777 24121
rect 11721 24067 11777 24069
rect 12004 24121 12060 24123
rect 12004 24069 12006 24121
rect 12006 24069 12058 24121
rect 12058 24069 12060 24121
rect 12004 24067 12060 24069
rect 11438 23903 11494 23905
rect 11438 23851 11440 23903
rect 11440 23851 11492 23903
rect 11492 23851 11494 23903
rect 11438 23849 11494 23851
rect 11721 23903 11777 23905
rect 11721 23851 11723 23903
rect 11723 23851 11775 23903
rect 11775 23851 11777 23903
rect 11721 23849 11777 23851
rect 12004 23903 12060 23905
rect 12004 23851 12006 23903
rect 12006 23851 12058 23903
rect 12058 23851 12060 23903
rect 12004 23849 12060 23851
rect 11438 23685 11494 23687
rect 11438 23633 11440 23685
rect 11440 23633 11492 23685
rect 11492 23633 11494 23685
rect 11438 23631 11494 23633
rect 11721 23685 11777 23687
rect 11721 23633 11723 23685
rect 11723 23633 11775 23685
rect 11775 23633 11777 23685
rect 11721 23631 11777 23633
rect 12004 23685 12060 23687
rect 12004 23633 12006 23685
rect 12006 23633 12058 23685
rect 12058 23633 12060 23685
rect 12004 23631 12060 23633
rect 11438 23467 11494 23469
rect 11438 23415 11440 23467
rect 11440 23415 11492 23467
rect 11492 23415 11494 23467
rect 11438 23413 11494 23415
rect 11721 23467 11777 23469
rect 11721 23415 11723 23467
rect 11723 23415 11775 23467
rect 11775 23415 11777 23467
rect 11721 23413 11777 23415
rect 12004 23467 12060 23469
rect 12004 23415 12006 23467
rect 12006 23415 12058 23467
rect 12058 23415 12060 23467
rect 12004 23413 12060 23415
rect 11438 23250 11494 23252
rect 11438 23198 11440 23250
rect 11440 23198 11492 23250
rect 11492 23198 11494 23250
rect 11438 23196 11494 23198
rect 11721 23250 11777 23252
rect 11721 23198 11723 23250
rect 11723 23198 11775 23250
rect 11775 23198 11777 23250
rect 11721 23196 11777 23198
rect 12004 23250 12060 23252
rect 12004 23198 12006 23250
rect 12006 23198 12058 23250
rect 12058 23198 12060 23250
rect 12004 23196 12060 23198
rect 11438 23032 11494 23034
rect 11438 22980 11440 23032
rect 11440 22980 11492 23032
rect 11492 22980 11494 23032
rect 11438 22978 11494 22980
rect 11721 23032 11777 23034
rect 11721 22980 11723 23032
rect 11723 22980 11775 23032
rect 11775 22980 11777 23032
rect 11721 22978 11777 22980
rect 12004 23032 12060 23034
rect 12004 22980 12006 23032
rect 12006 22980 12058 23032
rect 12058 22980 12060 23032
rect 12004 22978 12060 22980
rect 11438 22815 11494 22817
rect 11438 22763 11440 22815
rect 11440 22763 11492 22815
rect 11492 22763 11494 22815
rect 11438 22761 11494 22763
rect 11721 22815 11777 22817
rect 11721 22763 11723 22815
rect 11723 22763 11775 22815
rect 11775 22763 11777 22815
rect 11721 22761 11777 22763
rect 12004 22815 12060 22817
rect 12004 22763 12006 22815
rect 12006 22763 12058 22815
rect 12058 22763 12060 22815
rect 12004 22761 12060 22763
rect 12456 24773 12512 24775
rect 12456 24721 12458 24773
rect 12458 24721 12510 24773
rect 12510 24721 12512 24773
rect 12456 24719 12512 24721
rect 12456 24556 12512 24558
rect 12456 24504 12458 24556
rect 12458 24504 12510 24556
rect 12510 24504 12512 24556
rect 12456 24502 12512 24504
rect 12456 24338 12512 24340
rect 12456 24286 12458 24338
rect 12458 24286 12510 24338
rect 12510 24286 12512 24338
rect 12456 24284 12512 24286
rect 12456 24121 12512 24123
rect 12456 24069 12458 24121
rect 12458 24069 12510 24121
rect 12510 24069 12512 24121
rect 12456 24067 12512 24069
rect 12456 23903 12512 23905
rect 12456 23851 12458 23903
rect 12458 23851 12510 23903
rect 12510 23851 12512 23903
rect 12456 23849 12512 23851
rect 12456 23685 12512 23687
rect 12456 23633 12458 23685
rect 12458 23633 12510 23685
rect 12510 23633 12512 23685
rect 12456 23631 12512 23633
rect 12456 23467 12512 23469
rect 12456 23415 12458 23467
rect 12458 23415 12510 23467
rect 12510 23415 12512 23467
rect 12456 23413 12512 23415
rect 12456 23250 12512 23252
rect 12456 23198 12458 23250
rect 12458 23198 12510 23250
rect 12510 23198 12512 23250
rect 12456 23196 12512 23198
rect 12456 23032 12512 23034
rect 12456 22980 12458 23032
rect 12458 22980 12510 23032
rect 12510 22980 12512 23032
rect 12456 22978 12512 22980
rect 12456 22815 12512 22817
rect 12456 22763 12458 22815
rect 12458 22763 12510 22815
rect 12510 22763 12512 22815
rect 12456 22761 12512 22763
rect 8776 21987 8832 22043
rect 8776 21769 8832 21825
rect 9646 20364 9702 20366
rect 9646 20312 9648 20364
rect 9648 20312 9700 20364
rect 9700 20312 9702 20364
rect 9646 20310 9702 20312
rect 9929 20364 9985 20366
rect 9929 20312 9931 20364
rect 9931 20312 9983 20364
rect 9983 20312 9985 20364
rect 9929 20310 9985 20312
rect 10212 20364 10268 20366
rect 10212 20312 10214 20364
rect 10214 20312 10266 20364
rect 10266 20312 10268 20364
rect 10212 20310 10268 20312
rect 9646 20146 9702 20148
rect 9646 20094 9648 20146
rect 9648 20094 9700 20146
rect 9700 20094 9702 20146
rect 9646 20092 9702 20094
rect 9929 20146 9985 20148
rect 9929 20094 9931 20146
rect 9931 20094 9983 20146
rect 9983 20094 9985 20146
rect 9929 20092 9985 20094
rect 10212 20146 10268 20148
rect 10212 20094 10214 20146
rect 10214 20094 10266 20146
rect 10266 20094 10268 20146
rect 10212 20092 10268 20094
rect 9646 19929 9702 19930
rect 9646 19877 9648 19929
rect 9648 19877 9700 19929
rect 9700 19877 9702 19929
rect 9646 19874 9702 19877
rect 9929 19929 9985 19930
rect 9929 19877 9931 19929
rect 9931 19877 9983 19929
rect 9983 19877 9985 19929
rect 9929 19874 9985 19877
rect 10212 19929 10268 19930
rect 10212 19877 10214 19929
rect 10214 19877 10266 19929
rect 10266 19877 10268 19929
rect 10212 19874 10268 19877
rect 4059 18405 4115 18408
rect 4059 18353 4061 18405
rect 4061 18353 4113 18405
rect 4113 18353 4115 18405
rect 4059 18352 4115 18353
rect 4342 18405 4398 18408
rect 4342 18353 4344 18405
rect 4344 18353 4396 18405
rect 4396 18353 4398 18405
rect 4342 18352 4398 18353
rect 4625 18405 4681 18408
rect 4625 18353 4627 18405
rect 4627 18353 4679 18405
rect 4679 18353 4681 18405
rect 4625 18352 4681 18353
rect 4059 18188 4115 18190
rect 4059 18136 4061 18188
rect 4061 18136 4113 18188
rect 4113 18136 4115 18188
rect 4059 18134 4115 18136
rect 4342 18188 4398 18190
rect 4342 18136 4344 18188
rect 4344 18136 4396 18188
rect 4396 18136 4398 18188
rect 4342 18134 4398 18136
rect 4625 18188 4681 18190
rect 4625 18136 4627 18188
rect 4627 18136 4679 18188
rect 4679 18136 4681 18188
rect 4625 18134 4681 18136
rect 4059 17970 4115 17972
rect 4059 17918 4061 17970
rect 4061 17918 4113 17970
rect 4113 17918 4115 17970
rect 4059 17916 4115 17918
rect 4342 17970 4398 17972
rect 4342 17918 4344 17970
rect 4344 17918 4396 17970
rect 4396 17918 4398 17970
rect 4342 17916 4398 17918
rect 4625 17970 4681 17972
rect 4625 17918 4627 17970
rect 4627 17918 4679 17970
rect 4679 17918 4681 17970
rect 4625 17916 4681 17918
rect 11438 20364 11494 20366
rect 11438 20312 11440 20364
rect 11440 20312 11492 20364
rect 11492 20312 11494 20364
rect 11438 20310 11494 20312
rect 11721 20364 11777 20366
rect 11721 20312 11723 20364
rect 11723 20312 11775 20364
rect 11775 20312 11777 20364
rect 11721 20310 11777 20312
rect 12004 20364 12060 20366
rect 12004 20312 12006 20364
rect 12006 20312 12058 20364
rect 12058 20312 12060 20364
rect 12004 20310 12060 20312
rect 11438 20146 11494 20148
rect 11438 20094 11440 20146
rect 11440 20094 11492 20146
rect 11492 20094 11494 20146
rect 11438 20092 11494 20094
rect 11721 20146 11777 20148
rect 11721 20094 11723 20146
rect 11723 20094 11775 20146
rect 11775 20094 11777 20146
rect 11721 20092 11777 20094
rect 12004 20146 12060 20148
rect 12004 20094 12006 20146
rect 12006 20094 12058 20146
rect 12058 20094 12060 20146
rect 12004 20092 12060 20094
rect 11438 19929 11494 19930
rect 11438 19877 11440 19929
rect 11440 19877 11492 19929
rect 11492 19877 11494 19929
rect 11438 19874 11494 19877
rect 11721 19929 11777 19930
rect 11721 19877 11723 19929
rect 11723 19877 11775 19929
rect 11775 19877 11777 19929
rect 11721 19874 11777 19877
rect 12004 19929 12060 19930
rect 12004 19877 12006 19929
rect 12006 19877 12058 19929
rect 12058 19877 12060 19929
rect 12004 19874 12060 19877
rect 9646 18405 9702 18408
rect 9646 18353 9648 18405
rect 9648 18353 9700 18405
rect 9700 18353 9702 18405
rect 9646 18352 9702 18353
rect 9929 18405 9985 18408
rect 9929 18353 9931 18405
rect 9931 18353 9983 18405
rect 9983 18353 9985 18405
rect 9929 18352 9985 18353
rect 10212 18405 10268 18408
rect 10212 18353 10214 18405
rect 10214 18353 10266 18405
rect 10266 18353 10268 18405
rect 10212 18352 10268 18353
rect 9646 18188 9702 18190
rect 9646 18136 9648 18188
rect 9648 18136 9700 18188
rect 9700 18136 9702 18188
rect 9646 18134 9702 18136
rect 9929 18188 9985 18190
rect 9929 18136 9931 18188
rect 9931 18136 9983 18188
rect 9983 18136 9985 18188
rect 9929 18134 9985 18136
rect 10212 18188 10268 18190
rect 10212 18136 10214 18188
rect 10214 18136 10266 18188
rect 10266 18136 10268 18188
rect 10212 18134 10268 18136
rect 9646 17970 9702 17972
rect 9646 17918 9648 17970
rect 9648 17918 9700 17970
rect 9700 17918 9702 17970
rect 9646 17916 9702 17918
rect 9929 17970 9985 17972
rect 9929 17918 9931 17970
rect 9931 17918 9983 17970
rect 9983 17918 9985 17970
rect 9929 17916 9985 17918
rect 10212 17970 10268 17972
rect 10212 17918 10214 17970
rect 10214 17918 10266 17970
rect 10266 17918 10268 17970
rect 10212 17916 10268 17918
rect 4059 17698 4115 17754
rect 4342 17698 4398 17754
rect 4625 17698 4681 17754
rect 9646 17698 9702 17754
rect 9929 17698 9985 17754
rect 10212 17698 10268 17754
rect 13471 24802 13527 24804
rect 13471 24750 13473 24802
rect 13473 24750 13525 24802
rect 13525 24750 13527 24802
rect 13471 24748 13527 24750
rect 13471 24585 13527 24587
rect 13471 24533 13473 24585
rect 13473 24533 13525 24585
rect 13525 24533 13527 24585
rect 13471 24531 13527 24533
rect 13471 24367 13527 24369
rect 13471 24315 13473 24367
rect 13473 24315 13525 24367
rect 13525 24315 13527 24367
rect 13471 24313 13527 24315
rect 13471 24150 13527 24152
rect 13471 24098 13473 24150
rect 13473 24098 13525 24150
rect 13525 24098 13527 24150
rect 13471 24096 13527 24098
rect 13471 23932 13527 23934
rect 13471 23880 13473 23932
rect 13473 23880 13525 23932
rect 13525 23880 13527 23932
rect 13471 23878 13527 23880
rect 13471 23714 13527 23716
rect 13471 23662 13473 23714
rect 13473 23662 13525 23714
rect 13525 23662 13527 23714
rect 13471 23660 13527 23662
rect 13471 23496 13527 23498
rect 13471 23444 13473 23496
rect 13473 23444 13525 23496
rect 13525 23444 13527 23496
rect 13471 23442 13527 23444
rect 13471 23279 13527 23281
rect 13471 23227 13473 23279
rect 13473 23227 13525 23279
rect 13525 23227 13527 23279
rect 13471 23225 13527 23227
rect 13985 24811 14041 24813
rect 13985 24759 13987 24811
rect 13987 24759 14039 24811
rect 14039 24759 14041 24811
rect 13985 24757 14041 24759
rect 13985 24593 14041 24595
rect 13985 24541 13987 24593
rect 13987 24541 14039 24593
rect 14039 24541 14041 24593
rect 13985 24539 14041 24541
rect 13985 24376 14041 24378
rect 13985 24324 13987 24376
rect 13987 24324 14039 24376
rect 14039 24324 14041 24376
rect 13985 24322 14041 24324
rect 13985 24158 14041 24160
rect 13985 24106 13987 24158
rect 13987 24106 14039 24158
rect 14039 24106 14041 24158
rect 13985 24104 14041 24106
rect 13985 23940 14041 23942
rect 13985 23888 13987 23940
rect 13987 23888 14039 23940
rect 14039 23888 14041 23940
rect 13985 23886 14041 23888
rect 13985 23722 14041 23724
rect 13985 23670 13987 23722
rect 13987 23670 14039 23722
rect 14039 23670 14041 23722
rect 13985 23668 14041 23670
rect 13985 23505 14041 23507
rect 13985 23453 13987 23505
rect 13987 23453 14039 23505
rect 14039 23453 14041 23505
rect 13985 23451 14041 23453
rect 13985 23287 14041 23289
rect 13985 23235 13987 23287
rect 13987 23235 14039 23287
rect 14039 23235 14041 23287
rect 13985 23233 14041 23235
rect 13471 23061 13527 23063
rect 13471 23009 13473 23061
rect 13473 23009 13525 23061
rect 13525 23009 13527 23061
rect 13471 23007 13527 23009
rect 14942 26514 14998 26516
rect 14942 26462 14944 26514
rect 14944 26462 14996 26514
rect 14996 26462 14998 26514
rect 14942 26460 14998 26462
rect 15149 26514 15205 26516
rect 15149 26462 15151 26514
rect 15151 26462 15203 26514
rect 15203 26462 15205 26514
rect 15149 26460 15205 26462
rect 14942 26296 14998 26298
rect 14942 26244 14944 26296
rect 14944 26244 14996 26296
rect 14996 26244 14998 26296
rect 14942 26242 14998 26244
rect 15149 26296 15205 26298
rect 15149 26244 15151 26296
rect 15151 26244 15203 26296
rect 15203 26244 15205 26296
rect 15149 26242 15205 26244
rect 14942 26078 14998 26080
rect 14942 26026 14944 26078
rect 14944 26026 14996 26078
rect 14996 26026 14998 26078
rect 14942 26024 14998 26026
rect 15149 26078 15205 26080
rect 15149 26026 15151 26078
rect 15151 26026 15203 26078
rect 15203 26026 15205 26078
rect 15149 26024 15205 26026
rect 14942 25860 14998 25862
rect 14942 25808 14944 25860
rect 14944 25808 14996 25860
rect 14996 25808 14998 25860
rect 14942 25806 14998 25808
rect 15149 25860 15205 25862
rect 15149 25808 15151 25860
rect 15151 25808 15203 25860
rect 15203 25808 15205 25860
rect 15149 25806 15205 25808
rect 15669 26491 15725 26493
rect 15669 26439 15671 26491
rect 15671 26439 15723 26491
rect 15723 26439 15725 26491
rect 15669 26437 15725 26439
rect 15669 26273 15725 26275
rect 15669 26221 15671 26273
rect 15671 26221 15723 26273
rect 15723 26221 15725 26273
rect 15669 26219 15725 26221
rect 15669 26055 15725 26057
rect 15669 26003 15671 26055
rect 15671 26003 15723 26055
rect 15723 26003 15725 26055
rect 15669 26001 15725 26003
rect 15669 25837 15725 25839
rect 15669 25785 15671 25837
rect 15671 25785 15723 25837
rect 15723 25785 15725 25837
rect 15669 25783 15725 25785
rect 13471 22844 13527 22846
rect 13471 22792 13473 22844
rect 13473 22792 13525 22844
rect 13525 22792 13527 22844
rect 13471 22790 13527 22792
rect 13974 21511 14030 21567
rect 13974 21293 14030 21349
rect 14464 21987 14520 22043
rect 14464 21769 14520 21825
rect 15162 24802 15218 24804
rect 15162 24750 15164 24802
rect 15164 24750 15216 24802
rect 15216 24750 15218 24802
rect 15162 24748 15218 24750
rect 15162 24585 15218 24587
rect 15162 24533 15164 24585
rect 15164 24533 15216 24585
rect 15216 24533 15218 24585
rect 15162 24531 15218 24533
rect 15162 24367 15218 24369
rect 15162 24315 15164 24367
rect 15164 24315 15216 24367
rect 15216 24315 15218 24367
rect 15162 24313 15218 24315
rect 15162 24150 15218 24152
rect 15162 24098 15164 24150
rect 15164 24098 15216 24150
rect 15216 24098 15218 24150
rect 15162 24096 15218 24098
rect 15162 23932 15218 23934
rect 15162 23880 15164 23932
rect 15164 23880 15216 23932
rect 15216 23880 15218 23932
rect 15162 23878 15218 23880
rect 15162 23714 15218 23716
rect 15162 23662 15164 23714
rect 15164 23662 15216 23714
rect 15216 23662 15218 23714
rect 15162 23660 15218 23662
rect 15162 23496 15218 23498
rect 15162 23444 15164 23496
rect 15164 23444 15216 23496
rect 15216 23444 15218 23496
rect 15162 23442 15218 23444
rect 15162 23279 15218 23281
rect 15162 23227 15164 23279
rect 15164 23227 15216 23279
rect 15216 23227 15218 23279
rect 15162 23225 15218 23227
rect 15676 24811 15732 24813
rect 15676 24759 15678 24811
rect 15678 24759 15730 24811
rect 15730 24759 15732 24811
rect 15676 24757 15732 24759
rect 15676 24593 15732 24595
rect 15676 24541 15678 24593
rect 15678 24541 15730 24593
rect 15730 24541 15732 24593
rect 15676 24539 15732 24541
rect 15676 24376 15732 24378
rect 15676 24324 15678 24376
rect 15678 24324 15730 24376
rect 15730 24324 15732 24376
rect 15676 24322 15732 24324
rect 15676 24158 15732 24160
rect 15676 24106 15678 24158
rect 15678 24106 15730 24158
rect 15730 24106 15732 24158
rect 15676 24104 15732 24106
rect 15676 23940 15732 23942
rect 15676 23888 15678 23940
rect 15678 23888 15730 23940
rect 15730 23888 15732 23940
rect 15676 23886 15732 23888
rect 15676 23722 15732 23724
rect 15676 23670 15678 23722
rect 15678 23670 15730 23722
rect 15730 23670 15732 23722
rect 15676 23668 15732 23670
rect 15676 23505 15732 23507
rect 15676 23453 15678 23505
rect 15678 23453 15730 23505
rect 15730 23453 15732 23505
rect 15676 23451 15732 23453
rect 15676 23287 15732 23289
rect 15676 23235 15678 23287
rect 15678 23235 15730 23287
rect 15730 23235 15732 23287
rect 15676 23233 15732 23235
rect 15162 23061 15218 23063
rect 15162 23009 15164 23061
rect 15164 23009 15216 23061
rect 15216 23009 15218 23061
rect 15162 23007 15218 23009
rect 15162 22844 15218 22846
rect 15162 22792 15164 22844
rect 15164 22792 15216 22844
rect 15216 22792 15218 22844
rect 15162 22790 15218 22792
rect 15665 21511 15721 21567
rect 15665 21293 15721 21349
rect 23785 27378 23841 27380
rect 23785 27326 23787 27378
rect 23787 27326 23839 27378
rect 23839 27326 23841 27378
rect 23785 27324 23841 27326
rect 23785 27160 23841 27162
rect 23785 27108 23787 27160
rect 23787 27108 23839 27160
rect 23839 27108 23841 27160
rect 23785 27106 23841 27108
rect 24971 27437 25027 27439
rect 24971 27385 24973 27437
rect 24973 27385 25025 27437
rect 25025 27385 25027 27437
rect 24971 27383 25027 27385
rect 24971 27219 25027 27221
rect 24971 27167 24973 27219
rect 24973 27167 25025 27219
rect 25025 27167 25027 27219
rect 24971 27165 25027 27167
rect 25999 27392 26055 27394
rect 25999 27340 26001 27392
rect 26001 27340 26053 27392
rect 26053 27340 26055 27392
rect 25999 27338 26055 27340
rect 25999 27174 26055 27176
rect 25999 27122 26001 27174
rect 26001 27122 26053 27174
rect 26053 27122 26055 27174
rect 25999 27120 26055 27122
rect 23737 26535 23793 26537
rect 23737 26483 23739 26535
rect 23739 26483 23791 26535
rect 23791 26483 23793 26535
rect 23737 26481 23793 26483
rect 23944 26535 24000 26537
rect 23944 26483 23946 26535
rect 23946 26483 23998 26535
rect 23998 26483 24000 26535
rect 23944 26481 24000 26483
rect 23737 26317 23793 26319
rect 23737 26265 23739 26317
rect 23739 26265 23791 26317
rect 23791 26265 23793 26317
rect 23737 26263 23793 26265
rect 23944 26317 24000 26319
rect 23944 26265 23946 26317
rect 23946 26265 23998 26317
rect 23998 26265 24000 26317
rect 23944 26263 24000 26265
rect 23737 26099 23793 26101
rect 23737 26047 23739 26099
rect 23739 26047 23791 26099
rect 23791 26047 23793 26099
rect 23737 26045 23793 26047
rect 23944 26099 24000 26101
rect 23944 26047 23946 26099
rect 23946 26047 23998 26099
rect 23998 26047 24000 26099
rect 23944 26045 24000 26047
rect 23737 25881 23793 25883
rect 23737 25829 23739 25881
rect 23739 25829 23791 25881
rect 23791 25829 23793 25881
rect 23737 25827 23793 25829
rect 23944 25881 24000 25883
rect 23944 25829 23946 25881
rect 23946 25829 23998 25881
rect 23998 25829 24000 25881
rect 23944 25827 24000 25829
rect 24464 26535 24520 26537
rect 24464 26483 24466 26535
rect 24466 26483 24518 26535
rect 24518 26483 24520 26535
rect 24464 26481 24520 26483
rect 24464 26317 24520 26319
rect 24464 26265 24466 26317
rect 24466 26265 24518 26317
rect 24518 26265 24520 26317
rect 24464 26263 24520 26265
rect 24464 26099 24520 26101
rect 24464 26047 24466 26099
rect 24466 26047 24518 26099
rect 24518 26047 24520 26099
rect 24464 26045 24520 26047
rect 24464 25881 24520 25883
rect 24464 25829 24466 25881
rect 24466 25829 24518 25881
rect 24518 25829 24520 25881
rect 24464 25827 24520 25829
rect 16923 25300 16979 25302
rect 16923 25248 16925 25300
rect 16925 25248 16977 25300
rect 16977 25248 16979 25300
rect 16923 25246 16979 25248
rect 16923 25082 16979 25084
rect 16923 25030 16925 25082
rect 16925 25030 16977 25082
rect 16977 25030 16979 25082
rect 16923 25028 16979 25030
rect 16923 24864 16979 24866
rect 16923 24812 16925 24864
rect 16925 24812 16977 24864
rect 16977 24812 16979 24864
rect 16923 24810 16979 24812
rect 17371 25300 17427 25302
rect 17371 25248 17373 25300
rect 17373 25248 17425 25300
rect 17425 25248 17427 25300
rect 17371 25246 17427 25248
rect 17371 25082 17427 25084
rect 17371 25030 17373 25082
rect 17373 25030 17425 25082
rect 17425 25030 17427 25082
rect 17371 25028 17427 25030
rect 17371 24864 17427 24866
rect 17371 24812 17373 24864
rect 17373 24812 17425 24864
rect 17425 24812 17427 24864
rect 17371 24810 17427 24812
rect 17819 25300 17875 25302
rect 17819 25248 17821 25300
rect 17821 25248 17873 25300
rect 17873 25248 17875 25300
rect 17819 25246 17875 25248
rect 17819 25082 17875 25084
rect 17819 25030 17821 25082
rect 17821 25030 17873 25082
rect 17873 25030 17875 25082
rect 17819 25028 17875 25030
rect 17819 24864 17875 24866
rect 17819 24812 17821 24864
rect 17821 24812 17873 24864
rect 17873 24812 17875 24864
rect 17819 24810 17875 24812
rect 18557 25300 18613 25302
rect 18557 25248 18559 25300
rect 18559 25248 18611 25300
rect 18611 25248 18613 25300
rect 18557 25246 18613 25248
rect 18557 25082 18613 25084
rect 18557 25030 18559 25082
rect 18559 25030 18611 25082
rect 18611 25030 18613 25082
rect 18557 25028 18613 25030
rect 18557 24864 18613 24866
rect 18557 24812 18559 24864
rect 18559 24812 18611 24864
rect 18611 24812 18613 24864
rect 18557 24810 18613 24812
rect 19005 25300 19061 25302
rect 19005 25248 19007 25300
rect 19007 25248 19059 25300
rect 19059 25248 19061 25300
rect 19005 25246 19061 25248
rect 19005 25082 19061 25084
rect 19005 25030 19007 25082
rect 19007 25030 19059 25082
rect 19059 25030 19061 25082
rect 19005 25028 19061 25030
rect 19005 24864 19061 24866
rect 19005 24812 19007 24864
rect 19007 24812 19059 24864
rect 19059 24812 19061 24864
rect 19005 24810 19061 24812
rect 19453 25300 19509 25302
rect 19453 25248 19455 25300
rect 19455 25248 19507 25300
rect 19507 25248 19509 25300
rect 19453 25246 19509 25248
rect 19453 25082 19509 25084
rect 19453 25030 19455 25082
rect 19455 25030 19507 25082
rect 19507 25030 19509 25082
rect 19453 25028 19509 25030
rect 19453 24864 19509 24866
rect 19453 24812 19455 24864
rect 19455 24812 19507 24864
rect 19507 24812 19509 24864
rect 19453 24810 19509 24812
rect 20190 25300 20246 25302
rect 20190 25248 20192 25300
rect 20192 25248 20244 25300
rect 20244 25248 20246 25300
rect 20190 25246 20246 25248
rect 20190 25082 20246 25084
rect 20190 25030 20192 25082
rect 20192 25030 20244 25082
rect 20244 25030 20246 25082
rect 20190 25028 20246 25030
rect 20190 24864 20246 24866
rect 20190 24812 20192 24864
rect 20192 24812 20244 24864
rect 20244 24812 20246 24864
rect 20190 24810 20246 24812
rect 20638 25300 20694 25302
rect 20638 25248 20640 25300
rect 20640 25248 20692 25300
rect 20692 25248 20694 25300
rect 20638 25246 20694 25248
rect 20638 25082 20694 25084
rect 20638 25030 20640 25082
rect 20640 25030 20692 25082
rect 20692 25030 20694 25082
rect 20638 25028 20694 25030
rect 20638 24864 20694 24866
rect 20638 24812 20640 24864
rect 20640 24812 20692 24864
rect 20692 24812 20694 24864
rect 20638 24810 20694 24812
rect 21086 25300 21142 25302
rect 21086 25248 21088 25300
rect 21088 25248 21140 25300
rect 21140 25248 21142 25300
rect 21086 25246 21142 25248
rect 21086 25082 21142 25084
rect 21086 25030 21088 25082
rect 21088 25030 21140 25082
rect 21140 25030 21142 25082
rect 21086 25028 21142 25030
rect 21086 24864 21142 24866
rect 21086 24812 21088 24864
rect 21088 24812 21140 24864
rect 21140 24812 21142 24864
rect 21086 24810 21142 24812
rect 21824 25300 21880 25302
rect 21824 25248 21826 25300
rect 21826 25248 21878 25300
rect 21878 25248 21880 25300
rect 21824 25246 21880 25248
rect 21824 25082 21880 25084
rect 21824 25030 21826 25082
rect 21826 25030 21878 25082
rect 21878 25030 21880 25082
rect 21824 25028 21880 25030
rect 21824 24864 21880 24866
rect 21824 24812 21826 24864
rect 21826 24812 21878 24864
rect 21878 24812 21880 24864
rect 21824 24810 21880 24812
rect 22272 25300 22328 25302
rect 22272 25248 22274 25300
rect 22274 25248 22326 25300
rect 22326 25248 22328 25300
rect 22272 25246 22328 25248
rect 22272 25082 22328 25084
rect 22272 25030 22274 25082
rect 22274 25030 22326 25082
rect 22326 25030 22328 25082
rect 22272 25028 22328 25030
rect 22272 24864 22328 24866
rect 22272 24812 22274 24864
rect 22274 24812 22326 24864
rect 22326 24812 22328 24864
rect 22272 24810 22328 24812
rect 22720 25300 22776 25302
rect 22720 25248 22722 25300
rect 22722 25248 22774 25300
rect 22774 25248 22776 25300
rect 22720 25246 22776 25248
rect 22720 25082 22776 25084
rect 22720 25030 22722 25082
rect 22722 25030 22774 25082
rect 22774 25030 22776 25082
rect 22720 25028 22776 25030
rect 22720 24864 22776 24866
rect 22720 24812 22722 24864
rect 22722 24812 22774 24864
rect 22774 24812 22776 24864
rect 22720 24810 22776 24812
rect 16927 24180 16983 24182
rect 16927 24128 16929 24180
rect 16929 24128 16981 24180
rect 16981 24128 16983 24180
rect 16927 24126 16983 24128
rect 16927 23962 16983 23964
rect 16927 23910 16929 23962
rect 16929 23910 16981 23962
rect 16981 23910 16983 23962
rect 16927 23908 16983 23910
rect 16927 23745 16983 23747
rect 16927 23693 16929 23745
rect 16929 23693 16981 23745
rect 16981 23693 16983 23745
rect 16927 23691 16983 23693
rect 16927 23527 16983 23529
rect 16927 23475 16929 23527
rect 16929 23475 16981 23527
rect 16981 23475 16983 23527
rect 16927 23473 16983 23475
rect 16927 23309 16983 23311
rect 16927 23257 16929 23309
rect 16929 23257 16981 23309
rect 16981 23257 16983 23309
rect 16927 23255 16983 23257
rect 16927 23092 16983 23094
rect 16927 23040 16929 23092
rect 16929 23040 16981 23092
rect 16981 23040 16983 23092
rect 16927 23038 16983 23040
rect 16927 22874 16983 22876
rect 16927 22822 16929 22874
rect 16929 22822 16981 22874
rect 16981 22822 16983 22874
rect 16927 22820 16983 22822
rect 17371 24180 17427 24182
rect 17371 24128 17373 24180
rect 17373 24128 17425 24180
rect 17425 24128 17427 24180
rect 17371 24126 17427 24128
rect 17371 23962 17427 23964
rect 17371 23910 17373 23962
rect 17373 23910 17425 23962
rect 17425 23910 17427 23962
rect 17371 23908 17427 23910
rect 17371 23745 17427 23747
rect 17371 23693 17373 23745
rect 17373 23693 17425 23745
rect 17425 23693 17427 23745
rect 17371 23691 17427 23693
rect 17371 23527 17427 23529
rect 17371 23475 17373 23527
rect 17373 23475 17425 23527
rect 17425 23475 17427 23527
rect 17371 23473 17427 23475
rect 17371 23309 17427 23311
rect 17371 23257 17373 23309
rect 17373 23257 17425 23309
rect 17425 23257 17427 23309
rect 17371 23255 17427 23257
rect 17371 23092 17427 23094
rect 17371 23040 17373 23092
rect 17373 23040 17425 23092
rect 17425 23040 17427 23092
rect 17371 23038 17427 23040
rect 17371 22874 17427 22876
rect 17371 22822 17373 22874
rect 17373 22822 17425 22874
rect 17425 22822 17427 22874
rect 17371 22820 17427 22822
rect 17815 24180 17871 24182
rect 17815 24128 17817 24180
rect 17817 24128 17869 24180
rect 17869 24128 17871 24180
rect 17815 24126 17871 24128
rect 17815 23962 17871 23964
rect 17815 23910 17817 23962
rect 17817 23910 17869 23962
rect 17869 23910 17871 23962
rect 17815 23908 17871 23910
rect 17815 23745 17871 23747
rect 17815 23693 17817 23745
rect 17817 23693 17869 23745
rect 17869 23693 17871 23745
rect 17815 23691 17871 23693
rect 17815 23527 17871 23529
rect 17815 23475 17817 23527
rect 17817 23475 17869 23527
rect 17869 23475 17871 23527
rect 17815 23473 17871 23475
rect 17815 23309 17871 23311
rect 17815 23257 17817 23309
rect 17817 23257 17869 23309
rect 17869 23257 17871 23309
rect 17815 23255 17871 23257
rect 17815 23092 17871 23094
rect 17815 23040 17817 23092
rect 17817 23040 17869 23092
rect 17869 23040 17871 23092
rect 17815 23038 17871 23040
rect 17815 22874 17871 22876
rect 17815 22822 17817 22874
rect 17817 22822 17869 22874
rect 17869 22822 17871 22874
rect 17815 22820 17871 22822
rect 18561 24180 18617 24182
rect 18561 24128 18563 24180
rect 18563 24128 18615 24180
rect 18615 24128 18617 24180
rect 18561 24126 18617 24128
rect 18561 23962 18617 23964
rect 18561 23910 18563 23962
rect 18563 23910 18615 23962
rect 18615 23910 18617 23962
rect 18561 23908 18617 23910
rect 18561 23745 18617 23747
rect 18561 23693 18563 23745
rect 18563 23693 18615 23745
rect 18615 23693 18617 23745
rect 18561 23691 18617 23693
rect 18561 23527 18617 23529
rect 18561 23475 18563 23527
rect 18563 23475 18615 23527
rect 18615 23475 18617 23527
rect 18561 23473 18617 23475
rect 18561 23309 18617 23311
rect 18561 23257 18563 23309
rect 18563 23257 18615 23309
rect 18615 23257 18617 23309
rect 18561 23255 18617 23257
rect 18561 23092 18617 23094
rect 18561 23040 18563 23092
rect 18563 23040 18615 23092
rect 18615 23040 18617 23092
rect 18561 23038 18617 23040
rect 18561 22874 18617 22876
rect 18561 22822 18563 22874
rect 18563 22822 18615 22874
rect 18615 22822 18617 22874
rect 18561 22820 18617 22822
rect 19005 24180 19061 24182
rect 19005 24128 19007 24180
rect 19007 24128 19059 24180
rect 19059 24128 19061 24180
rect 19005 24126 19061 24128
rect 19005 23962 19061 23964
rect 19005 23910 19007 23962
rect 19007 23910 19059 23962
rect 19059 23910 19061 23962
rect 19005 23908 19061 23910
rect 19005 23745 19061 23747
rect 19005 23693 19007 23745
rect 19007 23693 19059 23745
rect 19059 23693 19061 23745
rect 19005 23691 19061 23693
rect 19005 23527 19061 23529
rect 19005 23475 19007 23527
rect 19007 23475 19059 23527
rect 19059 23475 19061 23527
rect 19005 23473 19061 23475
rect 19005 23309 19061 23311
rect 19005 23257 19007 23309
rect 19007 23257 19059 23309
rect 19059 23257 19061 23309
rect 19005 23255 19061 23257
rect 19005 23092 19061 23094
rect 19005 23040 19007 23092
rect 19007 23040 19059 23092
rect 19059 23040 19061 23092
rect 19005 23038 19061 23040
rect 19005 22874 19061 22876
rect 19005 22822 19007 22874
rect 19007 22822 19059 22874
rect 19059 22822 19061 22874
rect 19005 22820 19061 22822
rect 19449 24180 19505 24182
rect 19449 24128 19451 24180
rect 19451 24128 19503 24180
rect 19503 24128 19505 24180
rect 19449 24126 19505 24128
rect 19449 23962 19505 23964
rect 19449 23910 19451 23962
rect 19451 23910 19503 23962
rect 19503 23910 19505 23962
rect 19449 23908 19505 23910
rect 19449 23745 19505 23747
rect 19449 23693 19451 23745
rect 19451 23693 19503 23745
rect 19503 23693 19505 23745
rect 19449 23691 19505 23693
rect 19449 23527 19505 23529
rect 19449 23475 19451 23527
rect 19451 23475 19503 23527
rect 19503 23475 19505 23527
rect 19449 23473 19505 23475
rect 19449 23309 19505 23311
rect 19449 23257 19451 23309
rect 19451 23257 19503 23309
rect 19503 23257 19505 23309
rect 19449 23255 19505 23257
rect 19449 23092 19505 23094
rect 19449 23040 19451 23092
rect 19451 23040 19503 23092
rect 19503 23040 19505 23092
rect 19449 23038 19505 23040
rect 19449 22874 19505 22876
rect 19449 22822 19451 22874
rect 19451 22822 19503 22874
rect 19503 22822 19505 22874
rect 19449 22820 19505 22822
rect 20194 24180 20250 24182
rect 20194 24128 20196 24180
rect 20196 24128 20248 24180
rect 20248 24128 20250 24180
rect 20194 24126 20250 24128
rect 20194 23962 20250 23964
rect 20194 23910 20196 23962
rect 20196 23910 20248 23962
rect 20248 23910 20250 23962
rect 20194 23908 20250 23910
rect 20194 23745 20250 23747
rect 20194 23693 20196 23745
rect 20196 23693 20248 23745
rect 20248 23693 20250 23745
rect 20194 23691 20250 23693
rect 20194 23527 20250 23529
rect 20194 23475 20196 23527
rect 20196 23475 20248 23527
rect 20248 23475 20250 23527
rect 20194 23473 20250 23475
rect 20194 23309 20250 23311
rect 20194 23257 20196 23309
rect 20196 23257 20248 23309
rect 20248 23257 20250 23309
rect 20194 23255 20250 23257
rect 20194 23092 20250 23094
rect 20194 23040 20196 23092
rect 20196 23040 20248 23092
rect 20248 23040 20250 23092
rect 20194 23038 20250 23040
rect 20194 22874 20250 22876
rect 20194 22822 20196 22874
rect 20196 22822 20248 22874
rect 20248 22822 20250 22874
rect 20194 22820 20250 22822
rect 20638 24180 20694 24182
rect 20638 24128 20640 24180
rect 20640 24128 20692 24180
rect 20692 24128 20694 24180
rect 20638 24126 20694 24128
rect 20638 23962 20694 23964
rect 20638 23910 20640 23962
rect 20640 23910 20692 23962
rect 20692 23910 20694 23962
rect 20638 23908 20694 23910
rect 20638 23745 20694 23747
rect 20638 23693 20640 23745
rect 20640 23693 20692 23745
rect 20692 23693 20694 23745
rect 20638 23691 20694 23693
rect 20638 23527 20694 23529
rect 20638 23475 20640 23527
rect 20640 23475 20692 23527
rect 20692 23475 20694 23527
rect 20638 23473 20694 23475
rect 20638 23309 20694 23311
rect 20638 23257 20640 23309
rect 20640 23257 20692 23309
rect 20692 23257 20694 23309
rect 20638 23255 20694 23257
rect 20638 23092 20694 23094
rect 20638 23040 20640 23092
rect 20640 23040 20692 23092
rect 20692 23040 20694 23092
rect 20638 23038 20694 23040
rect 20638 22874 20694 22876
rect 20638 22822 20640 22874
rect 20640 22822 20692 22874
rect 20692 22822 20694 22874
rect 20638 22820 20694 22822
rect 21082 24180 21138 24182
rect 21082 24128 21084 24180
rect 21084 24128 21136 24180
rect 21136 24128 21138 24180
rect 21082 24126 21138 24128
rect 21082 23962 21138 23964
rect 21082 23910 21084 23962
rect 21084 23910 21136 23962
rect 21136 23910 21138 23962
rect 21082 23908 21138 23910
rect 21082 23745 21138 23747
rect 21082 23693 21084 23745
rect 21084 23693 21136 23745
rect 21136 23693 21138 23745
rect 21082 23691 21138 23693
rect 21082 23527 21138 23529
rect 21082 23475 21084 23527
rect 21084 23475 21136 23527
rect 21136 23475 21138 23527
rect 21082 23473 21138 23475
rect 21082 23309 21138 23311
rect 21082 23257 21084 23309
rect 21084 23257 21136 23309
rect 21136 23257 21138 23309
rect 21082 23255 21138 23257
rect 21082 23092 21138 23094
rect 21082 23040 21084 23092
rect 21084 23040 21136 23092
rect 21136 23040 21138 23092
rect 21082 23038 21138 23040
rect 21082 22874 21138 22876
rect 21082 22822 21084 22874
rect 21084 22822 21136 22874
rect 21136 22822 21138 22874
rect 21082 22820 21138 22822
rect 21828 24180 21884 24182
rect 21828 24128 21830 24180
rect 21830 24128 21882 24180
rect 21882 24128 21884 24180
rect 21828 24126 21884 24128
rect 21828 23962 21884 23964
rect 21828 23910 21830 23962
rect 21830 23910 21882 23962
rect 21882 23910 21884 23962
rect 21828 23908 21884 23910
rect 21828 23745 21884 23747
rect 21828 23693 21830 23745
rect 21830 23693 21882 23745
rect 21882 23693 21884 23745
rect 21828 23691 21884 23693
rect 21828 23527 21884 23529
rect 21828 23475 21830 23527
rect 21830 23475 21882 23527
rect 21882 23475 21884 23527
rect 21828 23473 21884 23475
rect 21828 23309 21884 23311
rect 21828 23257 21830 23309
rect 21830 23257 21882 23309
rect 21882 23257 21884 23309
rect 21828 23255 21884 23257
rect 21828 23092 21884 23094
rect 21828 23040 21830 23092
rect 21830 23040 21882 23092
rect 21882 23040 21884 23092
rect 21828 23038 21884 23040
rect 21828 22874 21884 22876
rect 21828 22822 21830 22874
rect 21830 22822 21882 22874
rect 21882 22822 21884 22874
rect 21828 22820 21884 22822
rect 22272 24180 22328 24182
rect 22272 24128 22274 24180
rect 22274 24128 22326 24180
rect 22326 24128 22328 24180
rect 22272 24126 22328 24128
rect 22272 23962 22328 23964
rect 22272 23910 22274 23962
rect 22274 23910 22326 23962
rect 22326 23910 22328 23962
rect 22272 23908 22328 23910
rect 22272 23745 22328 23747
rect 22272 23693 22274 23745
rect 22274 23693 22326 23745
rect 22326 23693 22328 23745
rect 22272 23691 22328 23693
rect 22272 23527 22328 23529
rect 22272 23475 22274 23527
rect 22274 23475 22326 23527
rect 22326 23475 22328 23527
rect 22272 23473 22328 23475
rect 22272 23309 22328 23311
rect 22272 23257 22274 23309
rect 22274 23257 22326 23309
rect 22326 23257 22328 23309
rect 22272 23255 22328 23257
rect 22272 23092 22328 23094
rect 22272 23040 22274 23092
rect 22274 23040 22326 23092
rect 22326 23040 22328 23092
rect 22272 23038 22328 23040
rect 22272 22874 22328 22876
rect 22272 22822 22274 22874
rect 22274 22822 22326 22874
rect 22326 22822 22328 22874
rect 22272 22820 22328 22822
rect 22716 24180 22772 24182
rect 22716 24128 22718 24180
rect 22718 24128 22770 24180
rect 22770 24128 22772 24180
rect 22716 24126 22772 24128
rect 22716 23962 22772 23964
rect 22716 23910 22718 23962
rect 22718 23910 22770 23962
rect 22770 23910 22772 23962
rect 22716 23908 22772 23910
rect 22716 23745 22772 23747
rect 22716 23693 22718 23745
rect 22718 23693 22770 23745
rect 22770 23693 22772 23745
rect 22716 23691 22772 23693
rect 22716 23527 22772 23529
rect 22716 23475 22718 23527
rect 22718 23475 22770 23527
rect 22770 23475 22772 23527
rect 22716 23473 22772 23475
rect 22716 23309 22772 23311
rect 22716 23257 22718 23309
rect 22718 23257 22770 23309
rect 22770 23257 22772 23309
rect 22716 23255 22772 23257
rect 22716 23092 22772 23094
rect 22716 23040 22718 23092
rect 22718 23040 22770 23092
rect 22770 23040 22772 23092
rect 22716 23038 22772 23040
rect 22716 22874 22772 22876
rect 22716 22822 22718 22874
rect 22718 22822 22770 22874
rect 22770 22822 22772 22874
rect 22716 22820 22772 22822
rect 16155 21987 16211 22043
rect 16155 21769 16211 21825
rect 17371 20385 17427 20387
rect 17371 20333 17373 20385
rect 17373 20333 17425 20385
rect 17425 20333 17427 20385
rect 17371 20331 17427 20333
rect 17371 20167 17427 20169
rect 17371 20115 17373 20167
rect 17373 20115 17425 20167
rect 17425 20115 17427 20167
rect 17371 20113 17427 20115
rect 17371 19950 17427 19951
rect 17371 19898 17373 19950
rect 17373 19898 17425 19950
rect 17425 19898 17427 19950
rect 17371 19895 17427 19898
rect 11438 18405 11494 18408
rect 11438 18353 11440 18405
rect 11440 18353 11492 18405
rect 11492 18353 11494 18405
rect 11438 18352 11494 18353
rect 11721 18405 11777 18408
rect 11721 18353 11723 18405
rect 11723 18353 11775 18405
rect 11775 18353 11777 18405
rect 11721 18352 11777 18353
rect 12004 18405 12060 18408
rect 12004 18353 12006 18405
rect 12006 18353 12058 18405
rect 12058 18353 12060 18405
rect 12004 18352 12060 18353
rect 11438 18188 11494 18190
rect 11438 18136 11440 18188
rect 11440 18136 11492 18188
rect 11492 18136 11494 18188
rect 11438 18134 11494 18136
rect 11721 18188 11777 18190
rect 11721 18136 11723 18188
rect 11723 18136 11775 18188
rect 11775 18136 11777 18188
rect 11721 18134 11777 18136
rect 12004 18188 12060 18190
rect 12004 18136 12006 18188
rect 12006 18136 12058 18188
rect 12058 18136 12060 18188
rect 12004 18134 12060 18136
rect 11438 17970 11494 17972
rect 11438 17918 11440 17970
rect 11440 17918 11492 17970
rect 11492 17918 11494 17970
rect 11438 17916 11494 17918
rect 11721 17970 11777 17972
rect 11721 17918 11723 17970
rect 11723 17918 11775 17970
rect 11775 17918 11777 17970
rect 11721 17916 11777 17918
rect 12004 17970 12060 17972
rect 12004 17918 12006 17970
rect 12006 17918 12058 17970
rect 12058 17918 12060 17970
rect 12004 17916 12060 17918
rect 19005 20385 19061 20387
rect 19005 20333 19007 20385
rect 19007 20333 19059 20385
rect 19059 20333 19061 20385
rect 19005 20331 19061 20333
rect 19005 20167 19061 20169
rect 19005 20115 19007 20167
rect 19007 20115 19059 20167
rect 19059 20115 19061 20167
rect 19005 20113 19061 20115
rect 19005 19950 19061 19951
rect 19005 19898 19007 19950
rect 19007 19898 19059 19950
rect 19059 19898 19061 19950
rect 19005 19895 19061 19898
rect 17371 18426 17427 18428
rect 17371 18374 17373 18426
rect 17373 18374 17425 18426
rect 17425 18374 17427 18426
rect 17371 18372 17427 18374
rect 17371 18208 17427 18210
rect 17371 18156 17373 18208
rect 17373 18156 17425 18208
rect 17425 18156 17427 18208
rect 17371 18154 17427 18156
rect 17371 17991 17427 17992
rect 17371 17939 17373 17991
rect 17373 17939 17425 17991
rect 17425 17939 17427 17991
rect 17371 17936 17427 17939
rect 11438 17698 11494 17754
rect 11721 17698 11777 17754
rect 12004 17698 12060 17754
rect 17371 17773 17427 17774
rect 17371 17721 17373 17773
rect 17373 17721 17425 17773
rect 17425 17721 17427 17773
rect 17371 17718 17427 17721
rect 20638 20385 20694 20387
rect 20638 20333 20640 20385
rect 20640 20333 20692 20385
rect 20692 20333 20694 20385
rect 20638 20331 20694 20333
rect 20638 20167 20694 20169
rect 20638 20115 20640 20167
rect 20640 20115 20692 20167
rect 20692 20115 20694 20167
rect 20638 20113 20694 20115
rect 20638 19950 20694 19951
rect 20638 19898 20640 19950
rect 20640 19898 20692 19950
rect 20692 19898 20694 19950
rect 20638 19895 20694 19898
rect 19005 18426 19061 18428
rect 19005 18374 19007 18426
rect 19007 18374 19059 18426
rect 19059 18374 19061 18426
rect 19005 18372 19061 18374
rect 19005 18208 19061 18210
rect 19005 18156 19007 18208
rect 19007 18156 19059 18208
rect 19059 18156 19061 18208
rect 19005 18154 19061 18156
rect 19005 17991 19061 17992
rect 19005 17939 19007 17991
rect 19007 17939 19059 17991
rect 19059 17939 19061 17991
rect 19005 17936 19061 17939
rect 19005 17773 19061 17774
rect 19005 17721 19007 17773
rect 19007 17721 19059 17773
rect 19059 17721 19061 17773
rect 19005 17718 19061 17721
rect 22272 20385 22328 20387
rect 22272 20333 22274 20385
rect 22274 20333 22326 20385
rect 22326 20333 22328 20385
rect 22272 20331 22328 20333
rect 22272 20167 22328 20169
rect 22272 20115 22274 20167
rect 22274 20115 22326 20167
rect 22326 20115 22328 20167
rect 22272 20113 22328 20115
rect 22272 19950 22328 19951
rect 22272 19898 22274 19950
rect 22274 19898 22326 19950
rect 22326 19898 22328 19950
rect 22272 19895 22328 19898
rect 20638 18426 20694 18428
rect 20638 18374 20640 18426
rect 20640 18374 20692 18426
rect 20692 18374 20694 18426
rect 20638 18372 20694 18374
rect 20638 18208 20694 18210
rect 20638 18156 20640 18208
rect 20640 18156 20692 18208
rect 20692 18156 20694 18208
rect 20638 18154 20694 18156
rect 20638 17991 20694 17992
rect 20638 17939 20640 17991
rect 20640 17939 20692 17991
rect 20692 17939 20694 17991
rect 20638 17936 20694 17939
rect 20638 17773 20694 17774
rect 20638 17721 20640 17773
rect 20640 17721 20692 17773
rect 20692 17721 20694 17773
rect 20638 17718 20694 17721
rect 23957 24997 24013 24999
rect 23957 24945 23959 24997
rect 23959 24945 24011 24997
rect 24011 24945 24013 24997
rect 23957 24943 24013 24945
rect 23957 24780 24013 24782
rect 23957 24728 23959 24780
rect 23959 24728 24011 24780
rect 24011 24728 24013 24780
rect 23957 24726 24013 24728
rect 23957 24562 24013 24564
rect 23957 24510 23959 24562
rect 23959 24510 24011 24562
rect 24011 24510 24013 24562
rect 23957 24508 24013 24510
rect 23957 24344 24013 24346
rect 23957 24292 23959 24344
rect 23959 24292 24011 24344
rect 24011 24292 24013 24344
rect 23957 24290 24013 24292
rect 23957 24126 24013 24128
rect 23957 24074 23959 24126
rect 23959 24074 24011 24126
rect 24011 24074 24013 24126
rect 23957 24072 24013 24074
rect 23957 23909 24013 23911
rect 23957 23857 23959 23909
rect 23959 23857 24011 23909
rect 24011 23857 24013 23909
rect 23957 23855 24013 23857
rect 24471 24997 24527 24999
rect 24471 24945 24473 24997
rect 24473 24945 24525 24997
rect 24525 24945 24527 24997
rect 24471 24943 24527 24945
rect 24471 24780 24527 24782
rect 24471 24728 24473 24780
rect 24473 24728 24525 24780
rect 24525 24728 24527 24780
rect 24471 24726 24527 24728
rect 24471 24562 24527 24564
rect 24471 24510 24473 24562
rect 24473 24510 24525 24562
rect 24525 24510 24527 24562
rect 24471 24508 24527 24510
rect 24471 24344 24527 24346
rect 24471 24292 24473 24344
rect 24473 24292 24525 24344
rect 24525 24292 24527 24344
rect 24471 24290 24527 24292
rect 24471 24126 24527 24128
rect 24471 24074 24473 24126
rect 24473 24074 24525 24126
rect 24525 24074 24527 24126
rect 24471 24072 24527 24074
rect 24471 23909 24527 23911
rect 24471 23857 24473 23909
rect 24473 23857 24525 23909
rect 24525 23857 24527 23909
rect 24471 23855 24527 23857
rect 25427 26535 25483 26537
rect 25427 26483 25429 26535
rect 25429 26483 25481 26535
rect 25481 26483 25483 26535
rect 25427 26481 25483 26483
rect 25634 26535 25690 26537
rect 25634 26483 25636 26535
rect 25636 26483 25688 26535
rect 25688 26483 25690 26535
rect 25634 26481 25690 26483
rect 25427 26317 25483 26319
rect 25427 26265 25429 26317
rect 25429 26265 25481 26317
rect 25481 26265 25483 26317
rect 25427 26263 25483 26265
rect 25634 26317 25690 26319
rect 25634 26265 25636 26317
rect 25636 26265 25688 26317
rect 25688 26265 25690 26317
rect 25634 26263 25690 26265
rect 25427 26099 25483 26101
rect 25427 26047 25429 26099
rect 25429 26047 25481 26099
rect 25481 26047 25483 26099
rect 25427 26045 25483 26047
rect 25634 26099 25690 26101
rect 25634 26047 25636 26099
rect 25636 26047 25688 26099
rect 25688 26047 25690 26099
rect 25634 26045 25690 26047
rect 25427 25881 25483 25883
rect 25427 25829 25429 25881
rect 25429 25829 25481 25881
rect 25481 25829 25483 25881
rect 25427 25827 25483 25829
rect 25634 25881 25690 25883
rect 25634 25829 25636 25881
rect 25636 25829 25688 25881
rect 25688 25829 25690 25881
rect 25634 25827 25690 25829
rect 26154 26535 26210 26537
rect 26154 26483 26156 26535
rect 26156 26483 26208 26535
rect 26208 26483 26210 26535
rect 26154 26481 26210 26483
rect 26154 26317 26210 26319
rect 26154 26265 26156 26317
rect 26156 26265 26208 26317
rect 26208 26265 26210 26317
rect 26154 26263 26210 26265
rect 26154 26099 26210 26101
rect 26154 26047 26156 26099
rect 26156 26047 26208 26099
rect 26208 26047 26210 26099
rect 26154 26045 26210 26047
rect 26154 25881 26210 25883
rect 26154 25829 26156 25881
rect 26156 25829 26208 25881
rect 26208 25829 26210 25881
rect 26154 25827 26210 25829
rect 24950 22390 25006 22446
rect 24460 21914 24516 21970
rect 24460 21696 24516 21752
rect 24950 22172 25006 22228
rect 25647 24997 25703 24999
rect 25647 24945 25649 24997
rect 25649 24945 25701 24997
rect 25701 24945 25703 24997
rect 25647 24943 25703 24945
rect 25647 24780 25703 24782
rect 25647 24728 25649 24780
rect 25649 24728 25701 24780
rect 25701 24728 25703 24780
rect 25647 24726 25703 24728
rect 25647 24562 25703 24564
rect 25647 24510 25649 24562
rect 25649 24510 25701 24562
rect 25701 24510 25703 24562
rect 25647 24508 25703 24510
rect 25647 24344 25703 24346
rect 25647 24292 25649 24344
rect 25649 24292 25701 24344
rect 25701 24292 25703 24344
rect 25647 24290 25703 24292
rect 25647 24126 25703 24128
rect 25647 24074 25649 24126
rect 25649 24074 25701 24126
rect 25701 24074 25703 24126
rect 25647 24072 25703 24074
rect 25647 23909 25703 23911
rect 25647 23857 25649 23909
rect 25649 23857 25701 23909
rect 25701 23857 25703 23909
rect 25647 23855 25703 23857
rect 26161 24997 26217 24999
rect 26161 24945 26163 24997
rect 26163 24945 26215 24997
rect 26215 24945 26217 24997
rect 26161 24943 26217 24945
rect 26161 24780 26217 24782
rect 26161 24728 26163 24780
rect 26163 24728 26215 24780
rect 26215 24728 26217 24780
rect 26161 24726 26217 24728
rect 26161 24562 26217 24564
rect 26161 24510 26163 24562
rect 26163 24510 26215 24562
rect 26215 24510 26217 24562
rect 26161 24508 26217 24510
rect 26161 24344 26217 24346
rect 26161 24292 26163 24344
rect 26163 24292 26215 24344
rect 26215 24292 26217 24344
rect 26161 24290 26217 24292
rect 26161 24126 26217 24128
rect 26161 24074 26163 24126
rect 26163 24074 26215 24126
rect 26215 24074 26217 24126
rect 26161 24072 26217 24074
rect 26161 23909 26217 23911
rect 26161 23857 26163 23909
rect 26163 23857 26215 23909
rect 26215 23857 26217 23909
rect 26161 23855 26217 23857
rect 27118 26535 27174 26537
rect 27118 26483 27120 26535
rect 27120 26483 27172 26535
rect 27172 26483 27174 26535
rect 27118 26481 27174 26483
rect 27325 26535 27381 26537
rect 27325 26483 27327 26535
rect 27327 26483 27379 26535
rect 27379 26483 27381 26535
rect 27325 26481 27381 26483
rect 27118 26317 27174 26319
rect 27118 26265 27120 26317
rect 27120 26265 27172 26317
rect 27172 26265 27174 26317
rect 27118 26263 27174 26265
rect 27325 26317 27381 26319
rect 27325 26265 27327 26317
rect 27327 26265 27379 26317
rect 27379 26265 27381 26317
rect 27325 26263 27381 26265
rect 27118 26099 27174 26101
rect 27118 26047 27120 26099
rect 27120 26047 27172 26099
rect 27172 26047 27174 26099
rect 27118 26045 27174 26047
rect 27325 26099 27381 26101
rect 27325 26047 27327 26099
rect 27327 26047 27379 26099
rect 27379 26047 27381 26099
rect 27325 26045 27381 26047
rect 27118 25881 27174 25883
rect 27118 25829 27120 25881
rect 27120 25829 27172 25881
rect 27172 25829 27174 25881
rect 27118 25827 27174 25829
rect 27325 25881 27381 25883
rect 27325 25829 27327 25881
rect 27327 25829 27379 25881
rect 27379 25829 27381 25881
rect 27325 25827 27381 25829
rect 27845 26535 27901 26537
rect 27845 26483 27847 26535
rect 27847 26483 27899 26535
rect 27899 26483 27901 26535
rect 27845 26481 27901 26483
rect 27845 26317 27901 26319
rect 27845 26265 27847 26317
rect 27847 26265 27899 26317
rect 27899 26265 27901 26317
rect 27845 26263 27901 26265
rect 27845 26099 27901 26101
rect 27845 26047 27847 26099
rect 27847 26047 27899 26099
rect 27899 26047 27901 26099
rect 27845 26045 27901 26047
rect 27845 25881 27901 25883
rect 27845 25829 27847 25881
rect 27847 25829 27899 25881
rect 27899 25829 27901 25881
rect 27845 25827 27901 25829
rect 26640 22390 26696 22446
rect 26150 21914 26206 21970
rect 26150 21696 26206 21752
rect 26640 22172 26696 22228
rect 27338 24997 27394 24999
rect 27338 24945 27340 24997
rect 27340 24945 27392 24997
rect 27392 24945 27394 24997
rect 27338 24943 27394 24945
rect 27338 24780 27394 24782
rect 27338 24728 27340 24780
rect 27340 24728 27392 24780
rect 27392 24728 27394 24780
rect 27338 24726 27394 24728
rect 27338 24562 27394 24564
rect 27338 24510 27340 24562
rect 27340 24510 27392 24562
rect 27392 24510 27394 24562
rect 27338 24508 27394 24510
rect 27338 24344 27394 24346
rect 27338 24292 27340 24344
rect 27340 24292 27392 24344
rect 27392 24292 27394 24344
rect 27338 24290 27394 24292
rect 27338 24126 27394 24128
rect 27338 24074 27340 24126
rect 27340 24074 27392 24126
rect 27392 24074 27394 24126
rect 27338 24072 27394 24074
rect 27338 23909 27394 23911
rect 27338 23857 27340 23909
rect 27340 23857 27392 23909
rect 27392 23857 27394 23909
rect 27338 23855 27394 23857
rect 27852 24997 27908 24999
rect 27852 24945 27854 24997
rect 27854 24945 27906 24997
rect 27906 24945 27908 24997
rect 27852 24943 27908 24945
rect 27852 24780 27908 24782
rect 27852 24728 27854 24780
rect 27854 24728 27906 24780
rect 27906 24728 27908 24780
rect 27852 24726 27908 24728
rect 27852 24562 27908 24564
rect 27852 24510 27854 24562
rect 27854 24510 27906 24562
rect 27906 24510 27908 24562
rect 27852 24508 27908 24510
rect 27852 24344 27908 24346
rect 27852 24292 27854 24344
rect 27854 24292 27906 24344
rect 27906 24292 27908 24344
rect 27852 24290 27908 24292
rect 27852 24126 27908 24128
rect 27852 24074 27854 24126
rect 27854 24074 27906 24126
rect 27906 24074 27908 24126
rect 27852 24072 27908 24074
rect 27852 23909 27908 23911
rect 27852 23857 27854 23909
rect 27854 23857 27906 23909
rect 27906 23857 27908 23909
rect 27852 23855 27908 23857
rect 28331 22390 28387 22446
rect 28331 22172 28387 22228
rect 27841 21914 27897 21970
rect 27841 21696 27897 21752
rect 22272 18426 22328 18428
rect 22272 18374 22274 18426
rect 22274 18374 22326 18426
rect 22326 18374 22328 18426
rect 22272 18372 22328 18374
rect 22272 18208 22328 18210
rect 22272 18156 22274 18208
rect 22274 18156 22326 18208
rect 22326 18156 22328 18208
rect 22272 18154 22328 18156
rect 22272 17991 22328 17992
rect 22272 17939 22274 17991
rect 22274 17939 22326 17991
rect 22326 17939 22328 17991
rect 22272 17936 22328 17939
rect 22272 17773 22328 17774
rect 22272 17721 22274 17773
rect 22274 17721 22326 17773
rect 22326 17721 22328 17773
rect 22272 17718 22328 17721
rect 1990 16902 2046 16904
rect 1990 16850 1992 16902
rect 1992 16850 2044 16902
rect 2044 16850 2046 16902
rect 1990 16848 2046 16850
rect 1990 16778 2046 16780
rect 1990 16726 1992 16778
rect 1992 16726 2044 16778
rect 2044 16726 2046 16778
rect 1990 16724 2046 16726
rect 1990 16654 2046 16656
rect 1990 16602 1992 16654
rect 1992 16602 2044 16654
rect 2044 16602 2046 16654
rect 1990 16600 2046 16602
rect 1990 16530 2046 16532
rect 1990 16478 1992 16530
rect 1992 16478 2044 16530
rect 2044 16478 2046 16530
rect 1990 16476 2046 16478
rect 1990 16406 2046 16408
rect 1990 16354 1992 16406
rect 1992 16354 2044 16406
rect 2044 16354 2046 16406
rect 1990 16352 2046 16354
rect 1990 16282 2046 16284
rect 1990 16230 1992 16282
rect 1992 16230 2044 16282
rect 2044 16230 2046 16282
rect 1990 16228 2046 16230
rect 1990 16158 2046 16160
rect 1990 16106 1992 16158
rect 1992 16106 2044 16158
rect 2044 16106 2046 16158
rect 1990 16104 2046 16106
rect 1990 16034 2046 16036
rect 1990 15982 1992 16034
rect 1992 15982 2044 16034
rect 2044 15982 2046 16034
rect 1990 15980 2046 15982
rect 1990 15910 2046 15912
rect 1990 15858 1992 15910
rect 1992 15858 2044 15910
rect 2044 15858 2046 15910
rect 1990 15856 2046 15858
rect 1990 15786 2046 15788
rect 1990 15734 1992 15786
rect 1992 15734 2044 15786
rect 2044 15734 2046 15786
rect 1990 15732 2046 15734
rect 1990 15662 2046 15664
rect 1990 15610 1992 15662
rect 1992 15610 2044 15662
rect 2044 15610 2046 15662
rect 1990 15608 2046 15610
rect 1990 15538 2046 15540
rect 1990 15486 1992 15538
rect 1992 15486 2044 15538
rect 2044 15486 2046 15538
rect 1990 15484 2046 15486
rect 2662 16902 2718 16904
rect 2662 16850 2664 16902
rect 2664 16850 2716 16902
rect 2716 16850 2718 16902
rect 2662 16848 2718 16850
rect 2662 16778 2718 16780
rect 2662 16726 2664 16778
rect 2664 16726 2716 16778
rect 2716 16726 2718 16778
rect 2662 16724 2718 16726
rect 2662 16654 2718 16656
rect 2662 16602 2664 16654
rect 2664 16602 2716 16654
rect 2716 16602 2718 16654
rect 2662 16600 2718 16602
rect 2662 16530 2718 16532
rect 2662 16478 2664 16530
rect 2664 16478 2716 16530
rect 2716 16478 2718 16530
rect 2662 16476 2718 16478
rect 2662 16406 2718 16408
rect 2662 16354 2664 16406
rect 2664 16354 2716 16406
rect 2716 16354 2718 16406
rect 2662 16352 2718 16354
rect 2662 16282 2718 16284
rect 2662 16230 2664 16282
rect 2664 16230 2716 16282
rect 2716 16230 2718 16282
rect 2662 16228 2718 16230
rect 2662 16158 2718 16160
rect 2662 16106 2664 16158
rect 2664 16106 2716 16158
rect 2716 16106 2718 16158
rect 2662 16104 2718 16106
rect 2662 16034 2718 16036
rect 2662 15982 2664 16034
rect 2664 15982 2716 16034
rect 2716 15982 2718 16034
rect 2662 15980 2718 15982
rect 2662 15910 2718 15912
rect 2662 15858 2664 15910
rect 2664 15858 2716 15910
rect 2716 15858 2718 15910
rect 2662 15856 2718 15858
rect 2662 15786 2718 15788
rect 2662 15734 2664 15786
rect 2664 15734 2716 15786
rect 2716 15734 2718 15786
rect 2662 15732 2718 15734
rect 2662 15662 2718 15664
rect 2662 15610 2664 15662
rect 2664 15610 2716 15662
rect 2716 15610 2718 15662
rect 2662 15608 2718 15610
rect 2662 15538 2718 15540
rect 2662 15486 2664 15538
rect 2664 15486 2716 15538
rect 2716 15486 2718 15538
rect 2662 15484 2718 15486
rect 3110 16902 3166 16904
rect 3110 16850 3112 16902
rect 3112 16850 3164 16902
rect 3164 16850 3166 16902
rect 3110 16848 3166 16850
rect 3110 16778 3166 16780
rect 3110 16726 3112 16778
rect 3112 16726 3164 16778
rect 3164 16726 3166 16778
rect 3110 16724 3166 16726
rect 3110 16654 3166 16656
rect 3110 16602 3112 16654
rect 3112 16602 3164 16654
rect 3164 16602 3166 16654
rect 3110 16600 3166 16602
rect 3110 16530 3166 16532
rect 3110 16478 3112 16530
rect 3112 16478 3164 16530
rect 3164 16478 3166 16530
rect 3110 16476 3166 16478
rect 3110 16406 3166 16408
rect 3110 16354 3112 16406
rect 3112 16354 3164 16406
rect 3164 16354 3166 16406
rect 3110 16352 3166 16354
rect 3110 16282 3166 16284
rect 3110 16230 3112 16282
rect 3112 16230 3164 16282
rect 3164 16230 3166 16282
rect 3110 16228 3166 16230
rect 3110 16158 3166 16160
rect 3110 16106 3112 16158
rect 3112 16106 3164 16158
rect 3164 16106 3166 16158
rect 3110 16104 3166 16106
rect 3110 16034 3166 16036
rect 3110 15982 3112 16034
rect 3112 15982 3164 16034
rect 3164 15982 3166 16034
rect 3110 15980 3166 15982
rect 3110 15910 3166 15912
rect 3110 15858 3112 15910
rect 3112 15858 3164 15910
rect 3164 15858 3166 15910
rect 3110 15856 3166 15858
rect 3110 15786 3166 15788
rect 3110 15734 3112 15786
rect 3112 15734 3164 15786
rect 3164 15734 3166 15786
rect 3110 15732 3166 15734
rect 3110 15662 3166 15664
rect 3110 15610 3112 15662
rect 3112 15610 3164 15662
rect 3164 15610 3166 15662
rect 3110 15608 3166 15610
rect 3110 15538 3166 15540
rect 3110 15486 3112 15538
rect 3112 15486 3164 15538
rect 3164 15486 3166 15538
rect 3110 15484 3166 15486
rect 3782 16902 3838 16904
rect 3782 16850 3784 16902
rect 3784 16850 3836 16902
rect 3836 16850 3838 16902
rect 3782 16848 3838 16850
rect 3782 16778 3838 16780
rect 3782 16726 3784 16778
rect 3784 16726 3836 16778
rect 3836 16726 3838 16778
rect 3782 16724 3838 16726
rect 3782 16654 3838 16656
rect 3782 16602 3784 16654
rect 3784 16602 3836 16654
rect 3836 16602 3838 16654
rect 3782 16600 3838 16602
rect 3782 16530 3838 16532
rect 3782 16478 3784 16530
rect 3784 16478 3836 16530
rect 3836 16478 3838 16530
rect 3782 16476 3838 16478
rect 3782 16406 3838 16408
rect 3782 16354 3784 16406
rect 3784 16354 3836 16406
rect 3836 16354 3838 16406
rect 3782 16352 3838 16354
rect 3782 16282 3838 16284
rect 3782 16230 3784 16282
rect 3784 16230 3836 16282
rect 3836 16230 3838 16282
rect 3782 16228 3838 16230
rect 3782 16158 3838 16160
rect 3782 16106 3784 16158
rect 3784 16106 3836 16158
rect 3836 16106 3838 16158
rect 3782 16104 3838 16106
rect 3782 16034 3838 16036
rect 3782 15982 3784 16034
rect 3784 15982 3836 16034
rect 3836 15982 3838 16034
rect 3782 15980 3838 15982
rect 3782 15910 3838 15912
rect 3782 15858 3784 15910
rect 3784 15858 3836 15910
rect 3836 15858 3838 15910
rect 3782 15856 3838 15858
rect 3782 15786 3838 15788
rect 3782 15734 3784 15786
rect 3784 15734 3836 15786
rect 3836 15734 3838 15786
rect 3782 15732 3838 15734
rect 3782 15662 3838 15664
rect 3782 15610 3784 15662
rect 3784 15610 3836 15662
rect 3836 15610 3838 15662
rect 3782 15608 3838 15610
rect 3782 15538 3838 15540
rect 3782 15486 3784 15538
rect 3784 15486 3836 15538
rect 3836 15486 3838 15538
rect 3782 15484 3838 15486
rect 4230 16902 4286 16904
rect 4230 16850 4232 16902
rect 4232 16850 4284 16902
rect 4284 16850 4286 16902
rect 4230 16848 4286 16850
rect 4230 16778 4286 16780
rect 4230 16726 4232 16778
rect 4232 16726 4284 16778
rect 4284 16726 4286 16778
rect 4230 16724 4286 16726
rect 4230 16654 4286 16656
rect 4230 16602 4232 16654
rect 4232 16602 4284 16654
rect 4284 16602 4286 16654
rect 4230 16600 4286 16602
rect 4230 16530 4286 16532
rect 4230 16478 4232 16530
rect 4232 16478 4284 16530
rect 4284 16478 4286 16530
rect 4230 16476 4286 16478
rect 4230 16406 4286 16408
rect 4230 16354 4232 16406
rect 4232 16354 4284 16406
rect 4284 16354 4286 16406
rect 4230 16352 4286 16354
rect 4230 16282 4286 16284
rect 4230 16230 4232 16282
rect 4232 16230 4284 16282
rect 4284 16230 4286 16282
rect 4230 16228 4286 16230
rect 4230 16158 4286 16160
rect 4230 16106 4232 16158
rect 4232 16106 4284 16158
rect 4284 16106 4286 16158
rect 4230 16104 4286 16106
rect 4230 16034 4286 16036
rect 4230 15982 4232 16034
rect 4232 15982 4284 16034
rect 4284 15982 4286 16034
rect 4230 15980 4286 15982
rect 4230 15910 4286 15912
rect 4230 15858 4232 15910
rect 4232 15858 4284 15910
rect 4284 15858 4286 15910
rect 4230 15856 4286 15858
rect 4230 15786 4286 15788
rect 4230 15734 4232 15786
rect 4232 15734 4284 15786
rect 4284 15734 4286 15786
rect 4230 15732 4286 15734
rect 4230 15662 4286 15664
rect 4230 15610 4232 15662
rect 4232 15610 4284 15662
rect 4284 15610 4286 15662
rect 4230 15608 4286 15610
rect 4230 15538 4286 15540
rect 4230 15486 4232 15538
rect 4232 15486 4284 15538
rect 4284 15486 4286 15538
rect 4230 15484 4286 15486
rect 4902 16902 4958 16904
rect 4902 16850 4904 16902
rect 4904 16850 4956 16902
rect 4956 16850 4958 16902
rect 4902 16848 4958 16850
rect 4902 16778 4958 16780
rect 4902 16726 4904 16778
rect 4904 16726 4956 16778
rect 4956 16726 4958 16778
rect 4902 16724 4958 16726
rect 4902 16654 4958 16656
rect 4902 16602 4904 16654
rect 4904 16602 4956 16654
rect 4956 16602 4958 16654
rect 4902 16600 4958 16602
rect 4902 16530 4958 16532
rect 4902 16478 4904 16530
rect 4904 16478 4956 16530
rect 4956 16478 4958 16530
rect 4902 16476 4958 16478
rect 4902 16406 4958 16408
rect 4902 16354 4904 16406
rect 4904 16354 4956 16406
rect 4956 16354 4958 16406
rect 4902 16352 4958 16354
rect 4902 16282 4958 16284
rect 4902 16230 4904 16282
rect 4904 16230 4956 16282
rect 4956 16230 4958 16282
rect 4902 16228 4958 16230
rect 4902 16158 4958 16160
rect 4902 16106 4904 16158
rect 4904 16106 4956 16158
rect 4956 16106 4958 16158
rect 4902 16104 4958 16106
rect 4902 16034 4958 16036
rect 4902 15982 4904 16034
rect 4904 15982 4956 16034
rect 4956 15982 4958 16034
rect 4902 15980 4958 15982
rect 4902 15910 4958 15912
rect 4902 15858 4904 15910
rect 4904 15858 4956 15910
rect 4956 15858 4958 15910
rect 4902 15856 4958 15858
rect 4902 15786 4958 15788
rect 4902 15734 4904 15786
rect 4904 15734 4956 15786
rect 4956 15734 4958 15786
rect 4902 15732 4958 15734
rect 4902 15662 4958 15664
rect 4902 15610 4904 15662
rect 4904 15610 4956 15662
rect 4956 15610 4958 15662
rect 4902 15608 4958 15610
rect 4902 15538 4958 15540
rect 4902 15486 4904 15538
rect 4904 15486 4956 15538
rect 4956 15486 4958 15538
rect 4902 15484 4958 15486
rect 5350 16902 5406 16904
rect 5350 16850 5352 16902
rect 5352 16850 5404 16902
rect 5404 16850 5406 16902
rect 5350 16848 5406 16850
rect 5350 16778 5406 16780
rect 5350 16726 5352 16778
rect 5352 16726 5404 16778
rect 5404 16726 5406 16778
rect 5350 16724 5406 16726
rect 5350 16654 5406 16656
rect 5350 16602 5352 16654
rect 5352 16602 5404 16654
rect 5404 16602 5406 16654
rect 5350 16600 5406 16602
rect 5350 16530 5406 16532
rect 5350 16478 5352 16530
rect 5352 16478 5404 16530
rect 5404 16478 5406 16530
rect 5350 16476 5406 16478
rect 5350 16406 5406 16408
rect 5350 16354 5352 16406
rect 5352 16354 5404 16406
rect 5404 16354 5406 16406
rect 5350 16352 5406 16354
rect 5350 16282 5406 16284
rect 5350 16230 5352 16282
rect 5352 16230 5404 16282
rect 5404 16230 5406 16282
rect 5350 16228 5406 16230
rect 5350 16158 5406 16160
rect 5350 16106 5352 16158
rect 5352 16106 5404 16158
rect 5404 16106 5406 16158
rect 5350 16104 5406 16106
rect 5350 16034 5406 16036
rect 5350 15982 5352 16034
rect 5352 15982 5404 16034
rect 5404 15982 5406 16034
rect 5350 15980 5406 15982
rect 5350 15910 5406 15912
rect 5350 15858 5352 15910
rect 5352 15858 5404 15910
rect 5404 15858 5406 15910
rect 5350 15856 5406 15858
rect 5350 15786 5406 15788
rect 5350 15734 5352 15786
rect 5352 15734 5404 15786
rect 5404 15734 5406 15786
rect 5350 15732 5406 15734
rect 5350 15662 5406 15664
rect 5350 15610 5352 15662
rect 5352 15610 5404 15662
rect 5404 15610 5406 15662
rect 5350 15608 5406 15610
rect 5350 15538 5406 15540
rect 5350 15486 5352 15538
rect 5352 15486 5404 15538
rect 5404 15486 5406 15538
rect 5350 15484 5406 15486
rect 6022 16902 6078 16904
rect 6022 16850 6024 16902
rect 6024 16850 6076 16902
rect 6076 16850 6078 16902
rect 6022 16848 6078 16850
rect 6022 16778 6078 16780
rect 6022 16726 6024 16778
rect 6024 16726 6076 16778
rect 6076 16726 6078 16778
rect 6022 16724 6078 16726
rect 6022 16654 6078 16656
rect 6022 16602 6024 16654
rect 6024 16602 6076 16654
rect 6076 16602 6078 16654
rect 6022 16600 6078 16602
rect 6022 16530 6078 16532
rect 6022 16478 6024 16530
rect 6024 16478 6076 16530
rect 6076 16478 6078 16530
rect 6022 16476 6078 16478
rect 6022 16406 6078 16408
rect 6022 16354 6024 16406
rect 6024 16354 6076 16406
rect 6076 16354 6078 16406
rect 6022 16352 6078 16354
rect 6022 16282 6078 16284
rect 6022 16230 6024 16282
rect 6024 16230 6076 16282
rect 6076 16230 6078 16282
rect 6022 16228 6078 16230
rect 6022 16158 6078 16160
rect 6022 16106 6024 16158
rect 6024 16106 6076 16158
rect 6076 16106 6078 16158
rect 6022 16104 6078 16106
rect 6022 16034 6078 16036
rect 6022 15982 6024 16034
rect 6024 15982 6076 16034
rect 6076 15982 6078 16034
rect 6022 15980 6078 15982
rect 6022 15910 6078 15912
rect 6022 15858 6024 15910
rect 6024 15858 6076 15910
rect 6076 15858 6078 15910
rect 6022 15856 6078 15858
rect 6022 15786 6078 15788
rect 6022 15734 6024 15786
rect 6024 15734 6076 15786
rect 6076 15734 6078 15786
rect 6022 15732 6078 15734
rect 6022 15662 6078 15664
rect 6022 15610 6024 15662
rect 6024 15610 6076 15662
rect 6076 15610 6078 15662
rect 6022 15608 6078 15610
rect 6022 15538 6078 15540
rect 6022 15486 6024 15538
rect 6024 15486 6076 15538
rect 6076 15486 6078 15538
rect 6022 15484 6078 15486
rect 6470 16902 6526 16904
rect 6470 16850 6472 16902
rect 6472 16850 6524 16902
rect 6524 16850 6526 16902
rect 6470 16848 6526 16850
rect 6470 16778 6526 16780
rect 6470 16726 6472 16778
rect 6472 16726 6524 16778
rect 6524 16726 6526 16778
rect 6470 16724 6526 16726
rect 6470 16654 6526 16656
rect 6470 16602 6472 16654
rect 6472 16602 6524 16654
rect 6524 16602 6526 16654
rect 6470 16600 6526 16602
rect 6470 16530 6526 16532
rect 6470 16478 6472 16530
rect 6472 16478 6524 16530
rect 6524 16478 6526 16530
rect 6470 16476 6526 16478
rect 6470 16406 6526 16408
rect 6470 16354 6472 16406
rect 6472 16354 6524 16406
rect 6524 16354 6526 16406
rect 6470 16352 6526 16354
rect 6470 16282 6526 16284
rect 6470 16230 6472 16282
rect 6472 16230 6524 16282
rect 6524 16230 6526 16282
rect 6470 16228 6526 16230
rect 6470 16158 6526 16160
rect 6470 16106 6472 16158
rect 6472 16106 6524 16158
rect 6524 16106 6526 16158
rect 6470 16104 6526 16106
rect 6470 16034 6526 16036
rect 6470 15982 6472 16034
rect 6472 15982 6524 16034
rect 6524 15982 6526 16034
rect 6470 15980 6526 15982
rect 6470 15910 6526 15912
rect 6470 15858 6472 15910
rect 6472 15858 6524 15910
rect 6524 15858 6526 15910
rect 6470 15856 6526 15858
rect 6470 15786 6526 15788
rect 6470 15734 6472 15786
rect 6472 15734 6524 15786
rect 6524 15734 6526 15786
rect 6470 15732 6526 15734
rect 6470 15662 6526 15664
rect 6470 15610 6472 15662
rect 6472 15610 6524 15662
rect 6524 15610 6526 15662
rect 6470 15608 6526 15610
rect 6470 15538 6526 15540
rect 6470 15486 6472 15538
rect 6472 15486 6524 15538
rect 6524 15486 6526 15538
rect 6470 15484 6526 15486
rect 7142 16902 7198 16904
rect 7142 16850 7144 16902
rect 7144 16850 7196 16902
rect 7196 16850 7198 16902
rect 7142 16848 7198 16850
rect 7142 16778 7198 16780
rect 7142 16726 7144 16778
rect 7144 16726 7196 16778
rect 7196 16726 7198 16778
rect 7142 16724 7198 16726
rect 7142 16654 7198 16656
rect 7142 16602 7144 16654
rect 7144 16602 7196 16654
rect 7196 16602 7198 16654
rect 7142 16600 7198 16602
rect 7142 16530 7198 16532
rect 7142 16478 7144 16530
rect 7144 16478 7196 16530
rect 7196 16478 7198 16530
rect 7142 16476 7198 16478
rect 7142 16406 7198 16408
rect 7142 16354 7144 16406
rect 7144 16354 7196 16406
rect 7196 16354 7198 16406
rect 7142 16352 7198 16354
rect 7142 16282 7198 16284
rect 7142 16230 7144 16282
rect 7144 16230 7196 16282
rect 7196 16230 7198 16282
rect 7142 16228 7198 16230
rect 7142 16158 7198 16160
rect 7142 16106 7144 16158
rect 7144 16106 7196 16158
rect 7196 16106 7198 16158
rect 7142 16104 7198 16106
rect 7142 16034 7198 16036
rect 7142 15982 7144 16034
rect 7144 15982 7196 16034
rect 7196 15982 7198 16034
rect 7142 15980 7198 15982
rect 7142 15910 7198 15912
rect 7142 15858 7144 15910
rect 7144 15858 7196 15910
rect 7196 15858 7198 15910
rect 7142 15856 7198 15858
rect 7142 15786 7198 15788
rect 7142 15734 7144 15786
rect 7144 15734 7196 15786
rect 7196 15734 7198 15786
rect 7142 15732 7198 15734
rect 7142 15662 7198 15664
rect 7142 15610 7144 15662
rect 7144 15610 7196 15662
rect 7196 15610 7198 15662
rect 7142 15608 7198 15610
rect 7142 15538 7198 15540
rect 7142 15486 7144 15538
rect 7144 15486 7196 15538
rect 7196 15486 7198 15538
rect 7142 15484 7198 15486
rect 7590 16902 7646 16904
rect 7590 16850 7592 16902
rect 7592 16850 7644 16902
rect 7644 16850 7646 16902
rect 7590 16848 7646 16850
rect 7590 16778 7646 16780
rect 7590 16726 7592 16778
rect 7592 16726 7644 16778
rect 7644 16726 7646 16778
rect 7590 16724 7646 16726
rect 7590 16654 7646 16656
rect 7590 16602 7592 16654
rect 7592 16602 7644 16654
rect 7644 16602 7646 16654
rect 7590 16600 7646 16602
rect 7590 16530 7646 16532
rect 7590 16478 7592 16530
rect 7592 16478 7644 16530
rect 7644 16478 7646 16530
rect 7590 16476 7646 16478
rect 7590 16406 7646 16408
rect 7590 16354 7592 16406
rect 7592 16354 7644 16406
rect 7644 16354 7646 16406
rect 7590 16352 7646 16354
rect 7590 16282 7646 16284
rect 7590 16230 7592 16282
rect 7592 16230 7644 16282
rect 7644 16230 7646 16282
rect 7590 16228 7646 16230
rect 7590 16158 7646 16160
rect 7590 16106 7592 16158
rect 7592 16106 7644 16158
rect 7644 16106 7646 16158
rect 7590 16104 7646 16106
rect 7590 16034 7646 16036
rect 7590 15982 7592 16034
rect 7592 15982 7644 16034
rect 7644 15982 7646 16034
rect 7590 15980 7646 15982
rect 7590 15910 7646 15912
rect 7590 15858 7592 15910
rect 7592 15858 7644 15910
rect 7644 15858 7646 15910
rect 7590 15856 7646 15858
rect 7590 15786 7646 15788
rect 7590 15734 7592 15786
rect 7592 15734 7644 15786
rect 7644 15734 7646 15786
rect 7590 15732 7646 15734
rect 7590 15662 7646 15664
rect 7590 15610 7592 15662
rect 7592 15610 7644 15662
rect 7644 15610 7646 15662
rect 7590 15608 7646 15610
rect 7590 15538 7646 15540
rect 7590 15486 7592 15538
rect 7592 15486 7644 15538
rect 7644 15486 7646 15538
rect 7590 15484 7646 15486
rect 8262 16902 8318 16904
rect 8262 16850 8264 16902
rect 8264 16850 8316 16902
rect 8316 16850 8318 16902
rect 8262 16848 8318 16850
rect 8262 16778 8318 16780
rect 8262 16726 8264 16778
rect 8264 16726 8316 16778
rect 8316 16726 8318 16778
rect 8262 16724 8318 16726
rect 8262 16654 8318 16656
rect 8262 16602 8264 16654
rect 8264 16602 8316 16654
rect 8316 16602 8318 16654
rect 8262 16600 8318 16602
rect 8262 16530 8318 16532
rect 8262 16478 8264 16530
rect 8264 16478 8316 16530
rect 8316 16478 8318 16530
rect 8262 16476 8318 16478
rect 8262 16406 8318 16408
rect 8262 16354 8264 16406
rect 8264 16354 8316 16406
rect 8316 16354 8318 16406
rect 8262 16352 8318 16354
rect 8262 16282 8318 16284
rect 8262 16230 8264 16282
rect 8264 16230 8316 16282
rect 8316 16230 8318 16282
rect 8262 16228 8318 16230
rect 8262 16158 8318 16160
rect 8262 16106 8264 16158
rect 8264 16106 8316 16158
rect 8316 16106 8318 16158
rect 8262 16104 8318 16106
rect 8262 16034 8318 16036
rect 8262 15982 8264 16034
rect 8264 15982 8316 16034
rect 8316 15982 8318 16034
rect 8262 15980 8318 15982
rect 8262 15910 8318 15912
rect 8262 15858 8264 15910
rect 8264 15858 8316 15910
rect 8316 15858 8318 15910
rect 8262 15856 8318 15858
rect 8262 15786 8318 15788
rect 8262 15734 8264 15786
rect 8264 15734 8316 15786
rect 8316 15734 8318 15786
rect 8262 15732 8318 15734
rect 8262 15662 8318 15664
rect 8262 15610 8264 15662
rect 8264 15610 8316 15662
rect 8316 15610 8318 15662
rect 8262 15608 8318 15610
rect 8262 15538 8318 15540
rect 8262 15486 8264 15538
rect 8264 15486 8316 15538
rect 8316 15486 8318 15538
rect 8262 15484 8318 15486
rect 8710 16902 8766 16904
rect 8710 16850 8712 16902
rect 8712 16850 8764 16902
rect 8764 16850 8766 16902
rect 8710 16848 8766 16850
rect 8710 16778 8766 16780
rect 8710 16726 8712 16778
rect 8712 16726 8764 16778
rect 8764 16726 8766 16778
rect 8710 16724 8766 16726
rect 8710 16654 8766 16656
rect 8710 16602 8712 16654
rect 8712 16602 8764 16654
rect 8764 16602 8766 16654
rect 8710 16600 8766 16602
rect 8710 16530 8766 16532
rect 8710 16478 8712 16530
rect 8712 16478 8764 16530
rect 8764 16478 8766 16530
rect 8710 16476 8766 16478
rect 8710 16406 8766 16408
rect 8710 16354 8712 16406
rect 8712 16354 8764 16406
rect 8764 16354 8766 16406
rect 8710 16352 8766 16354
rect 8710 16282 8766 16284
rect 8710 16230 8712 16282
rect 8712 16230 8764 16282
rect 8764 16230 8766 16282
rect 8710 16228 8766 16230
rect 8710 16158 8766 16160
rect 8710 16106 8712 16158
rect 8712 16106 8764 16158
rect 8764 16106 8766 16158
rect 8710 16104 8766 16106
rect 8710 16034 8766 16036
rect 8710 15982 8712 16034
rect 8712 15982 8764 16034
rect 8764 15982 8766 16034
rect 8710 15980 8766 15982
rect 8710 15910 8766 15912
rect 8710 15858 8712 15910
rect 8712 15858 8764 15910
rect 8764 15858 8766 15910
rect 8710 15856 8766 15858
rect 8710 15786 8766 15788
rect 8710 15734 8712 15786
rect 8712 15734 8764 15786
rect 8764 15734 8766 15786
rect 8710 15732 8766 15734
rect 8710 15662 8766 15664
rect 8710 15610 8712 15662
rect 8712 15610 8764 15662
rect 8764 15610 8766 15662
rect 8710 15608 8766 15610
rect 8710 15538 8766 15540
rect 8710 15486 8712 15538
rect 8712 15486 8764 15538
rect 8764 15486 8766 15538
rect 8710 15484 8766 15486
rect 9382 16902 9438 16904
rect 9382 16850 9384 16902
rect 9384 16850 9436 16902
rect 9436 16850 9438 16902
rect 9382 16848 9438 16850
rect 9382 16778 9438 16780
rect 9382 16726 9384 16778
rect 9384 16726 9436 16778
rect 9436 16726 9438 16778
rect 9382 16724 9438 16726
rect 9382 16654 9438 16656
rect 9382 16602 9384 16654
rect 9384 16602 9436 16654
rect 9436 16602 9438 16654
rect 9382 16600 9438 16602
rect 9382 16530 9438 16532
rect 9382 16478 9384 16530
rect 9384 16478 9436 16530
rect 9436 16478 9438 16530
rect 9382 16476 9438 16478
rect 9382 16406 9438 16408
rect 9382 16354 9384 16406
rect 9384 16354 9436 16406
rect 9436 16354 9438 16406
rect 9382 16352 9438 16354
rect 9382 16282 9438 16284
rect 9382 16230 9384 16282
rect 9384 16230 9436 16282
rect 9436 16230 9438 16282
rect 9382 16228 9438 16230
rect 9382 16158 9438 16160
rect 9382 16106 9384 16158
rect 9384 16106 9436 16158
rect 9436 16106 9438 16158
rect 9382 16104 9438 16106
rect 9382 16034 9438 16036
rect 9382 15982 9384 16034
rect 9384 15982 9436 16034
rect 9436 15982 9438 16034
rect 9382 15980 9438 15982
rect 9382 15910 9438 15912
rect 9382 15858 9384 15910
rect 9384 15858 9436 15910
rect 9436 15858 9438 15910
rect 9382 15856 9438 15858
rect 9382 15786 9438 15788
rect 9382 15734 9384 15786
rect 9384 15734 9436 15786
rect 9436 15734 9438 15786
rect 9382 15732 9438 15734
rect 9382 15662 9438 15664
rect 9382 15610 9384 15662
rect 9384 15610 9436 15662
rect 9436 15610 9438 15662
rect 9382 15608 9438 15610
rect 9382 15538 9438 15540
rect 9382 15486 9384 15538
rect 9384 15486 9436 15538
rect 9436 15486 9438 15538
rect 9382 15484 9438 15486
rect 9830 16902 9886 16904
rect 9830 16850 9832 16902
rect 9832 16850 9884 16902
rect 9884 16850 9886 16902
rect 9830 16848 9886 16850
rect 9830 16778 9886 16780
rect 9830 16726 9832 16778
rect 9832 16726 9884 16778
rect 9884 16726 9886 16778
rect 9830 16724 9886 16726
rect 9830 16654 9886 16656
rect 9830 16602 9832 16654
rect 9832 16602 9884 16654
rect 9884 16602 9886 16654
rect 9830 16600 9886 16602
rect 9830 16530 9886 16532
rect 9830 16478 9832 16530
rect 9832 16478 9884 16530
rect 9884 16478 9886 16530
rect 9830 16476 9886 16478
rect 9830 16406 9886 16408
rect 9830 16354 9832 16406
rect 9832 16354 9884 16406
rect 9884 16354 9886 16406
rect 9830 16352 9886 16354
rect 9830 16282 9886 16284
rect 9830 16230 9832 16282
rect 9832 16230 9884 16282
rect 9884 16230 9886 16282
rect 9830 16228 9886 16230
rect 9830 16158 9886 16160
rect 9830 16106 9832 16158
rect 9832 16106 9884 16158
rect 9884 16106 9886 16158
rect 9830 16104 9886 16106
rect 9830 16034 9886 16036
rect 9830 15982 9832 16034
rect 9832 15982 9884 16034
rect 9884 15982 9886 16034
rect 9830 15980 9886 15982
rect 9830 15910 9886 15912
rect 9830 15858 9832 15910
rect 9832 15858 9884 15910
rect 9884 15858 9886 15910
rect 9830 15856 9886 15858
rect 9830 15786 9886 15788
rect 9830 15734 9832 15786
rect 9832 15734 9884 15786
rect 9884 15734 9886 15786
rect 9830 15732 9886 15734
rect 9830 15662 9886 15664
rect 9830 15610 9832 15662
rect 9832 15610 9884 15662
rect 9884 15610 9886 15662
rect 9830 15608 9886 15610
rect 9830 15538 9886 15540
rect 9830 15486 9832 15538
rect 9832 15486 9884 15538
rect 9884 15486 9886 15538
rect 9830 15484 9886 15486
rect 10502 16902 10558 16904
rect 10502 16850 10504 16902
rect 10504 16850 10556 16902
rect 10556 16850 10558 16902
rect 10502 16848 10558 16850
rect 10502 16778 10558 16780
rect 10502 16726 10504 16778
rect 10504 16726 10556 16778
rect 10556 16726 10558 16778
rect 10502 16724 10558 16726
rect 10502 16654 10558 16656
rect 10502 16602 10504 16654
rect 10504 16602 10556 16654
rect 10556 16602 10558 16654
rect 10502 16600 10558 16602
rect 10502 16530 10558 16532
rect 10502 16478 10504 16530
rect 10504 16478 10556 16530
rect 10556 16478 10558 16530
rect 10502 16476 10558 16478
rect 10502 16406 10558 16408
rect 10502 16354 10504 16406
rect 10504 16354 10556 16406
rect 10556 16354 10558 16406
rect 10502 16352 10558 16354
rect 10502 16282 10558 16284
rect 10502 16230 10504 16282
rect 10504 16230 10556 16282
rect 10556 16230 10558 16282
rect 10502 16228 10558 16230
rect 10502 16158 10558 16160
rect 10502 16106 10504 16158
rect 10504 16106 10556 16158
rect 10556 16106 10558 16158
rect 10502 16104 10558 16106
rect 10502 16034 10558 16036
rect 10502 15982 10504 16034
rect 10504 15982 10556 16034
rect 10556 15982 10558 16034
rect 10502 15980 10558 15982
rect 10502 15910 10558 15912
rect 10502 15858 10504 15910
rect 10504 15858 10556 15910
rect 10556 15858 10558 15910
rect 10502 15856 10558 15858
rect 10502 15786 10558 15788
rect 10502 15734 10504 15786
rect 10504 15734 10556 15786
rect 10556 15734 10558 15786
rect 10502 15732 10558 15734
rect 10502 15662 10558 15664
rect 10502 15610 10504 15662
rect 10504 15610 10556 15662
rect 10556 15610 10558 15662
rect 10502 15608 10558 15610
rect 10502 15538 10558 15540
rect 10502 15486 10504 15538
rect 10504 15486 10556 15538
rect 10556 15486 10558 15538
rect 10502 15484 10558 15486
rect 10950 16902 11006 16904
rect 10950 16850 10952 16902
rect 10952 16850 11004 16902
rect 11004 16850 11006 16902
rect 10950 16848 11006 16850
rect 10950 16778 11006 16780
rect 10950 16726 10952 16778
rect 10952 16726 11004 16778
rect 11004 16726 11006 16778
rect 10950 16724 11006 16726
rect 10950 16654 11006 16656
rect 10950 16602 10952 16654
rect 10952 16602 11004 16654
rect 11004 16602 11006 16654
rect 10950 16600 11006 16602
rect 10950 16530 11006 16532
rect 10950 16478 10952 16530
rect 10952 16478 11004 16530
rect 11004 16478 11006 16530
rect 10950 16476 11006 16478
rect 10950 16406 11006 16408
rect 10950 16354 10952 16406
rect 10952 16354 11004 16406
rect 11004 16354 11006 16406
rect 10950 16352 11006 16354
rect 10950 16282 11006 16284
rect 10950 16230 10952 16282
rect 10952 16230 11004 16282
rect 11004 16230 11006 16282
rect 10950 16228 11006 16230
rect 10950 16158 11006 16160
rect 10950 16106 10952 16158
rect 10952 16106 11004 16158
rect 11004 16106 11006 16158
rect 10950 16104 11006 16106
rect 10950 16034 11006 16036
rect 10950 15982 10952 16034
rect 10952 15982 11004 16034
rect 11004 15982 11006 16034
rect 10950 15980 11006 15982
rect 10950 15910 11006 15912
rect 10950 15858 10952 15910
rect 10952 15858 11004 15910
rect 11004 15858 11006 15910
rect 10950 15856 11006 15858
rect 10950 15786 11006 15788
rect 10950 15734 10952 15786
rect 10952 15734 11004 15786
rect 11004 15734 11006 15786
rect 10950 15732 11006 15734
rect 10950 15662 11006 15664
rect 10950 15610 10952 15662
rect 10952 15610 11004 15662
rect 11004 15610 11006 15662
rect 10950 15608 11006 15610
rect 10950 15538 11006 15540
rect 10950 15486 10952 15538
rect 10952 15486 11004 15538
rect 11004 15486 11006 15538
rect 10950 15484 11006 15486
rect 11622 16902 11678 16904
rect 11622 16850 11624 16902
rect 11624 16850 11676 16902
rect 11676 16850 11678 16902
rect 11622 16848 11678 16850
rect 11622 16778 11678 16780
rect 11622 16726 11624 16778
rect 11624 16726 11676 16778
rect 11676 16726 11678 16778
rect 11622 16724 11678 16726
rect 11622 16654 11678 16656
rect 11622 16602 11624 16654
rect 11624 16602 11676 16654
rect 11676 16602 11678 16654
rect 11622 16600 11678 16602
rect 11622 16530 11678 16532
rect 11622 16478 11624 16530
rect 11624 16478 11676 16530
rect 11676 16478 11678 16530
rect 11622 16476 11678 16478
rect 11622 16406 11678 16408
rect 11622 16354 11624 16406
rect 11624 16354 11676 16406
rect 11676 16354 11678 16406
rect 11622 16352 11678 16354
rect 11622 16282 11678 16284
rect 11622 16230 11624 16282
rect 11624 16230 11676 16282
rect 11676 16230 11678 16282
rect 11622 16228 11678 16230
rect 11622 16158 11678 16160
rect 11622 16106 11624 16158
rect 11624 16106 11676 16158
rect 11676 16106 11678 16158
rect 11622 16104 11678 16106
rect 11622 16034 11678 16036
rect 11622 15982 11624 16034
rect 11624 15982 11676 16034
rect 11676 15982 11678 16034
rect 11622 15980 11678 15982
rect 11622 15910 11678 15912
rect 11622 15858 11624 15910
rect 11624 15858 11676 15910
rect 11676 15858 11678 15910
rect 11622 15856 11678 15858
rect 11622 15786 11678 15788
rect 11622 15734 11624 15786
rect 11624 15734 11676 15786
rect 11676 15734 11678 15786
rect 11622 15732 11678 15734
rect 11622 15662 11678 15664
rect 11622 15610 11624 15662
rect 11624 15610 11676 15662
rect 11676 15610 11678 15662
rect 11622 15608 11678 15610
rect 11622 15538 11678 15540
rect 11622 15486 11624 15538
rect 11624 15486 11676 15538
rect 11676 15486 11678 15538
rect 11622 15484 11678 15486
rect 12070 16902 12126 16904
rect 12070 16850 12072 16902
rect 12072 16850 12124 16902
rect 12124 16850 12126 16902
rect 12070 16848 12126 16850
rect 12070 16778 12126 16780
rect 12070 16726 12072 16778
rect 12072 16726 12124 16778
rect 12124 16726 12126 16778
rect 12070 16724 12126 16726
rect 12070 16654 12126 16656
rect 12070 16602 12072 16654
rect 12072 16602 12124 16654
rect 12124 16602 12126 16654
rect 12070 16600 12126 16602
rect 12070 16530 12126 16532
rect 12070 16478 12072 16530
rect 12072 16478 12124 16530
rect 12124 16478 12126 16530
rect 12070 16476 12126 16478
rect 12070 16406 12126 16408
rect 12070 16354 12072 16406
rect 12072 16354 12124 16406
rect 12124 16354 12126 16406
rect 12070 16352 12126 16354
rect 12070 16282 12126 16284
rect 12070 16230 12072 16282
rect 12072 16230 12124 16282
rect 12124 16230 12126 16282
rect 12070 16228 12126 16230
rect 12070 16158 12126 16160
rect 12070 16106 12072 16158
rect 12072 16106 12124 16158
rect 12124 16106 12126 16158
rect 12070 16104 12126 16106
rect 12070 16034 12126 16036
rect 12070 15982 12072 16034
rect 12072 15982 12124 16034
rect 12124 15982 12126 16034
rect 12070 15980 12126 15982
rect 12070 15910 12126 15912
rect 12070 15858 12072 15910
rect 12072 15858 12124 15910
rect 12124 15858 12126 15910
rect 12070 15856 12126 15858
rect 12070 15786 12126 15788
rect 12070 15734 12072 15786
rect 12072 15734 12124 15786
rect 12124 15734 12126 15786
rect 12070 15732 12126 15734
rect 12070 15662 12126 15664
rect 12070 15610 12072 15662
rect 12072 15610 12124 15662
rect 12124 15610 12126 15662
rect 12070 15608 12126 15610
rect 12070 15538 12126 15540
rect 12070 15486 12072 15538
rect 12072 15486 12124 15538
rect 12124 15486 12126 15538
rect 12070 15484 12126 15486
rect 12742 16902 12798 16904
rect 12742 16850 12744 16902
rect 12744 16850 12796 16902
rect 12796 16850 12798 16902
rect 12742 16848 12798 16850
rect 12742 16778 12798 16780
rect 12742 16726 12744 16778
rect 12744 16726 12796 16778
rect 12796 16726 12798 16778
rect 12742 16724 12798 16726
rect 12742 16654 12798 16656
rect 12742 16602 12744 16654
rect 12744 16602 12796 16654
rect 12796 16602 12798 16654
rect 12742 16600 12798 16602
rect 12742 16530 12798 16532
rect 12742 16478 12744 16530
rect 12744 16478 12796 16530
rect 12796 16478 12798 16530
rect 12742 16476 12798 16478
rect 12742 16406 12798 16408
rect 12742 16354 12744 16406
rect 12744 16354 12796 16406
rect 12796 16354 12798 16406
rect 12742 16352 12798 16354
rect 12742 16282 12798 16284
rect 12742 16230 12744 16282
rect 12744 16230 12796 16282
rect 12796 16230 12798 16282
rect 12742 16228 12798 16230
rect 12742 16158 12798 16160
rect 12742 16106 12744 16158
rect 12744 16106 12796 16158
rect 12796 16106 12798 16158
rect 12742 16104 12798 16106
rect 12742 16034 12798 16036
rect 12742 15982 12744 16034
rect 12744 15982 12796 16034
rect 12796 15982 12798 16034
rect 12742 15980 12798 15982
rect 12742 15910 12798 15912
rect 12742 15858 12744 15910
rect 12744 15858 12796 15910
rect 12796 15858 12798 15910
rect 12742 15856 12798 15858
rect 12742 15786 12798 15788
rect 12742 15734 12744 15786
rect 12744 15734 12796 15786
rect 12796 15734 12798 15786
rect 12742 15732 12798 15734
rect 12742 15662 12798 15664
rect 12742 15610 12744 15662
rect 12744 15610 12796 15662
rect 12796 15610 12798 15662
rect 12742 15608 12798 15610
rect 12742 15538 12798 15540
rect 12742 15486 12744 15538
rect 12744 15486 12796 15538
rect 12796 15486 12798 15538
rect 12742 15484 12798 15486
rect 13190 16902 13246 16904
rect 13190 16850 13192 16902
rect 13192 16850 13244 16902
rect 13244 16850 13246 16902
rect 13190 16848 13246 16850
rect 13190 16778 13246 16780
rect 13190 16726 13192 16778
rect 13192 16726 13244 16778
rect 13244 16726 13246 16778
rect 13190 16724 13246 16726
rect 13190 16654 13246 16656
rect 13190 16602 13192 16654
rect 13192 16602 13244 16654
rect 13244 16602 13246 16654
rect 13190 16600 13246 16602
rect 13190 16530 13246 16532
rect 13190 16478 13192 16530
rect 13192 16478 13244 16530
rect 13244 16478 13246 16530
rect 13190 16476 13246 16478
rect 13190 16406 13246 16408
rect 13190 16354 13192 16406
rect 13192 16354 13244 16406
rect 13244 16354 13246 16406
rect 13190 16352 13246 16354
rect 13190 16282 13246 16284
rect 13190 16230 13192 16282
rect 13192 16230 13244 16282
rect 13244 16230 13246 16282
rect 13190 16228 13246 16230
rect 13190 16158 13246 16160
rect 13190 16106 13192 16158
rect 13192 16106 13244 16158
rect 13244 16106 13246 16158
rect 13190 16104 13246 16106
rect 13190 16034 13246 16036
rect 13190 15982 13192 16034
rect 13192 15982 13244 16034
rect 13244 15982 13246 16034
rect 13190 15980 13246 15982
rect 13190 15910 13246 15912
rect 13190 15858 13192 15910
rect 13192 15858 13244 15910
rect 13244 15858 13246 15910
rect 13190 15856 13246 15858
rect 13190 15786 13246 15788
rect 13190 15734 13192 15786
rect 13192 15734 13244 15786
rect 13244 15734 13246 15786
rect 13190 15732 13246 15734
rect 13190 15662 13246 15664
rect 13190 15610 13192 15662
rect 13192 15610 13244 15662
rect 13244 15610 13246 15662
rect 13190 15608 13246 15610
rect 13190 15538 13246 15540
rect 13190 15486 13192 15538
rect 13192 15486 13244 15538
rect 13244 15486 13246 15538
rect 13190 15484 13246 15486
rect 13862 16902 13918 16904
rect 13862 16850 13864 16902
rect 13864 16850 13916 16902
rect 13916 16850 13918 16902
rect 13862 16848 13918 16850
rect 13862 16778 13918 16780
rect 13862 16726 13864 16778
rect 13864 16726 13916 16778
rect 13916 16726 13918 16778
rect 13862 16724 13918 16726
rect 13862 16654 13918 16656
rect 13862 16602 13864 16654
rect 13864 16602 13916 16654
rect 13916 16602 13918 16654
rect 13862 16600 13918 16602
rect 13862 16530 13918 16532
rect 13862 16478 13864 16530
rect 13864 16478 13916 16530
rect 13916 16478 13918 16530
rect 13862 16476 13918 16478
rect 13862 16406 13918 16408
rect 13862 16354 13864 16406
rect 13864 16354 13916 16406
rect 13916 16354 13918 16406
rect 13862 16352 13918 16354
rect 13862 16282 13918 16284
rect 13862 16230 13864 16282
rect 13864 16230 13916 16282
rect 13916 16230 13918 16282
rect 13862 16228 13918 16230
rect 13862 16158 13918 16160
rect 13862 16106 13864 16158
rect 13864 16106 13916 16158
rect 13916 16106 13918 16158
rect 13862 16104 13918 16106
rect 13862 16034 13918 16036
rect 13862 15982 13864 16034
rect 13864 15982 13916 16034
rect 13916 15982 13918 16034
rect 13862 15980 13918 15982
rect 13862 15910 13918 15912
rect 13862 15858 13864 15910
rect 13864 15858 13916 15910
rect 13916 15858 13918 15910
rect 13862 15856 13918 15858
rect 13862 15786 13918 15788
rect 13862 15734 13864 15786
rect 13864 15734 13916 15786
rect 13916 15734 13918 15786
rect 13862 15732 13918 15734
rect 13862 15662 13918 15664
rect 13862 15610 13864 15662
rect 13864 15610 13916 15662
rect 13916 15610 13918 15662
rect 13862 15608 13918 15610
rect 13862 15538 13918 15540
rect 13862 15486 13864 15538
rect 13864 15486 13916 15538
rect 13916 15486 13918 15538
rect 13862 15484 13918 15486
rect 14310 16902 14366 16904
rect 14310 16850 14312 16902
rect 14312 16850 14364 16902
rect 14364 16850 14366 16902
rect 14310 16848 14366 16850
rect 14310 16778 14366 16780
rect 14310 16726 14312 16778
rect 14312 16726 14364 16778
rect 14364 16726 14366 16778
rect 14310 16724 14366 16726
rect 14310 16654 14366 16656
rect 14310 16602 14312 16654
rect 14312 16602 14364 16654
rect 14364 16602 14366 16654
rect 14310 16600 14366 16602
rect 14310 16530 14366 16532
rect 14310 16478 14312 16530
rect 14312 16478 14364 16530
rect 14364 16478 14366 16530
rect 14310 16476 14366 16478
rect 14310 16406 14366 16408
rect 14310 16354 14312 16406
rect 14312 16354 14364 16406
rect 14364 16354 14366 16406
rect 14310 16352 14366 16354
rect 14310 16282 14366 16284
rect 14310 16230 14312 16282
rect 14312 16230 14364 16282
rect 14364 16230 14366 16282
rect 14310 16228 14366 16230
rect 14310 16158 14366 16160
rect 14310 16106 14312 16158
rect 14312 16106 14364 16158
rect 14364 16106 14366 16158
rect 14310 16104 14366 16106
rect 14310 16034 14366 16036
rect 14310 15982 14312 16034
rect 14312 15982 14364 16034
rect 14364 15982 14366 16034
rect 14310 15980 14366 15982
rect 14310 15910 14366 15912
rect 14310 15858 14312 15910
rect 14312 15858 14364 15910
rect 14364 15858 14366 15910
rect 14310 15856 14366 15858
rect 14310 15786 14366 15788
rect 14310 15734 14312 15786
rect 14312 15734 14364 15786
rect 14364 15734 14366 15786
rect 14310 15732 14366 15734
rect 14310 15662 14366 15664
rect 14310 15610 14312 15662
rect 14312 15610 14364 15662
rect 14364 15610 14366 15662
rect 14310 15608 14366 15610
rect 14310 15538 14366 15540
rect 14310 15486 14312 15538
rect 14312 15486 14364 15538
rect 14364 15486 14366 15538
rect 14310 15484 14366 15486
rect 14982 16902 15038 16904
rect 14982 16850 14984 16902
rect 14984 16850 15036 16902
rect 15036 16850 15038 16902
rect 14982 16848 15038 16850
rect 14982 16778 15038 16780
rect 14982 16726 14984 16778
rect 14984 16726 15036 16778
rect 15036 16726 15038 16778
rect 14982 16724 15038 16726
rect 14982 16654 15038 16656
rect 14982 16602 14984 16654
rect 14984 16602 15036 16654
rect 15036 16602 15038 16654
rect 14982 16600 15038 16602
rect 14982 16530 15038 16532
rect 14982 16478 14984 16530
rect 14984 16478 15036 16530
rect 15036 16478 15038 16530
rect 14982 16476 15038 16478
rect 14982 16406 15038 16408
rect 14982 16354 14984 16406
rect 14984 16354 15036 16406
rect 15036 16354 15038 16406
rect 14982 16352 15038 16354
rect 14982 16282 15038 16284
rect 14982 16230 14984 16282
rect 14984 16230 15036 16282
rect 15036 16230 15038 16282
rect 14982 16228 15038 16230
rect 14982 16158 15038 16160
rect 14982 16106 14984 16158
rect 14984 16106 15036 16158
rect 15036 16106 15038 16158
rect 14982 16104 15038 16106
rect 14982 16034 15038 16036
rect 14982 15982 14984 16034
rect 14984 15982 15036 16034
rect 15036 15982 15038 16034
rect 14982 15980 15038 15982
rect 14982 15910 15038 15912
rect 14982 15858 14984 15910
rect 14984 15858 15036 15910
rect 15036 15858 15038 15910
rect 14982 15856 15038 15858
rect 14982 15786 15038 15788
rect 14982 15734 14984 15786
rect 14984 15734 15036 15786
rect 15036 15734 15038 15786
rect 14982 15732 15038 15734
rect 14982 15662 15038 15664
rect 14982 15610 14984 15662
rect 14984 15610 15036 15662
rect 15036 15610 15038 15662
rect 14982 15608 15038 15610
rect 14982 15538 15038 15540
rect 14982 15486 14984 15538
rect 14984 15486 15036 15538
rect 15036 15486 15038 15538
rect 14982 15484 15038 15486
rect 15430 16902 15486 16904
rect 15430 16850 15432 16902
rect 15432 16850 15484 16902
rect 15484 16850 15486 16902
rect 15430 16848 15486 16850
rect 15430 16778 15486 16780
rect 15430 16726 15432 16778
rect 15432 16726 15484 16778
rect 15484 16726 15486 16778
rect 15430 16724 15486 16726
rect 15430 16654 15486 16656
rect 15430 16602 15432 16654
rect 15432 16602 15484 16654
rect 15484 16602 15486 16654
rect 15430 16600 15486 16602
rect 15430 16530 15486 16532
rect 15430 16478 15432 16530
rect 15432 16478 15484 16530
rect 15484 16478 15486 16530
rect 15430 16476 15486 16478
rect 15430 16406 15486 16408
rect 15430 16354 15432 16406
rect 15432 16354 15484 16406
rect 15484 16354 15486 16406
rect 15430 16352 15486 16354
rect 15430 16282 15486 16284
rect 15430 16230 15432 16282
rect 15432 16230 15484 16282
rect 15484 16230 15486 16282
rect 15430 16228 15486 16230
rect 15430 16158 15486 16160
rect 15430 16106 15432 16158
rect 15432 16106 15484 16158
rect 15484 16106 15486 16158
rect 15430 16104 15486 16106
rect 15430 16034 15486 16036
rect 15430 15982 15432 16034
rect 15432 15982 15484 16034
rect 15484 15982 15486 16034
rect 15430 15980 15486 15982
rect 15430 15910 15486 15912
rect 15430 15858 15432 15910
rect 15432 15858 15484 15910
rect 15484 15858 15486 15910
rect 15430 15856 15486 15858
rect 15430 15786 15486 15788
rect 15430 15734 15432 15786
rect 15432 15734 15484 15786
rect 15484 15734 15486 15786
rect 15430 15732 15486 15734
rect 15430 15662 15486 15664
rect 15430 15610 15432 15662
rect 15432 15610 15484 15662
rect 15484 15610 15486 15662
rect 15430 15608 15486 15610
rect 15430 15538 15486 15540
rect 15430 15486 15432 15538
rect 15432 15486 15484 15538
rect 15484 15486 15486 15538
rect 15430 15484 15486 15486
rect 16102 16902 16158 16904
rect 16102 16850 16104 16902
rect 16104 16850 16156 16902
rect 16156 16850 16158 16902
rect 16102 16848 16158 16850
rect 16102 16778 16158 16780
rect 16102 16726 16104 16778
rect 16104 16726 16156 16778
rect 16156 16726 16158 16778
rect 16102 16724 16158 16726
rect 16102 16654 16158 16656
rect 16102 16602 16104 16654
rect 16104 16602 16156 16654
rect 16156 16602 16158 16654
rect 16102 16600 16158 16602
rect 16102 16530 16158 16532
rect 16102 16478 16104 16530
rect 16104 16478 16156 16530
rect 16156 16478 16158 16530
rect 16102 16476 16158 16478
rect 16102 16406 16158 16408
rect 16102 16354 16104 16406
rect 16104 16354 16156 16406
rect 16156 16354 16158 16406
rect 16102 16352 16158 16354
rect 16102 16282 16158 16284
rect 16102 16230 16104 16282
rect 16104 16230 16156 16282
rect 16156 16230 16158 16282
rect 16102 16228 16158 16230
rect 16102 16158 16158 16160
rect 16102 16106 16104 16158
rect 16104 16106 16156 16158
rect 16156 16106 16158 16158
rect 16102 16104 16158 16106
rect 16102 16034 16158 16036
rect 16102 15982 16104 16034
rect 16104 15982 16156 16034
rect 16156 15982 16158 16034
rect 16102 15980 16158 15982
rect 16102 15910 16158 15912
rect 16102 15858 16104 15910
rect 16104 15858 16156 15910
rect 16156 15858 16158 15910
rect 16102 15856 16158 15858
rect 16102 15786 16158 15788
rect 16102 15734 16104 15786
rect 16104 15734 16156 15786
rect 16156 15734 16158 15786
rect 16102 15732 16158 15734
rect 16102 15662 16158 15664
rect 16102 15610 16104 15662
rect 16104 15610 16156 15662
rect 16156 15610 16158 15662
rect 16102 15608 16158 15610
rect 16102 15538 16158 15540
rect 16102 15486 16104 15538
rect 16104 15486 16156 15538
rect 16156 15486 16158 15538
rect 16102 15484 16158 15486
rect 16550 16902 16606 16904
rect 16550 16850 16552 16902
rect 16552 16850 16604 16902
rect 16604 16850 16606 16902
rect 16550 16848 16606 16850
rect 16550 16778 16606 16780
rect 16550 16726 16552 16778
rect 16552 16726 16604 16778
rect 16604 16726 16606 16778
rect 16550 16724 16606 16726
rect 16550 16654 16606 16656
rect 16550 16602 16552 16654
rect 16552 16602 16604 16654
rect 16604 16602 16606 16654
rect 16550 16600 16606 16602
rect 16550 16530 16606 16532
rect 16550 16478 16552 16530
rect 16552 16478 16604 16530
rect 16604 16478 16606 16530
rect 16550 16476 16606 16478
rect 16550 16406 16606 16408
rect 16550 16354 16552 16406
rect 16552 16354 16604 16406
rect 16604 16354 16606 16406
rect 16550 16352 16606 16354
rect 16550 16282 16606 16284
rect 16550 16230 16552 16282
rect 16552 16230 16604 16282
rect 16604 16230 16606 16282
rect 16550 16228 16606 16230
rect 16550 16158 16606 16160
rect 16550 16106 16552 16158
rect 16552 16106 16604 16158
rect 16604 16106 16606 16158
rect 16550 16104 16606 16106
rect 16550 16034 16606 16036
rect 16550 15982 16552 16034
rect 16552 15982 16604 16034
rect 16604 15982 16606 16034
rect 16550 15980 16606 15982
rect 16550 15910 16606 15912
rect 16550 15858 16552 15910
rect 16552 15858 16604 15910
rect 16604 15858 16606 15910
rect 16550 15856 16606 15858
rect 16550 15786 16606 15788
rect 16550 15734 16552 15786
rect 16552 15734 16604 15786
rect 16604 15734 16606 15786
rect 16550 15732 16606 15734
rect 16550 15662 16606 15664
rect 16550 15610 16552 15662
rect 16552 15610 16604 15662
rect 16604 15610 16606 15662
rect 16550 15608 16606 15610
rect 16550 15538 16606 15540
rect 16550 15486 16552 15538
rect 16552 15486 16604 15538
rect 16604 15486 16606 15538
rect 16550 15484 16606 15486
rect 17222 16902 17278 16904
rect 17222 16850 17224 16902
rect 17224 16850 17276 16902
rect 17276 16850 17278 16902
rect 17222 16848 17278 16850
rect 17222 16778 17278 16780
rect 17222 16726 17224 16778
rect 17224 16726 17276 16778
rect 17276 16726 17278 16778
rect 17222 16724 17278 16726
rect 17222 16654 17278 16656
rect 17222 16602 17224 16654
rect 17224 16602 17276 16654
rect 17276 16602 17278 16654
rect 17222 16600 17278 16602
rect 17222 16530 17278 16532
rect 17222 16478 17224 16530
rect 17224 16478 17276 16530
rect 17276 16478 17278 16530
rect 17222 16476 17278 16478
rect 17222 16406 17278 16408
rect 17222 16354 17224 16406
rect 17224 16354 17276 16406
rect 17276 16354 17278 16406
rect 17222 16352 17278 16354
rect 17222 16282 17278 16284
rect 17222 16230 17224 16282
rect 17224 16230 17276 16282
rect 17276 16230 17278 16282
rect 17222 16228 17278 16230
rect 17222 16158 17278 16160
rect 17222 16106 17224 16158
rect 17224 16106 17276 16158
rect 17276 16106 17278 16158
rect 17222 16104 17278 16106
rect 17222 16034 17278 16036
rect 17222 15982 17224 16034
rect 17224 15982 17276 16034
rect 17276 15982 17278 16034
rect 17222 15980 17278 15982
rect 17222 15910 17278 15912
rect 17222 15858 17224 15910
rect 17224 15858 17276 15910
rect 17276 15858 17278 15910
rect 17222 15856 17278 15858
rect 17222 15786 17278 15788
rect 17222 15734 17224 15786
rect 17224 15734 17276 15786
rect 17276 15734 17278 15786
rect 17222 15732 17278 15734
rect 17222 15662 17278 15664
rect 17222 15610 17224 15662
rect 17224 15610 17276 15662
rect 17276 15610 17278 15662
rect 17222 15608 17278 15610
rect 17222 15538 17278 15540
rect 17222 15486 17224 15538
rect 17224 15486 17276 15538
rect 17276 15486 17278 15538
rect 17222 15484 17278 15486
rect 17670 16902 17726 16904
rect 17670 16850 17672 16902
rect 17672 16850 17724 16902
rect 17724 16850 17726 16902
rect 17670 16848 17726 16850
rect 17670 16778 17726 16780
rect 17670 16726 17672 16778
rect 17672 16726 17724 16778
rect 17724 16726 17726 16778
rect 17670 16724 17726 16726
rect 17670 16654 17726 16656
rect 17670 16602 17672 16654
rect 17672 16602 17724 16654
rect 17724 16602 17726 16654
rect 17670 16600 17726 16602
rect 17670 16530 17726 16532
rect 17670 16478 17672 16530
rect 17672 16478 17724 16530
rect 17724 16478 17726 16530
rect 17670 16476 17726 16478
rect 17670 16406 17726 16408
rect 17670 16354 17672 16406
rect 17672 16354 17724 16406
rect 17724 16354 17726 16406
rect 17670 16352 17726 16354
rect 17670 16282 17726 16284
rect 17670 16230 17672 16282
rect 17672 16230 17724 16282
rect 17724 16230 17726 16282
rect 17670 16228 17726 16230
rect 17670 16158 17726 16160
rect 17670 16106 17672 16158
rect 17672 16106 17724 16158
rect 17724 16106 17726 16158
rect 17670 16104 17726 16106
rect 17670 16034 17726 16036
rect 17670 15982 17672 16034
rect 17672 15982 17724 16034
rect 17724 15982 17726 16034
rect 17670 15980 17726 15982
rect 17670 15910 17726 15912
rect 17670 15858 17672 15910
rect 17672 15858 17724 15910
rect 17724 15858 17726 15910
rect 17670 15856 17726 15858
rect 17670 15786 17726 15788
rect 17670 15734 17672 15786
rect 17672 15734 17724 15786
rect 17724 15734 17726 15786
rect 17670 15732 17726 15734
rect 17670 15662 17726 15664
rect 17670 15610 17672 15662
rect 17672 15610 17724 15662
rect 17724 15610 17726 15662
rect 17670 15608 17726 15610
rect 17670 15538 17726 15540
rect 17670 15486 17672 15538
rect 17672 15486 17724 15538
rect 17724 15486 17726 15538
rect 17670 15484 17726 15486
rect 18342 16902 18398 16904
rect 18342 16850 18344 16902
rect 18344 16850 18396 16902
rect 18396 16850 18398 16902
rect 18342 16848 18398 16850
rect 18342 16778 18398 16780
rect 18342 16726 18344 16778
rect 18344 16726 18396 16778
rect 18396 16726 18398 16778
rect 18342 16724 18398 16726
rect 18342 16654 18398 16656
rect 18342 16602 18344 16654
rect 18344 16602 18396 16654
rect 18396 16602 18398 16654
rect 18342 16600 18398 16602
rect 18342 16530 18398 16532
rect 18342 16478 18344 16530
rect 18344 16478 18396 16530
rect 18396 16478 18398 16530
rect 18342 16476 18398 16478
rect 18342 16406 18398 16408
rect 18342 16354 18344 16406
rect 18344 16354 18396 16406
rect 18396 16354 18398 16406
rect 18342 16352 18398 16354
rect 18342 16282 18398 16284
rect 18342 16230 18344 16282
rect 18344 16230 18396 16282
rect 18396 16230 18398 16282
rect 18342 16228 18398 16230
rect 18342 16158 18398 16160
rect 18342 16106 18344 16158
rect 18344 16106 18396 16158
rect 18396 16106 18398 16158
rect 18342 16104 18398 16106
rect 18342 16034 18398 16036
rect 18342 15982 18344 16034
rect 18344 15982 18396 16034
rect 18396 15982 18398 16034
rect 18342 15980 18398 15982
rect 18342 15910 18398 15912
rect 18342 15858 18344 15910
rect 18344 15858 18396 15910
rect 18396 15858 18398 15910
rect 18342 15856 18398 15858
rect 18342 15786 18398 15788
rect 18342 15734 18344 15786
rect 18344 15734 18396 15786
rect 18396 15734 18398 15786
rect 18342 15732 18398 15734
rect 18342 15662 18398 15664
rect 18342 15610 18344 15662
rect 18344 15610 18396 15662
rect 18396 15610 18398 15662
rect 18342 15608 18398 15610
rect 18342 15538 18398 15540
rect 18342 15486 18344 15538
rect 18344 15486 18396 15538
rect 18396 15486 18398 15538
rect 18342 15484 18398 15486
rect 18790 16902 18846 16904
rect 18790 16850 18792 16902
rect 18792 16850 18844 16902
rect 18844 16850 18846 16902
rect 18790 16848 18846 16850
rect 18790 16778 18846 16780
rect 18790 16726 18792 16778
rect 18792 16726 18844 16778
rect 18844 16726 18846 16778
rect 18790 16724 18846 16726
rect 18790 16654 18846 16656
rect 18790 16602 18792 16654
rect 18792 16602 18844 16654
rect 18844 16602 18846 16654
rect 18790 16600 18846 16602
rect 18790 16530 18846 16532
rect 18790 16478 18792 16530
rect 18792 16478 18844 16530
rect 18844 16478 18846 16530
rect 18790 16476 18846 16478
rect 18790 16406 18846 16408
rect 18790 16354 18792 16406
rect 18792 16354 18844 16406
rect 18844 16354 18846 16406
rect 18790 16352 18846 16354
rect 18790 16282 18846 16284
rect 18790 16230 18792 16282
rect 18792 16230 18844 16282
rect 18844 16230 18846 16282
rect 18790 16228 18846 16230
rect 18790 16158 18846 16160
rect 18790 16106 18792 16158
rect 18792 16106 18844 16158
rect 18844 16106 18846 16158
rect 18790 16104 18846 16106
rect 18790 16034 18846 16036
rect 18790 15982 18792 16034
rect 18792 15982 18844 16034
rect 18844 15982 18846 16034
rect 18790 15980 18846 15982
rect 18790 15910 18846 15912
rect 18790 15858 18792 15910
rect 18792 15858 18844 15910
rect 18844 15858 18846 15910
rect 18790 15856 18846 15858
rect 18790 15786 18846 15788
rect 18790 15734 18792 15786
rect 18792 15734 18844 15786
rect 18844 15734 18846 15786
rect 18790 15732 18846 15734
rect 18790 15662 18846 15664
rect 18790 15610 18792 15662
rect 18792 15610 18844 15662
rect 18844 15610 18846 15662
rect 18790 15608 18846 15610
rect 18790 15538 18846 15540
rect 18790 15486 18792 15538
rect 18792 15486 18844 15538
rect 18844 15486 18846 15538
rect 18790 15484 18846 15486
rect 19462 16902 19518 16904
rect 19462 16850 19464 16902
rect 19464 16850 19516 16902
rect 19516 16850 19518 16902
rect 19462 16848 19518 16850
rect 19462 16778 19518 16780
rect 19462 16726 19464 16778
rect 19464 16726 19516 16778
rect 19516 16726 19518 16778
rect 19462 16724 19518 16726
rect 19462 16654 19518 16656
rect 19462 16602 19464 16654
rect 19464 16602 19516 16654
rect 19516 16602 19518 16654
rect 19462 16600 19518 16602
rect 19462 16530 19518 16532
rect 19462 16478 19464 16530
rect 19464 16478 19516 16530
rect 19516 16478 19518 16530
rect 19462 16476 19518 16478
rect 19462 16406 19518 16408
rect 19462 16354 19464 16406
rect 19464 16354 19516 16406
rect 19516 16354 19518 16406
rect 19462 16352 19518 16354
rect 19462 16282 19518 16284
rect 19462 16230 19464 16282
rect 19464 16230 19516 16282
rect 19516 16230 19518 16282
rect 19462 16228 19518 16230
rect 19462 16158 19518 16160
rect 19462 16106 19464 16158
rect 19464 16106 19516 16158
rect 19516 16106 19518 16158
rect 19462 16104 19518 16106
rect 19462 16034 19518 16036
rect 19462 15982 19464 16034
rect 19464 15982 19516 16034
rect 19516 15982 19518 16034
rect 19462 15980 19518 15982
rect 19462 15910 19518 15912
rect 19462 15858 19464 15910
rect 19464 15858 19516 15910
rect 19516 15858 19518 15910
rect 19462 15856 19518 15858
rect 19462 15786 19518 15788
rect 19462 15734 19464 15786
rect 19464 15734 19516 15786
rect 19516 15734 19518 15786
rect 19462 15732 19518 15734
rect 19462 15662 19518 15664
rect 19462 15610 19464 15662
rect 19464 15610 19516 15662
rect 19516 15610 19518 15662
rect 19462 15608 19518 15610
rect 19462 15538 19518 15540
rect 19462 15486 19464 15538
rect 19464 15486 19516 15538
rect 19516 15486 19518 15538
rect 19462 15484 19518 15486
rect 19910 16902 19966 16904
rect 19910 16850 19912 16902
rect 19912 16850 19964 16902
rect 19964 16850 19966 16902
rect 19910 16848 19966 16850
rect 19910 16778 19966 16780
rect 19910 16726 19912 16778
rect 19912 16726 19964 16778
rect 19964 16726 19966 16778
rect 19910 16724 19966 16726
rect 19910 16654 19966 16656
rect 19910 16602 19912 16654
rect 19912 16602 19964 16654
rect 19964 16602 19966 16654
rect 19910 16600 19966 16602
rect 19910 16530 19966 16532
rect 19910 16478 19912 16530
rect 19912 16478 19964 16530
rect 19964 16478 19966 16530
rect 19910 16476 19966 16478
rect 19910 16406 19966 16408
rect 19910 16354 19912 16406
rect 19912 16354 19964 16406
rect 19964 16354 19966 16406
rect 19910 16352 19966 16354
rect 19910 16282 19966 16284
rect 19910 16230 19912 16282
rect 19912 16230 19964 16282
rect 19964 16230 19966 16282
rect 19910 16228 19966 16230
rect 19910 16158 19966 16160
rect 19910 16106 19912 16158
rect 19912 16106 19964 16158
rect 19964 16106 19966 16158
rect 19910 16104 19966 16106
rect 19910 16034 19966 16036
rect 19910 15982 19912 16034
rect 19912 15982 19964 16034
rect 19964 15982 19966 16034
rect 19910 15980 19966 15982
rect 19910 15910 19966 15912
rect 19910 15858 19912 15910
rect 19912 15858 19964 15910
rect 19964 15858 19966 15910
rect 19910 15856 19966 15858
rect 19910 15786 19966 15788
rect 19910 15734 19912 15786
rect 19912 15734 19964 15786
rect 19964 15734 19966 15786
rect 19910 15732 19966 15734
rect 19910 15662 19966 15664
rect 19910 15610 19912 15662
rect 19912 15610 19964 15662
rect 19964 15610 19966 15662
rect 19910 15608 19966 15610
rect 19910 15538 19966 15540
rect 19910 15486 19912 15538
rect 19912 15486 19964 15538
rect 19964 15486 19966 15538
rect 19910 15484 19966 15486
rect 10277 14878 10333 14934
rect 10725 14878 10781 14934
rect 9158 14572 9160 14594
rect 9160 14572 9212 14594
rect 9212 14572 9214 14594
rect 9158 14538 9214 14572
rect 9605 14572 9608 14594
rect 9608 14572 9660 14594
rect 9660 14572 9661 14594
rect 9605 14538 9661 14572
rect 8038 14252 8094 14253
rect 8038 14200 8040 14252
rect 8040 14200 8092 14252
rect 8092 14200 8094 14252
rect 8038 14197 8094 14200
rect 8486 14252 8542 14253
rect 8486 14200 8488 14252
rect 8488 14200 8540 14252
rect 8540 14200 8542 14252
rect 8486 14197 8542 14200
rect 6918 13880 6974 13913
rect 6918 13857 6920 13880
rect 6920 13857 6972 13880
rect 6972 13857 6974 13880
rect 7366 13880 7422 13913
rect 7366 13857 7368 13880
rect 7368 13857 7420 13880
rect 7420 13857 7422 13880
rect 5798 13517 5854 13573
rect 6246 13517 6302 13573
rect 4678 13208 4680 13233
rect 4680 13208 4732 13233
rect 4732 13208 4734 13233
rect 4678 13177 4734 13208
rect 5126 13208 5128 13233
rect 5128 13208 5180 13233
rect 5180 13208 5182 13233
rect 5126 13177 5182 13208
rect 3558 12888 3614 12893
rect 3558 12837 3560 12888
rect 3560 12837 3612 12888
rect 3612 12837 3614 12888
rect 4006 12888 4062 12893
rect 4006 12837 4008 12888
rect 4008 12837 4060 12888
rect 4060 12837 4062 12888
rect 2438 12497 2494 12553
rect 2886 12497 2942 12553
rect 2005 12096 2061 12152
rect 2005 11911 2061 11934
rect 2005 11878 2008 11911
rect 2008 11878 2060 11911
rect 2060 11878 2061 11911
rect 3125 11794 3181 11850
rect 3337 11794 3393 11850
rect 4245 11566 4301 11622
rect 4245 11348 4301 11404
rect 5364 11377 5420 11433
rect 5576 11377 5632 11433
rect 6379 11169 6435 11225
rect 6591 11169 6647 11225
rect 7499 10960 7555 11016
rect 7711 10960 7767 11016
rect 9317 10960 9373 11016
rect 9529 10960 9585 11016
rect 8426 10752 8482 10808
rect 8638 10752 8694 10808
rect 7789 10543 7845 10599
rect 8001 10543 8057 10599
rect 2402 9364 2458 9366
rect 2402 9312 2404 9364
rect 2404 9312 2456 9364
rect 2456 9312 2458 9364
rect 2402 9310 2458 9312
rect 2609 9364 2665 9366
rect 2609 9312 2611 9364
rect 2611 9312 2663 9364
rect 2663 9312 2665 9364
rect 2609 9310 2665 9312
rect 2402 9146 2458 9148
rect 2402 9094 2404 9146
rect 2404 9094 2456 9146
rect 2456 9094 2458 9146
rect 2402 9092 2458 9094
rect 2609 9146 2665 9148
rect 2609 9094 2611 9146
rect 2611 9094 2663 9146
rect 2663 9094 2665 9146
rect 2609 9092 2665 9094
rect 2402 8928 2458 8930
rect 2402 8876 2404 8928
rect 2404 8876 2456 8928
rect 2456 8876 2458 8928
rect 2402 8874 2458 8876
rect 2609 8928 2665 8930
rect 2609 8876 2611 8928
rect 2611 8876 2663 8928
rect 2663 8876 2665 8928
rect 2609 8874 2665 8876
rect 2402 8710 2458 8712
rect 2402 8658 2404 8710
rect 2404 8658 2456 8710
rect 2456 8658 2458 8710
rect 2402 8656 2458 8658
rect 2609 8710 2665 8712
rect 2609 8658 2611 8710
rect 2611 8658 2663 8710
rect 2663 8658 2665 8710
rect 2609 8656 2665 8658
rect 3129 9364 3185 9366
rect 3129 9312 3131 9364
rect 3131 9312 3183 9364
rect 3183 9312 3185 9364
rect 3129 9310 3185 9312
rect 3129 9146 3185 9148
rect 3129 9094 3131 9146
rect 3131 9094 3183 9146
rect 3183 9094 3185 9146
rect 3129 9092 3185 9094
rect 3129 8928 3185 8930
rect 3129 8876 3131 8928
rect 3131 8876 3183 8928
rect 3183 8876 3185 8928
rect 3129 8874 3185 8876
rect 3129 8710 3185 8712
rect 3129 8658 3131 8710
rect 3131 8658 3183 8710
rect 3183 8658 3185 8710
rect 3129 8656 3185 8658
rect 4093 9364 4149 9366
rect 4093 9312 4095 9364
rect 4095 9312 4147 9364
rect 4147 9312 4149 9364
rect 4093 9310 4149 9312
rect 4300 9364 4356 9366
rect 4300 9312 4302 9364
rect 4302 9312 4354 9364
rect 4354 9312 4356 9364
rect 4300 9310 4356 9312
rect 4093 9146 4149 9148
rect 4093 9094 4095 9146
rect 4095 9094 4147 9146
rect 4147 9094 4149 9146
rect 4093 9092 4149 9094
rect 4300 9146 4356 9148
rect 4300 9094 4302 9146
rect 4302 9094 4354 9146
rect 4354 9094 4356 9146
rect 4300 9092 4356 9094
rect 4093 8928 4149 8930
rect 4093 8876 4095 8928
rect 4095 8876 4147 8928
rect 4147 8876 4149 8928
rect 4093 8874 4149 8876
rect 4300 8928 4356 8930
rect 4300 8876 4302 8928
rect 4302 8876 4354 8928
rect 4354 8876 4356 8928
rect 4300 8874 4356 8876
rect 4093 8710 4149 8712
rect 4093 8658 4095 8710
rect 4095 8658 4147 8710
rect 4147 8658 4149 8710
rect 4093 8656 4149 8658
rect 4300 8710 4356 8712
rect 4300 8658 4302 8710
rect 4302 8658 4354 8710
rect 4354 8658 4356 8710
rect 4300 8656 4356 8658
rect 4820 9364 4876 9366
rect 4820 9312 4822 9364
rect 4822 9312 4874 9364
rect 4874 9312 4876 9364
rect 4820 9310 4876 9312
rect 4820 9146 4876 9148
rect 4820 9094 4822 9146
rect 4822 9094 4874 9146
rect 4874 9094 4876 9146
rect 4820 9092 4876 9094
rect 4820 8928 4876 8930
rect 4820 8876 4822 8928
rect 4822 8876 4874 8928
rect 4874 8876 4876 8928
rect 4820 8874 4876 8876
rect 4820 8710 4876 8712
rect 4820 8658 4822 8710
rect 4822 8658 4874 8710
rect 4874 8658 4876 8710
rect 4820 8656 4876 8658
rect 5784 9364 5840 9366
rect 5784 9312 5786 9364
rect 5786 9312 5838 9364
rect 5838 9312 5840 9364
rect 5784 9310 5840 9312
rect 5991 9364 6047 9366
rect 5991 9312 5993 9364
rect 5993 9312 6045 9364
rect 6045 9312 6047 9364
rect 5991 9310 6047 9312
rect 5784 9146 5840 9148
rect 5784 9094 5786 9146
rect 5786 9094 5838 9146
rect 5838 9094 5840 9146
rect 5784 9092 5840 9094
rect 5991 9146 6047 9148
rect 5991 9094 5993 9146
rect 5993 9094 6045 9146
rect 6045 9094 6047 9146
rect 5991 9092 6047 9094
rect 5784 8928 5840 8930
rect 5784 8876 5786 8928
rect 5786 8876 5838 8928
rect 5838 8876 5840 8928
rect 5784 8874 5840 8876
rect 5991 8928 6047 8930
rect 5991 8876 5993 8928
rect 5993 8876 6045 8928
rect 6045 8876 6047 8928
rect 5991 8874 6047 8876
rect 5784 8710 5840 8712
rect 5784 8658 5786 8710
rect 5786 8658 5838 8710
rect 5838 8658 5840 8710
rect 5784 8656 5840 8658
rect 5991 8710 6047 8712
rect 5991 8658 5993 8710
rect 5993 8658 6045 8710
rect 6045 8658 6047 8710
rect 5991 8656 6047 8658
rect 6511 9364 6567 9366
rect 6511 9312 6513 9364
rect 6513 9312 6565 9364
rect 6565 9312 6567 9364
rect 6511 9310 6567 9312
rect 6511 9146 6567 9148
rect 6511 9094 6513 9146
rect 6513 9094 6565 9146
rect 6565 9094 6567 9146
rect 6511 9092 6567 9094
rect 6511 8928 6567 8930
rect 6511 8876 6513 8928
rect 6513 8876 6565 8928
rect 6565 8876 6567 8928
rect 6511 8874 6567 8876
rect 6511 8710 6567 8712
rect 6511 8658 6513 8710
rect 6513 8658 6565 8710
rect 6565 8658 6567 8710
rect 6511 8656 6567 8658
rect 7669 9324 7725 9326
rect 7669 9272 7671 9324
rect 7671 9272 7723 9324
rect 7723 9272 7725 9324
rect 7669 9270 7725 9272
rect 7669 9106 7725 9108
rect 7669 9054 7671 9106
rect 7671 9054 7723 9106
rect 7723 9054 7725 9106
rect 7669 9052 7725 9054
rect 7669 8888 7725 8890
rect 7669 8836 7671 8888
rect 7671 8836 7723 8888
rect 7723 8836 7725 8888
rect 7669 8834 7725 8836
rect 7669 8670 7725 8672
rect 7669 8618 7671 8670
rect 7671 8618 7723 8670
rect 7723 8618 7725 8670
rect 7669 8616 7725 8618
rect 8117 9324 8173 9326
rect 8117 9272 8119 9324
rect 8119 9272 8171 9324
rect 8171 9272 8173 9324
rect 8117 9270 8173 9272
rect 8117 9106 8173 9108
rect 8117 9054 8119 9106
rect 8119 9054 8171 9106
rect 8171 9054 8173 9106
rect 8117 9052 8173 9054
rect 8117 8888 8173 8890
rect 8117 8836 8119 8888
rect 8119 8836 8171 8888
rect 8171 8836 8173 8888
rect 8117 8834 8173 8836
rect 8117 8670 8173 8672
rect 8117 8618 8119 8670
rect 8119 8618 8171 8670
rect 8171 8618 8173 8670
rect 8117 8616 8173 8618
rect 8565 9324 8621 9326
rect 8565 9272 8567 9324
rect 8567 9272 8619 9324
rect 8619 9272 8621 9324
rect 8565 9270 8621 9272
rect 8565 9106 8621 9108
rect 8565 9054 8567 9106
rect 8567 9054 8619 9106
rect 8619 9054 8621 9106
rect 8565 9052 8621 9054
rect 8565 8888 8621 8890
rect 8565 8836 8567 8888
rect 8567 8836 8619 8888
rect 8619 8836 8621 8888
rect 8565 8834 8621 8836
rect 8565 8670 8621 8672
rect 8565 8618 8567 8670
rect 8567 8618 8619 8670
rect 8619 8618 8621 8670
rect 8565 8616 8621 8618
rect 9302 9324 9358 9326
rect 9302 9272 9304 9324
rect 9304 9272 9356 9324
rect 9356 9272 9358 9324
rect 9302 9270 9358 9272
rect 9302 9106 9358 9108
rect 9302 9054 9304 9106
rect 9304 9054 9356 9106
rect 9356 9054 9358 9106
rect 9302 9052 9358 9054
rect 9302 8888 9358 8890
rect 9302 8836 9304 8888
rect 9304 8836 9356 8888
rect 9356 8836 9358 8888
rect 9302 8834 9358 8836
rect 9302 8670 9358 8672
rect 9302 8618 9304 8670
rect 9304 8618 9356 8670
rect 9356 8618 9358 8670
rect 9302 8616 9358 8618
rect 19237 14878 19293 14934
rect 19685 14878 19741 14934
rect 18117 14572 18120 14594
rect 18120 14572 18172 14594
rect 18172 14572 18173 14594
rect 18117 14538 18173 14572
rect 18565 14572 18568 14594
rect 18568 14572 18620 14594
rect 18620 14572 18621 14594
rect 18565 14538 18621 14572
rect 16997 14252 17053 14253
rect 16997 14200 17000 14252
rect 17000 14200 17052 14252
rect 17052 14200 17053 14252
rect 16997 14197 17053 14200
rect 17445 14252 17501 14253
rect 17445 14200 17448 14252
rect 17448 14200 17500 14252
rect 17500 14200 17501 14252
rect 17445 14197 17501 14200
rect 15877 13880 15933 13913
rect 15877 13857 15880 13880
rect 15880 13857 15932 13880
rect 15932 13857 15933 13880
rect 16325 13880 16381 13913
rect 16325 13857 16328 13880
rect 16328 13857 16380 13880
rect 16380 13857 16381 13880
rect 14757 13517 14813 13573
rect 15205 13517 15261 13573
rect 13637 13208 13640 13233
rect 13640 13208 13692 13233
rect 13692 13208 13693 13233
rect 13637 13177 13693 13208
rect 14085 13208 14088 13233
rect 14088 13208 14140 13233
rect 14140 13208 14141 13233
rect 14085 13177 14141 13208
rect 12517 12888 12573 12893
rect 12517 12837 12520 12888
rect 12520 12837 12572 12888
rect 12572 12837 12573 12888
rect 12965 12888 13021 12893
rect 12965 12837 12968 12888
rect 12968 12837 13020 12888
rect 13020 12837 13021 12888
rect 11397 12497 11453 12553
rect 11845 12497 11901 12553
rect 10964 12003 11020 12059
rect 11176 12003 11232 12059
rect 11619 11586 11675 11642
rect 10951 11377 11007 11433
rect 11163 11377 11219 11433
rect 10268 11169 10324 11225
rect 10480 11169 10536 11225
rect 9844 10543 9900 10599
rect 10056 10543 10112 10599
rect 9750 9324 9806 9326
rect 9750 9272 9752 9324
rect 9752 9272 9804 9324
rect 9804 9272 9806 9324
rect 9750 9270 9806 9272
rect 9750 9106 9806 9108
rect 9750 9054 9752 9106
rect 9752 9054 9804 9106
rect 9804 9054 9806 9106
rect 9750 9052 9806 9054
rect 9750 8888 9806 8890
rect 9750 8836 9752 8888
rect 9752 8836 9804 8888
rect 9804 8836 9806 8888
rect 9750 8834 9806 8836
rect 9750 8670 9806 8672
rect 9750 8618 9752 8670
rect 9752 8618 9804 8670
rect 9804 8618 9806 8670
rect 9750 8616 9806 8618
rect 10198 9324 10254 9326
rect 10198 9272 10200 9324
rect 10200 9272 10252 9324
rect 10252 9272 10254 9324
rect 10198 9270 10254 9272
rect 10198 9106 10254 9108
rect 10198 9054 10200 9106
rect 10200 9054 10252 9106
rect 10252 9054 10254 9106
rect 10198 9052 10254 9054
rect 10198 8888 10254 8890
rect 10198 8836 10200 8888
rect 10200 8836 10252 8888
rect 10252 8836 10254 8888
rect 10198 8834 10254 8836
rect 10198 8670 10254 8672
rect 10198 8618 10200 8670
rect 10200 8618 10252 8670
rect 10252 8618 10254 8670
rect 10198 8616 10254 8618
rect 10936 9324 10992 9326
rect 10936 9272 10938 9324
rect 10938 9272 10990 9324
rect 10990 9272 10992 9324
rect 10936 9270 10992 9272
rect 10936 9106 10992 9108
rect 10936 9054 10938 9106
rect 10938 9054 10990 9106
rect 10990 9054 10992 9106
rect 10936 9052 10992 9054
rect 10936 8888 10992 8890
rect 10936 8836 10938 8888
rect 10938 8836 10990 8888
rect 10990 8836 10992 8888
rect 10936 8834 10992 8836
rect 10936 8670 10992 8672
rect 10936 8618 10938 8670
rect 10938 8618 10990 8670
rect 10990 8618 10992 8670
rect 10936 8616 10992 8618
rect 12084 11794 12140 11850
rect 12296 11794 12352 11850
rect 12741 12112 12797 12168
rect 12741 11894 12797 11950
rect 13204 11593 13260 11649
rect 13416 11593 13472 11649
rect 14325 11616 14381 11672
rect 14325 11398 14381 11454
rect 15445 11407 15501 11463
rect 15445 11189 15501 11245
rect 16565 11198 16621 11254
rect 16565 10980 16621 11036
rect 17685 10990 17741 11046
rect 17685 10772 17741 10828
rect 18805 10781 18861 10837
rect 18805 10563 18861 10619
rect 11384 9324 11440 9326
rect 11384 9272 11386 9324
rect 11386 9272 11438 9324
rect 11438 9272 11440 9324
rect 11384 9270 11440 9272
rect 11384 9106 11440 9108
rect 11384 9054 11386 9106
rect 11386 9054 11438 9106
rect 11438 9054 11440 9106
rect 11384 9052 11440 9054
rect 11384 8888 11440 8890
rect 11384 8836 11386 8888
rect 11386 8836 11438 8888
rect 11438 8836 11440 8888
rect 11384 8834 11440 8836
rect 11384 8670 11440 8672
rect 11384 8618 11386 8670
rect 11386 8618 11438 8670
rect 11438 8618 11440 8670
rect 11384 8616 11440 8618
rect 11832 9324 11888 9326
rect 11832 9272 11834 9324
rect 11834 9272 11886 9324
rect 11886 9272 11888 9324
rect 11832 9270 11888 9272
rect 11832 9106 11888 9108
rect 11832 9054 11834 9106
rect 11834 9054 11886 9106
rect 11886 9054 11888 9106
rect 11832 9052 11888 9054
rect 11832 8888 11888 8890
rect 11832 8836 11834 8888
rect 11834 8836 11886 8888
rect 11886 8836 11888 8888
rect 11832 8834 11888 8836
rect 11832 8670 11888 8672
rect 11832 8618 11834 8670
rect 11834 8618 11886 8670
rect 11886 8618 11888 8670
rect 11832 8616 11888 8618
rect 12570 9324 12626 9326
rect 12570 9272 12572 9324
rect 12572 9272 12624 9324
rect 12624 9272 12626 9324
rect 12570 9270 12626 9272
rect 12570 9106 12626 9108
rect 12570 9054 12572 9106
rect 12572 9054 12624 9106
rect 12624 9054 12626 9106
rect 12570 9052 12626 9054
rect 12570 8888 12626 8890
rect 12570 8836 12572 8888
rect 12572 8836 12624 8888
rect 12624 8836 12626 8888
rect 12570 8834 12626 8836
rect 12570 8670 12626 8672
rect 12570 8618 12572 8670
rect 12572 8618 12624 8670
rect 12624 8618 12626 8670
rect 12570 8616 12626 8618
rect 13018 9324 13074 9326
rect 13018 9272 13020 9324
rect 13020 9272 13072 9324
rect 13072 9272 13074 9324
rect 13018 9270 13074 9272
rect 13018 9106 13074 9108
rect 13018 9054 13020 9106
rect 13020 9054 13072 9106
rect 13072 9054 13074 9106
rect 13018 9052 13074 9054
rect 13018 8888 13074 8890
rect 13018 8836 13020 8888
rect 13020 8836 13072 8888
rect 13072 8836 13074 8888
rect 13018 8834 13074 8836
rect 13018 8670 13074 8672
rect 13018 8618 13020 8670
rect 13020 8618 13072 8670
rect 13072 8618 13074 8670
rect 13018 8616 13074 8618
rect 29559 28996 29615 28998
rect 29559 28944 29561 28996
rect 29561 28944 29613 28996
rect 29613 28944 29615 28996
rect 29559 28942 29615 28944
rect 29559 28778 29615 28780
rect 29559 28726 29561 28778
rect 29561 28726 29613 28778
rect 29613 28726 29615 28778
rect 29559 28724 29615 28726
rect 28627 9988 28683 10044
rect 28838 9988 28894 10044
rect 29050 9988 29106 10044
rect 29261 9988 29317 10044
rect 28627 9770 28683 9826
rect 28838 9770 28894 9826
rect 29050 9770 29106 9826
rect 29261 9770 29317 9826
rect 28627 9552 28683 9608
rect 28838 9552 28894 9608
rect 29050 9552 29106 9608
rect 29261 9552 29317 9608
rect 13466 9324 13522 9326
rect 13466 9272 13468 9324
rect 13468 9272 13520 9324
rect 13520 9272 13522 9324
rect 13466 9270 13522 9272
rect 13466 9106 13522 9108
rect 13466 9054 13468 9106
rect 13468 9054 13520 9106
rect 13520 9054 13522 9106
rect 13466 9052 13522 9054
rect 13466 8888 13522 8890
rect 13466 8836 13468 8888
rect 13468 8836 13520 8888
rect 13520 8836 13522 8888
rect 13466 8834 13522 8836
rect 13466 8670 13522 8672
rect 13466 8618 13468 8670
rect 13468 8618 13520 8670
rect 13520 8618 13522 8670
rect 13466 8616 13522 8618
rect 28627 9334 28683 9390
rect 28838 9334 28894 9390
rect 29050 9334 29106 9390
rect 29261 9334 29317 9390
rect 2622 7879 2678 7881
rect 2622 7827 2624 7879
rect 2624 7827 2676 7879
rect 2676 7827 2678 7879
rect 2622 7825 2678 7827
rect 2622 7662 2678 7664
rect 2622 7610 2624 7662
rect 2624 7610 2676 7662
rect 2676 7610 2678 7662
rect 2622 7608 2678 7610
rect 2622 7444 2678 7446
rect 2622 7392 2624 7444
rect 2624 7392 2676 7444
rect 2676 7392 2678 7444
rect 2622 7390 2678 7392
rect 2622 7226 2678 7228
rect 2622 7174 2624 7226
rect 2624 7174 2676 7226
rect 2676 7174 2678 7226
rect 2622 7172 2678 7174
rect 2622 7008 2678 7010
rect 2622 6956 2624 7008
rect 2624 6956 2676 7008
rect 2676 6956 2678 7008
rect 2622 6954 2678 6956
rect 2622 6791 2678 6793
rect 2622 6739 2624 6791
rect 2624 6739 2676 6791
rect 2676 6739 2678 6791
rect 2622 6737 2678 6739
rect 3136 7879 3192 7881
rect 3136 7827 3138 7879
rect 3138 7827 3190 7879
rect 3190 7827 3192 7879
rect 3136 7825 3192 7827
rect 3136 7662 3192 7664
rect 3136 7610 3138 7662
rect 3138 7610 3190 7662
rect 3190 7610 3192 7662
rect 3136 7608 3192 7610
rect 3136 7444 3192 7446
rect 3136 7392 3138 7444
rect 3138 7392 3190 7444
rect 3190 7392 3192 7444
rect 3136 7390 3192 7392
rect 3136 7226 3192 7228
rect 3136 7174 3138 7226
rect 3138 7174 3190 7226
rect 3190 7174 3192 7226
rect 3136 7172 3192 7174
rect 3136 7008 3192 7010
rect 3136 6956 3138 7008
rect 3138 6956 3190 7008
rect 3190 6956 3192 7008
rect 3136 6954 3192 6956
rect 3136 6791 3192 6793
rect 3136 6739 3138 6791
rect 3138 6739 3190 6791
rect 3190 6739 3192 6791
rect 3136 6737 3192 6739
rect 3615 5764 3671 5820
rect 3125 5288 3181 5344
rect 3125 5070 3181 5126
rect 3615 5546 3671 5602
rect 4313 7879 4369 7881
rect 4313 7827 4315 7879
rect 4315 7827 4367 7879
rect 4367 7827 4369 7879
rect 4313 7825 4369 7827
rect 4313 7662 4369 7664
rect 4313 7610 4315 7662
rect 4315 7610 4367 7662
rect 4367 7610 4369 7662
rect 4313 7608 4369 7610
rect 4313 7444 4369 7446
rect 4313 7392 4315 7444
rect 4315 7392 4367 7444
rect 4367 7392 4369 7444
rect 4313 7390 4369 7392
rect 4313 7226 4369 7228
rect 4313 7174 4315 7226
rect 4315 7174 4367 7226
rect 4367 7174 4369 7226
rect 4313 7172 4369 7174
rect 4313 7008 4369 7010
rect 4313 6956 4315 7008
rect 4315 6956 4367 7008
rect 4367 6956 4369 7008
rect 4313 6954 4369 6956
rect 4313 6791 4369 6793
rect 4313 6739 4315 6791
rect 4315 6739 4367 6791
rect 4367 6739 4369 6791
rect 4313 6737 4369 6739
rect 4827 7879 4883 7881
rect 4827 7827 4829 7879
rect 4829 7827 4881 7879
rect 4881 7827 4883 7879
rect 4827 7825 4883 7827
rect 4827 7662 4883 7664
rect 4827 7610 4829 7662
rect 4829 7610 4881 7662
rect 4881 7610 4883 7662
rect 4827 7608 4883 7610
rect 4827 7444 4883 7446
rect 4827 7392 4829 7444
rect 4829 7392 4881 7444
rect 4881 7392 4883 7444
rect 4827 7390 4883 7392
rect 4827 7226 4883 7228
rect 4827 7174 4829 7226
rect 4829 7174 4881 7226
rect 4881 7174 4883 7226
rect 4827 7172 4883 7174
rect 4827 7008 4883 7010
rect 4827 6956 4829 7008
rect 4829 6956 4881 7008
rect 4881 6956 4883 7008
rect 4827 6954 4883 6956
rect 4827 6791 4883 6793
rect 4827 6739 4829 6791
rect 4829 6739 4881 6791
rect 4881 6739 4883 6791
rect 4827 6737 4883 6739
rect 5306 5764 5362 5820
rect 4816 5288 4872 5344
rect 4816 5070 4872 5126
rect 5306 5546 5362 5602
rect 6004 7879 6060 7881
rect 6004 7827 6006 7879
rect 6006 7827 6058 7879
rect 6058 7827 6060 7879
rect 6004 7825 6060 7827
rect 6004 7662 6060 7664
rect 6004 7610 6006 7662
rect 6006 7610 6058 7662
rect 6058 7610 6060 7662
rect 6004 7608 6060 7610
rect 6004 7444 6060 7446
rect 6004 7392 6006 7444
rect 6006 7392 6058 7444
rect 6058 7392 6060 7444
rect 6004 7390 6060 7392
rect 6004 7226 6060 7228
rect 6004 7174 6006 7226
rect 6006 7174 6058 7226
rect 6058 7174 6060 7226
rect 6004 7172 6060 7174
rect 6004 7008 6060 7010
rect 6004 6956 6006 7008
rect 6006 6956 6058 7008
rect 6058 6956 6060 7008
rect 6004 6954 6060 6956
rect 6004 6791 6060 6793
rect 6004 6739 6006 6791
rect 6006 6739 6058 6791
rect 6058 6739 6060 6791
rect 6004 6737 6060 6739
rect 6518 7879 6574 7881
rect 6518 7827 6520 7879
rect 6520 7827 6572 7879
rect 6572 7827 6574 7879
rect 6518 7825 6574 7827
rect 6518 7662 6574 7664
rect 6518 7610 6520 7662
rect 6520 7610 6572 7662
rect 6572 7610 6574 7662
rect 6518 7608 6574 7610
rect 6518 7444 6574 7446
rect 6518 7392 6520 7444
rect 6520 7392 6572 7444
rect 6572 7392 6574 7444
rect 6518 7390 6574 7392
rect 7669 7819 7725 7821
rect 7669 7767 7671 7819
rect 7671 7767 7723 7819
rect 7723 7767 7725 7819
rect 7669 7765 7725 7767
rect 7669 7601 7725 7603
rect 7669 7549 7671 7601
rect 7671 7549 7723 7601
rect 7723 7549 7725 7601
rect 7669 7547 7725 7549
rect 7669 7383 7725 7385
rect 7669 7331 7671 7383
rect 7671 7331 7723 7383
rect 7723 7331 7725 7383
rect 7669 7329 7725 7331
rect 8117 7819 8173 7821
rect 8117 7767 8119 7819
rect 8119 7767 8171 7819
rect 8171 7767 8173 7819
rect 8117 7765 8173 7767
rect 8117 7601 8173 7603
rect 8117 7549 8119 7601
rect 8119 7549 8171 7601
rect 8171 7549 8173 7601
rect 8117 7547 8173 7549
rect 8117 7383 8173 7385
rect 8117 7331 8119 7383
rect 8119 7331 8171 7383
rect 8171 7331 8173 7383
rect 8117 7329 8173 7331
rect 8565 7819 8621 7821
rect 8565 7767 8567 7819
rect 8567 7767 8619 7819
rect 8619 7767 8621 7819
rect 8565 7765 8621 7767
rect 8565 7601 8621 7603
rect 8565 7549 8567 7601
rect 8567 7549 8619 7601
rect 8619 7549 8621 7601
rect 8565 7547 8621 7549
rect 8565 7383 8621 7385
rect 8565 7331 8567 7383
rect 8567 7331 8619 7383
rect 8619 7331 8621 7383
rect 8565 7329 8621 7331
rect 9302 7819 9358 7821
rect 9302 7767 9304 7819
rect 9304 7767 9356 7819
rect 9356 7767 9358 7819
rect 9302 7765 9358 7767
rect 9302 7601 9358 7603
rect 9302 7549 9304 7601
rect 9304 7549 9356 7601
rect 9356 7549 9358 7601
rect 9302 7547 9358 7549
rect 9302 7383 9358 7385
rect 9302 7331 9304 7383
rect 9304 7331 9356 7383
rect 9356 7331 9358 7383
rect 9302 7329 9358 7331
rect 9750 7819 9806 7821
rect 9750 7767 9752 7819
rect 9752 7767 9804 7819
rect 9804 7767 9806 7819
rect 9750 7765 9806 7767
rect 9750 7601 9806 7603
rect 9750 7549 9752 7601
rect 9752 7549 9804 7601
rect 9804 7549 9806 7601
rect 9750 7547 9806 7549
rect 9750 7383 9806 7385
rect 9750 7331 9752 7383
rect 9752 7331 9804 7383
rect 9804 7331 9806 7383
rect 9750 7329 9806 7331
rect 10198 7819 10254 7821
rect 10198 7767 10200 7819
rect 10200 7767 10252 7819
rect 10252 7767 10254 7819
rect 10198 7765 10254 7767
rect 10198 7601 10254 7603
rect 10198 7549 10200 7601
rect 10200 7549 10252 7601
rect 10252 7549 10254 7601
rect 10198 7547 10254 7549
rect 10198 7383 10254 7385
rect 10198 7331 10200 7383
rect 10200 7331 10252 7383
rect 10252 7331 10254 7383
rect 10198 7329 10254 7331
rect 10936 7819 10992 7821
rect 10936 7767 10938 7819
rect 10938 7767 10990 7819
rect 10990 7767 10992 7819
rect 10936 7765 10992 7767
rect 10936 7601 10992 7603
rect 10936 7549 10938 7601
rect 10938 7549 10990 7601
rect 10990 7549 10992 7601
rect 10936 7547 10992 7549
rect 10936 7383 10992 7385
rect 10936 7331 10938 7383
rect 10938 7331 10990 7383
rect 10990 7331 10992 7383
rect 10936 7329 10992 7331
rect 11384 7819 11440 7821
rect 11384 7767 11386 7819
rect 11386 7767 11438 7819
rect 11438 7767 11440 7819
rect 11384 7765 11440 7767
rect 11384 7601 11440 7603
rect 11384 7549 11386 7601
rect 11386 7549 11438 7601
rect 11438 7549 11440 7601
rect 11384 7547 11440 7549
rect 11384 7383 11440 7385
rect 11384 7331 11386 7383
rect 11386 7331 11438 7383
rect 11438 7331 11440 7383
rect 11384 7329 11440 7331
rect 11832 7819 11888 7821
rect 11832 7767 11834 7819
rect 11834 7767 11886 7819
rect 11886 7767 11888 7819
rect 11832 7765 11888 7767
rect 11832 7601 11888 7603
rect 11832 7549 11834 7601
rect 11834 7549 11886 7601
rect 11886 7549 11888 7601
rect 11832 7547 11888 7549
rect 11832 7383 11888 7385
rect 11832 7331 11834 7383
rect 11834 7331 11886 7383
rect 11886 7331 11888 7383
rect 11832 7329 11888 7331
rect 12570 7819 12626 7821
rect 12570 7767 12572 7819
rect 12572 7767 12624 7819
rect 12624 7767 12626 7819
rect 12570 7765 12626 7767
rect 12570 7601 12626 7603
rect 12570 7549 12572 7601
rect 12572 7549 12624 7601
rect 12624 7549 12626 7601
rect 12570 7547 12626 7549
rect 12570 7383 12626 7385
rect 12570 7331 12572 7383
rect 12572 7331 12624 7383
rect 12624 7331 12626 7383
rect 12570 7329 12626 7331
rect 13018 7819 13074 7821
rect 13018 7767 13020 7819
rect 13020 7767 13072 7819
rect 13072 7767 13074 7819
rect 13018 7765 13074 7767
rect 13018 7601 13074 7603
rect 13018 7549 13020 7601
rect 13020 7549 13072 7601
rect 13072 7549 13074 7601
rect 13018 7547 13074 7549
rect 13018 7383 13074 7385
rect 13018 7331 13020 7383
rect 13020 7331 13072 7383
rect 13072 7331 13074 7383
rect 13018 7329 13074 7331
rect 13466 7819 13522 7821
rect 13466 7767 13468 7819
rect 13468 7767 13520 7819
rect 13520 7767 13522 7819
rect 13466 7765 13522 7767
rect 13466 7601 13522 7603
rect 13466 7549 13468 7601
rect 13468 7549 13520 7601
rect 13520 7549 13522 7601
rect 13466 7547 13522 7549
rect 13466 7383 13522 7385
rect 13466 7331 13468 7383
rect 13468 7331 13520 7383
rect 13520 7331 13522 7383
rect 13466 7329 13522 7331
rect 6518 7226 6574 7228
rect 6518 7174 6520 7226
rect 6520 7174 6572 7226
rect 6572 7174 6574 7226
rect 6518 7172 6574 7174
rect 6518 7008 6574 7010
rect 6518 6956 6520 7008
rect 6520 6956 6572 7008
rect 6572 6956 6574 7008
rect 6518 6954 6574 6956
rect 6518 6791 6574 6793
rect 6518 6739 6520 6791
rect 6520 6739 6572 6791
rect 6572 6739 6574 6791
rect 6518 6737 6574 6739
rect 7673 6709 7729 6711
rect 7673 6657 7675 6709
rect 7675 6657 7727 6709
rect 7727 6657 7729 6709
rect 7673 6655 7729 6657
rect 7673 6492 7729 6494
rect 7673 6440 7675 6492
rect 7675 6440 7727 6492
rect 7727 6440 7729 6492
rect 7673 6438 7729 6440
rect 7673 6274 7729 6276
rect 7673 6222 7675 6274
rect 7675 6222 7727 6274
rect 7727 6222 7729 6274
rect 7673 6220 7729 6222
rect 7673 6056 7729 6058
rect 7673 6004 7675 6056
rect 7675 6004 7727 6056
rect 7727 6004 7729 6056
rect 7673 6002 7729 6004
rect 6997 5764 7053 5820
rect 7673 5839 7729 5841
rect 7673 5787 7675 5839
rect 7675 5787 7727 5839
rect 7727 5787 7729 5839
rect 7673 5785 7729 5787
rect 8117 6710 8173 6712
rect 8117 6658 8119 6710
rect 8119 6658 8171 6710
rect 8171 6658 8173 6710
rect 8117 6656 8173 6658
rect 8117 6492 8173 6494
rect 8117 6440 8119 6492
rect 8119 6440 8171 6492
rect 8171 6440 8173 6492
rect 8117 6438 8173 6440
rect 8117 6275 8173 6277
rect 8117 6223 8119 6275
rect 8119 6223 8171 6275
rect 8171 6223 8173 6275
rect 8117 6221 8173 6223
rect 8117 6057 8173 6059
rect 8117 6005 8119 6057
rect 8119 6005 8171 6057
rect 8171 6005 8173 6057
rect 8117 6003 8173 6005
rect 8117 5839 8173 5841
rect 8117 5787 8119 5839
rect 8119 5787 8171 5839
rect 8171 5787 8173 5839
rect 8117 5785 8173 5787
rect 6997 5546 7053 5602
rect 6507 5288 6563 5344
rect 6507 5070 6563 5126
rect 8561 6709 8617 6711
rect 8561 6657 8563 6709
rect 8563 6657 8615 6709
rect 8615 6657 8617 6709
rect 8561 6655 8617 6657
rect 8561 6492 8617 6494
rect 8561 6440 8563 6492
rect 8563 6440 8615 6492
rect 8615 6440 8617 6492
rect 8561 6438 8617 6440
rect 8561 6274 8617 6276
rect 8561 6222 8563 6274
rect 8563 6222 8615 6274
rect 8615 6222 8617 6274
rect 8561 6220 8617 6222
rect 8561 6056 8617 6058
rect 8561 6004 8563 6056
rect 8563 6004 8615 6056
rect 8615 6004 8617 6056
rect 8561 6002 8617 6004
rect 8561 5839 8617 5841
rect 8561 5787 8563 5839
rect 8563 5787 8615 5839
rect 8615 5787 8617 5839
rect 8561 5785 8617 5787
rect 9306 6709 9362 6711
rect 9306 6657 9308 6709
rect 9308 6657 9360 6709
rect 9360 6657 9362 6709
rect 9306 6655 9362 6657
rect 9306 6492 9362 6494
rect 9306 6440 9308 6492
rect 9308 6440 9360 6492
rect 9360 6440 9362 6492
rect 9306 6438 9362 6440
rect 9306 6274 9362 6276
rect 9306 6222 9308 6274
rect 9308 6222 9360 6274
rect 9360 6222 9362 6274
rect 9306 6220 9362 6222
rect 9306 6056 9362 6058
rect 9306 6004 9308 6056
rect 9308 6004 9360 6056
rect 9360 6004 9362 6056
rect 9306 6002 9362 6004
rect 9306 5839 9362 5841
rect 9306 5787 9308 5839
rect 9308 5787 9360 5839
rect 9360 5787 9362 5839
rect 9306 5785 9362 5787
rect 9750 6710 9806 6712
rect 9750 6658 9752 6710
rect 9752 6658 9804 6710
rect 9804 6658 9806 6710
rect 9750 6656 9806 6658
rect 9750 6492 9806 6494
rect 9750 6440 9752 6492
rect 9752 6440 9804 6492
rect 9804 6440 9806 6492
rect 9750 6438 9806 6440
rect 9750 6275 9806 6277
rect 9750 6223 9752 6275
rect 9752 6223 9804 6275
rect 9804 6223 9806 6275
rect 9750 6221 9806 6223
rect 9750 6057 9806 6059
rect 9750 6005 9752 6057
rect 9752 6005 9804 6057
rect 9804 6005 9806 6057
rect 9750 6003 9806 6005
rect 9750 5839 9806 5841
rect 9750 5787 9752 5839
rect 9752 5787 9804 5839
rect 9804 5787 9806 5839
rect 9750 5785 9806 5787
rect 8117 5622 8173 5624
rect 8117 5570 8119 5622
rect 8119 5570 8171 5622
rect 8171 5570 8173 5622
rect 8117 5568 8173 5570
rect 8117 5404 8173 5406
rect 8117 5352 8119 5404
rect 8119 5352 8171 5404
rect 8171 5352 8173 5404
rect 8117 5350 8173 5352
rect 10194 6709 10250 6711
rect 10194 6657 10196 6709
rect 10196 6657 10248 6709
rect 10248 6657 10250 6709
rect 10194 6655 10250 6657
rect 10194 6492 10250 6494
rect 10194 6440 10196 6492
rect 10196 6440 10248 6492
rect 10248 6440 10250 6492
rect 10194 6438 10250 6440
rect 10194 6274 10250 6276
rect 10194 6222 10196 6274
rect 10196 6222 10248 6274
rect 10248 6222 10250 6274
rect 10194 6220 10250 6222
rect 10194 6056 10250 6058
rect 10194 6004 10196 6056
rect 10196 6004 10248 6056
rect 10248 6004 10250 6056
rect 10194 6002 10250 6004
rect 10194 5839 10250 5841
rect 10194 5787 10196 5839
rect 10196 5787 10248 5839
rect 10248 5787 10250 5839
rect 10194 5785 10250 5787
rect 10940 6709 10996 6711
rect 10940 6657 10942 6709
rect 10942 6657 10994 6709
rect 10994 6657 10996 6709
rect 10940 6655 10996 6657
rect 10940 6492 10996 6494
rect 10940 6440 10942 6492
rect 10942 6440 10994 6492
rect 10994 6440 10996 6492
rect 10940 6438 10996 6440
rect 10940 6274 10996 6276
rect 10940 6222 10942 6274
rect 10942 6222 10994 6274
rect 10994 6222 10996 6274
rect 10940 6220 10996 6222
rect 10940 6056 10996 6058
rect 10940 6004 10942 6056
rect 10942 6004 10994 6056
rect 10994 6004 10996 6056
rect 10940 6002 10996 6004
rect 10940 5839 10996 5841
rect 10940 5787 10942 5839
rect 10942 5787 10994 5839
rect 10994 5787 10996 5839
rect 10940 5785 10996 5787
rect 11384 6710 11440 6712
rect 11384 6658 11386 6710
rect 11386 6658 11438 6710
rect 11438 6658 11440 6710
rect 11384 6656 11440 6658
rect 11384 6492 11440 6494
rect 11384 6440 11386 6492
rect 11386 6440 11438 6492
rect 11438 6440 11440 6492
rect 11384 6438 11440 6440
rect 11384 6275 11440 6277
rect 11384 6223 11386 6275
rect 11386 6223 11438 6275
rect 11438 6223 11440 6275
rect 11384 6221 11440 6223
rect 11384 6057 11440 6059
rect 11384 6005 11386 6057
rect 11386 6005 11438 6057
rect 11438 6005 11440 6057
rect 11384 6003 11440 6005
rect 11384 5839 11440 5841
rect 11384 5787 11386 5839
rect 11386 5787 11438 5839
rect 11438 5787 11440 5839
rect 11384 5785 11440 5787
rect 9750 5622 9806 5624
rect 9750 5570 9752 5622
rect 9752 5570 9804 5622
rect 9804 5570 9806 5622
rect 9750 5568 9806 5570
rect 9750 5404 9806 5406
rect 9750 5352 9752 5404
rect 9752 5352 9804 5404
rect 9804 5352 9806 5404
rect 9750 5350 9806 5352
rect 336 -1388 392 -1332
rect 548 -1388 604 -1332
rect 8117 3584 8173 3586
rect 8117 2596 8119 3584
rect 8119 2596 8171 3584
rect 8171 2596 8173 3584
rect 8117 2594 8173 2596
rect 11828 6709 11884 6711
rect 11828 6657 11830 6709
rect 11830 6657 11882 6709
rect 11882 6657 11884 6709
rect 11828 6655 11884 6657
rect 11828 6492 11884 6494
rect 11828 6440 11830 6492
rect 11830 6440 11882 6492
rect 11882 6440 11884 6492
rect 11828 6438 11884 6440
rect 11828 6274 11884 6276
rect 11828 6222 11830 6274
rect 11830 6222 11882 6274
rect 11882 6222 11884 6274
rect 11828 6220 11884 6222
rect 11828 6056 11884 6058
rect 11828 6004 11830 6056
rect 11830 6004 11882 6056
rect 11882 6004 11884 6056
rect 11828 6002 11884 6004
rect 11828 5839 11884 5841
rect 11828 5787 11830 5839
rect 11830 5787 11882 5839
rect 11882 5787 11884 5839
rect 11828 5785 11884 5787
rect 12574 6709 12630 6711
rect 12574 6657 12576 6709
rect 12576 6657 12628 6709
rect 12628 6657 12630 6709
rect 12574 6655 12630 6657
rect 12574 6492 12630 6494
rect 12574 6440 12576 6492
rect 12576 6440 12628 6492
rect 12628 6440 12630 6492
rect 12574 6438 12630 6440
rect 12574 6274 12630 6276
rect 12574 6222 12576 6274
rect 12576 6222 12628 6274
rect 12628 6222 12630 6274
rect 12574 6220 12630 6222
rect 12574 6056 12630 6058
rect 12574 6004 12576 6056
rect 12576 6004 12628 6056
rect 12628 6004 12630 6056
rect 12574 6002 12630 6004
rect 12574 5839 12630 5841
rect 12574 5787 12576 5839
rect 12576 5787 12628 5839
rect 12628 5787 12630 5839
rect 12574 5785 12630 5787
rect 13018 6710 13074 6712
rect 13018 6658 13020 6710
rect 13020 6658 13072 6710
rect 13072 6658 13074 6710
rect 13018 6656 13074 6658
rect 13018 6492 13074 6494
rect 13018 6440 13020 6492
rect 13020 6440 13072 6492
rect 13072 6440 13074 6492
rect 13018 6438 13074 6440
rect 13018 6275 13074 6277
rect 13018 6223 13020 6275
rect 13020 6223 13072 6275
rect 13072 6223 13074 6275
rect 13018 6221 13074 6223
rect 13018 6057 13074 6059
rect 13018 6005 13020 6057
rect 13020 6005 13072 6057
rect 13072 6005 13074 6057
rect 13018 6003 13074 6005
rect 13018 5839 13074 5841
rect 13018 5787 13020 5839
rect 13020 5787 13072 5839
rect 13072 5787 13074 5839
rect 13018 5785 13074 5787
rect 11384 5622 11440 5624
rect 11384 5570 11386 5622
rect 11386 5570 11438 5622
rect 11438 5570 11440 5622
rect 11384 5568 11440 5570
rect 11384 5404 11440 5406
rect 11384 5352 11386 5404
rect 11386 5352 11438 5404
rect 11438 5352 11440 5404
rect 11384 5350 11440 5352
rect 9751 3584 9807 3586
rect 9751 2596 9753 3584
rect 9753 2596 9805 3584
rect 9805 2596 9807 3584
rect 9751 2594 9807 2596
rect 13462 6709 13518 6711
rect 13462 6657 13464 6709
rect 13464 6657 13516 6709
rect 13516 6657 13518 6709
rect 13462 6655 13518 6657
rect 13462 6492 13518 6494
rect 13462 6440 13464 6492
rect 13464 6440 13516 6492
rect 13516 6440 13518 6492
rect 13462 6438 13518 6440
rect 13462 6274 13518 6276
rect 13462 6222 13464 6274
rect 13464 6222 13516 6274
rect 13516 6222 13518 6274
rect 13462 6220 13518 6222
rect 13462 6056 13518 6058
rect 13462 6004 13464 6056
rect 13464 6004 13516 6056
rect 13516 6004 13518 6056
rect 13462 6002 13518 6004
rect 13462 5839 13518 5841
rect 13462 5787 13464 5839
rect 13464 5787 13516 5839
rect 13516 5787 13518 5839
rect 13462 5785 13518 5787
rect 13018 5622 13074 5624
rect 13018 5570 13020 5622
rect 13020 5570 13072 5622
rect 13072 5570 13074 5622
rect 13018 5568 13074 5570
rect 13018 5404 13074 5406
rect 13018 5352 13020 5404
rect 13020 5352 13072 5404
rect 13072 5352 13074 5404
rect 13018 5350 13074 5352
rect 11384 3584 11440 3586
rect 11384 2596 11386 3584
rect 11386 2596 11438 3584
rect 11438 2596 11440 3584
rect 11384 2594 11440 2596
rect 13018 3584 13074 3586
rect 13018 2596 13020 3584
rect 13020 2596 13072 3584
rect 13072 2596 13074 3584
rect 13018 2594 13074 2596
rect 7836 1876 7892 1878
rect 7836 1824 7838 1876
rect 7838 1824 7890 1876
rect 7890 1824 7892 1876
rect 7836 1822 7892 1824
rect 7836 1658 7892 1660
rect 7836 1606 7838 1658
rect 7838 1606 7890 1658
rect 7890 1606 7892 1658
rect 7836 1604 7892 1606
rect 9898 2008 9954 2010
rect 9898 1956 9900 2008
rect 9900 1956 9952 2008
rect 9952 1956 9954 2008
rect 9898 1954 9954 1956
rect 10109 2008 10165 2010
rect 10109 1956 10111 2008
rect 10111 1956 10163 2008
rect 10163 1956 10165 2008
rect 10109 1954 10165 1956
rect 10319 2008 10375 2010
rect 10319 1956 10321 2008
rect 10321 1956 10373 2008
rect 10373 1956 10375 2008
rect 10319 1954 10375 1956
rect 10530 2008 10586 2010
rect 10530 1956 10532 2008
rect 10532 1956 10584 2008
rect 10584 1956 10586 2008
rect 10530 1954 10586 1956
rect 10741 2008 10797 2010
rect 10741 1956 10743 2008
rect 10743 1956 10795 2008
rect 10795 1956 10797 2008
rect 10741 1954 10797 1956
rect 10952 2008 11008 2010
rect 10952 1956 10954 2008
rect 10954 1956 11006 2008
rect 11006 1956 11008 2008
rect 10952 1954 11008 1956
rect 11163 2008 11219 2010
rect 11163 1956 11165 2008
rect 11165 1956 11217 2008
rect 11217 1956 11219 2008
rect 11163 1954 11219 1956
rect 11373 2008 11429 2010
rect 11373 1956 11375 2008
rect 11375 1956 11427 2008
rect 11427 1956 11429 2008
rect 11373 1954 11429 1956
rect 11584 2008 11640 2010
rect 11584 1956 11586 2008
rect 11586 1956 11638 2008
rect 11638 1956 11640 2008
rect 11584 1954 11640 1956
rect 11796 2008 11852 2010
rect 11796 1956 11798 2008
rect 11798 1956 11850 2008
rect 11850 1956 11852 2008
rect 11796 1954 11852 1956
rect 12007 2008 12063 2010
rect 12007 1956 12009 2008
rect 12009 1956 12061 2008
rect 12061 1956 12063 2008
rect 12007 1954 12063 1956
rect 12217 2008 12273 2010
rect 12217 1956 12219 2008
rect 12219 1956 12271 2008
rect 12271 1956 12273 2008
rect 12217 1954 12273 1956
rect 12428 2008 12484 2010
rect 12428 1956 12430 2008
rect 12430 1956 12482 2008
rect 12482 1956 12484 2008
rect 12428 1954 12484 1956
rect 12639 2008 12695 2010
rect 12639 1956 12641 2008
rect 12641 1956 12693 2008
rect 12693 1956 12695 2008
rect 12639 1954 12695 1956
rect 12850 2008 12906 2010
rect 12850 1956 12852 2008
rect 12852 1956 12904 2008
rect 12904 1956 12906 2008
rect 12850 1954 12906 1956
rect 13061 2008 13117 2010
rect 13061 1956 13063 2008
rect 13063 1956 13115 2008
rect 13115 1956 13117 2008
rect 13061 1954 13117 1956
rect 13271 2008 13327 2010
rect 13271 1956 13273 2008
rect 13273 1956 13325 2008
rect 13325 1956 13327 2008
rect 13271 1954 13327 1956
rect 13482 2008 13538 2010
rect 13482 1956 13484 2008
rect 13484 1956 13536 2008
rect 13536 1956 13538 2008
rect 13482 1954 13538 1956
rect 9898 1790 9954 1792
rect 9898 1738 9900 1790
rect 9900 1738 9952 1790
rect 9952 1738 9954 1790
rect 9898 1736 9954 1738
rect 10109 1790 10165 1792
rect 10109 1738 10111 1790
rect 10111 1738 10163 1790
rect 10163 1738 10165 1790
rect 10109 1736 10165 1738
rect 10319 1790 10375 1792
rect 10319 1738 10321 1790
rect 10321 1738 10373 1790
rect 10373 1738 10375 1790
rect 10319 1736 10375 1738
rect 10530 1790 10586 1792
rect 10530 1738 10532 1790
rect 10532 1738 10584 1790
rect 10584 1738 10586 1790
rect 10530 1736 10586 1738
rect 10741 1790 10797 1792
rect 10741 1738 10743 1790
rect 10743 1738 10795 1790
rect 10795 1738 10797 1790
rect 10741 1736 10797 1738
rect 10952 1790 11008 1792
rect 10952 1738 10954 1790
rect 10954 1738 11006 1790
rect 11006 1738 11008 1790
rect 10952 1736 11008 1738
rect 11163 1790 11219 1792
rect 11163 1738 11165 1790
rect 11165 1738 11217 1790
rect 11217 1738 11219 1790
rect 11163 1736 11219 1738
rect 11373 1790 11429 1792
rect 11373 1738 11375 1790
rect 11375 1738 11427 1790
rect 11427 1738 11429 1790
rect 11373 1736 11429 1738
rect 11584 1790 11640 1792
rect 11584 1738 11586 1790
rect 11586 1738 11638 1790
rect 11638 1738 11640 1790
rect 11584 1736 11640 1738
rect 11796 1790 11852 1792
rect 11796 1738 11798 1790
rect 11798 1738 11850 1790
rect 11850 1738 11852 1790
rect 11796 1736 11852 1738
rect 12007 1790 12063 1792
rect 12007 1738 12009 1790
rect 12009 1738 12061 1790
rect 12061 1738 12063 1790
rect 12007 1736 12063 1738
rect 12217 1790 12273 1792
rect 12217 1738 12219 1790
rect 12219 1738 12271 1790
rect 12271 1738 12273 1790
rect 12217 1736 12273 1738
rect 12428 1790 12484 1792
rect 12428 1738 12430 1790
rect 12430 1738 12482 1790
rect 12482 1738 12484 1790
rect 12428 1736 12484 1738
rect 12639 1790 12695 1792
rect 12639 1738 12641 1790
rect 12641 1738 12693 1790
rect 12693 1738 12695 1790
rect 12639 1736 12695 1738
rect 12850 1790 12906 1792
rect 12850 1738 12852 1790
rect 12852 1738 12904 1790
rect 12904 1738 12906 1790
rect 12850 1736 12906 1738
rect 13061 1790 13117 1792
rect 13061 1738 13063 1790
rect 13063 1738 13115 1790
rect 13115 1738 13117 1790
rect 13061 1736 13117 1738
rect 13271 1790 13327 1792
rect 13271 1738 13273 1790
rect 13273 1738 13325 1790
rect 13325 1738 13327 1790
rect 13271 1736 13327 1738
rect 13482 1790 13538 1792
rect 13482 1738 13484 1790
rect 13484 1738 13536 1790
rect 13536 1738 13538 1790
rect 13482 1736 13538 1738
rect 7445 1160 7501 1162
rect 7445 1108 7447 1160
rect 7447 1108 7499 1160
rect 7499 1108 7501 1160
rect 7445 1106 7501 1108
rect 7445 942 7501 944
rect 7445 890 7447 942
rect 7447 890 7499 942
rect 7499 890 7501 942
rect 7445 888 7501 890
rect 8472 1178 8528 1180
rect 8472 1126 8474 1178
rect 8474 1126 8526 1178
rect 8526 1126 8528 1178
rect 8472 1124 8528 1126
rect 8472 960 8528 962
rect 8472 908 8474 960
rect 8474 908 8526 960
rect 8526 908 8528 960
rect 8472 906 8528 908
rect 9658 1173 9714 1175
rect 9658 1121 9660 1173
rect 9660 1121 9712 1173
rect 9712 1121 9714 1173
rect 9658 1119 9714 1121
rect 9869 1173 9925 1175
rect 9869 1121 9871 1173
rect 9871 1121 9923 1173
rect 9923 1121 9925 1173
rect 9869 1119 9925 1121
rect 10080 1173 10136 1175
rect 10080 1121 10082 1173
rect 10082 1121 10134 1173
rect 10134 1121 10136 1173
rect 10080 1119 10136 1121
rect 10291 1173 10347 1175
rect 10291 1121 10293 1173
rect 10293 1121 10345 1173
rect 10345 1121 10347 1173
rect 10291 1119 10347 1121
rect 10502 1173 10558 1175
rect 10502 1121 10504 1173
rect 10504 1121 10556 1173
rect 10556 1121 10558 1173
rect 10502 1119 10558 1121
rect 10712 1173 10768 1175
rect 10712 1121 10714 1173
rect 10714 1121 10766 1173
rect 10766 1121 10768 1173
rect 10712 1119 10768 1121
rect 10923 1173 10979 1175
rect 10923 1121 10925 1173
rect 10925 1121 10977 1173
rect 10977 1121 10979 1173
rect 10923 1119 10979 1121
rect 11134 1173 11190 1175
rect 11134 1121 11136 1173
rect 11136 1121 11188 1173
rect 11188 1121 11190 1173
rect 11134 1119 11190 1121
rect 11345 1173 11401 1175
rect 11345 1121 11347 1173
rect 11347 1121 11399 1173
rect 11399 1121 11401 1173
rect 11345 1119 11401 1121
rect 11556 1173 11612 1175
rect 11556 1121 11558 1173
rect 11558 1121 11610 1173
rect 11610 1121 11612 1173
rect 11556 1119 11612 1121
rect 11767 1173 11823 1175
rect 11767 1121 11769 1173
rect 11769 1121 11821 1173
rect 11821 1121 11823 1173
rect 11767 1119 11823 1121
rect 11978 1173 12034 1175
rect 11978 1121 11980 1173
rect 11980 1121 12032 1173
rect 12032 1121 12034 1173
rect 11978 1119 12034 1121
rect 12189 1173 12245 1175
rect 12189 1121 12191 1173
rect 12191 1121 12243 1173
rect 12243 1121 12245 1173
rect 12189 1119 12245 1121
rect 12400 1173 12456 1175
rect 12400 1121 12402 1173
rect 12402 1121 12454 1173
rect 12454 1121 12456 1173
rect 12400 1119 12456 1121
rect 12610 1173 12666 1175
rect 12610 1121 12612 1173
rect 12612 1121 12664 1173
rect 12664 1121 12666 1173
rect 12610 1119 12666 1121
rect 12821 1173 12877 1175
rect 12821 1121 12823 1173
rect 12823 1121 12875 1173
rect 12875 1121 12877 1173
rect 12821 1119 12877 1121
rect 13032 1173 13088 1175
rect 13032 1121 13034 1173
rect 13034 1121 13086 1173
rect 13086 1121 13088 1173
rect 13032 1119 13088 1121
rect 13243 1173 13299 1175
rect 13243 1121 13245 1173
rect 13245 1121 13297 1173
rect 13297 1121 13299 1173
rect 13243 1119 13299 1121
rect 13454 1173 13510 1175
rect 13454 1121 13456 1173
rect 13456 1121 13508 1173
rect 13508 1121 13510 1173
rect 13454 1119 13510 1121
rect 9658 955 9714 957
rect 9658 903 9660 955
rect 9660 903 9712 955
rect 9712 903 9714 955
rect 9658 901 9714 903
rect 9869 955 9925 957
rect 9869 903 9871 955
rect 9871 903 9923 955
rect 9923 903 9925 955
rect 9869 901 9925 903
rect 10080 955 10136 957
rect 10080 903 10082 955
rect 10082 903 10134 955
rect 10134 903 10136 955
rect 10080 901 10136 903
rect 10291 955 10347 957
rect 10291 903 10293 955
rect 10293 903 10345 955
rect 10345 903 10347 955
rect 10291 901 10347 903
rect 10502 955 10558 957
rect 10502 903 10504 955
rect 10504 903 10556 955
rect 10556 903 10558 955
rect 10502 901 10558 903
rect 10712 955 10768 957
rect 10712 903 10714 955
rect 10714 903 10766 955
rect 10766 903 10768 955
rect 10712 901 10768 903
rect 10923 955 10979 957
rect 10923 903 10925 955
rect 10925 903 10977 955
rect 10977 903 10979 955
rect 10923 901 10979 903
rect 11134 955 11190 957
rect 11134 903 11136 955
rect 11136 903 11188 955
rect 11188 903 11190 955
rect 11134 901 11190 903
rect 11345 955 11401 957
rect 11345 903 11347 955
rect 11347 903 11399 955
rect 11399 903 11401 955
rect 11345 901 11401 903
rect 11556 955 11612 957
rect 11556 903 11558 955
rect 11558 903 11610 955
rect 11610 903 11612 955
rect 11556 901 11612 903
rect 11767 955 11823 957
rect 11767 903 11769 955
rect 11769 903 11821 955
rect 11821 903 11823 955
rect 11767 901 11823 903
rect 11978 955 12034 957
rect 11978 903 11980 955
rect 11980 903 12032 955
rect 12032 903 12034 955
rect 11978 901 12034 903
rect 12189 955 12245 957
rect 12189 903 12191 955
rect 12191 903 12243 955
rect 12243 903 12245 955
rect 12189 901 12245 903
rect 12400 955 12456 957
rect 12400 903 12402 955
rect 12402 903 12454 955
rect 12454 903 12456 955
rect 12400 901 12456 903
rect 12610 955 12666 957
rect 12610 903 12612 955
rect 12612 903 12664 955
rect 12664 903 12666 955
rect 12610 901 12666 903
rect 12821 955 12877 957
rect 12821 903 12823 955
rect 12823 903 12875 955
rect 12875 903 12877 955
rect 12821 901 12877 903
rect 13032 955 13088 957
rect 13032 903 13034 955
rect 13034 903 13086 955
rect 13086 903 13088 955
rect 13032 901 13088 903
rect 13243 955 13299 957
rect 13243 903 13245 955
rect 13245 903 13297 955
rect 13297 903 13299 955
rect 13243 901 13299 903
rect 13454 955 13510 957
rect 13454 903 13456 955
rect 13456 903 13508 955
rect 13508 903 13510 955
rect 13454 901 13510 903
rect 8064 -1388 8120 -1332
rect 8276 -1388 8332 -1332
rect 21660 615 21924 879
rect 21660 -453 21924 -189
rect 29453 -1388 29509 -1332
rect 29665 -1388 29721 -1332
<< metal3 >>
rect 645 30026 29412 30125
rect 645 29970 740 30026
rect 796 29970 951 30026
rect 1007 29970 1163 30026
rect 1219 29970 1374 30026
rect 1430 29970 5479 30026
rect 5535 29970 5691 30026
rect 5747 29970 16395 30026
rect 16451 29970 16607 30026
rect 16663 29970 23343 30026
rect 23399 29970 23555 30026
rect 23611 29970 28627 30026
rect 28683 29970 28838 30026
rect 28894 29970 29050 30026
rect 29106 29970 29261 30026
rect 29317 29970 29412 30026
rect 645 29808 29412 29970
rect 645 29752 740 29808
rect 796 29752 951 29808
rect 1007 29752 1163 29808
rect 1219 29752 1374 29808
rect 1430 29752 5479 29808
rect 5535 29752 5691 29808
rect 5747 29752 16395 29808
rect 16451 29752 16607 29808
rect 16663 29752 23343 29808
rect 23399 29752 23555 29808
rect 23611 29752 28627 29808
rect 28683 29752 28838 29808
rect 28894 29752 29050 29808
rect 29106 29752 29261 29808
rect 29317 29752 29412 29808
rect 645 29590 29412 29752
rect 645 29534 740 29590
rect 796 29534 951 29590
rect 1007 29534 1163 29590
rect 1219 29534 1374 29590
rect 1430 29534 5479 29590
rect 5535 29534 5691 29590
rect 5747 29534 16395 29590
rect 16451 29534 16607 29590
rect 16663 29534 23343 29590
rect 23399 29534 23555 29590
rect 23611 29534 28627 29590
rect 28683 29534 28838 29590
rect 28894 29534 29050 29590
rect 29106 29534 29261 29590
rect 29317 29534 29412 29590
rect 645 29372 29412 29534
rect 645 29316 740 29372
rect 796 29316 951 29372
rect 1007 29316 1163 29372
rect 1219 29316 1374 29372
rect 1430 29316 5479 29372
rect 5535 29316 5691 29372
rect 5747 29316 16395 29372
rect 16451 29316 16607 29372
rect 16663 29316 23343 29372
rect 23399 29316 23555 29372
rect 23611 29316 28627 29372
rect 28683 29316 28838 29372
rect 28894 29316 29050 29372
rect 29106 29316 29261 29372
rect 29317 29316 29412 29372
rect 645 29216 29412 29316
rect 6545 29037 6671 29038
rect 13923 29037 14049 29038
rect 24409 29037 24535 29038
rect 403 28999 29654 29037
rect 403 28998 6580 28999
rect 403 28942 442 28998
rect 498 28943 6580 28998
rect 6636 28943 13958 28999
rect 14014 28943 24444 28999
rect 24500 28998 29654 28999
rect 24500 28943 29559 28998
rect 498 28942 29559 28943
rect 29615 28942 29654 28998
rect 403 28781 29654 28942
rect 403 28780 6580 28781
rect 403 28724 442 28780
rect 498 28725 6580 28780
rect 6636 28725 13958 28781
rect 14014 28725 24444 28781
rect 24500 28780 29654 28781
rect 24500 28725 29559 28780
rect 498 28724 29559 28725
rect 29615 28724 29654 28780
rect 403 28686 29654 28724
rect 407 28685 533 28686
rect 29524 28685 29650 28686
rect 1393 28502 28604 28552
rect 1393 28446 1654 28502
rect 1710 28446 2094 28502
rect 2150 28446 3006 28502
rect 3062 28446 3446 28502
rect 3502 28446 3886 28502
rect 3942 28446 4798 28502
rect 4854 28446 5238 28502
rect 5294 28446 9033 28502
rect 9089 28446 9473 28502
rect 9529 28446 10385 28502
rect 10441 28446 10825 28502
rect 10881 28446 11265 28502
rect 11321 28446 12177 28502
rect 12233 28446 12617 28502
rect 12673 28446 28604 28502
rect 1393 28403 28604 28446
rect 1393 28347 5921 28403
rect 5977 28347 6360 28403
rect 6416 28347 13300 28403
rect 13356 28347 13739 28403
rect 13795 28394 23785 28403
rect 13795 28347 16916 28394
rect 1393 28346 16916 28347
rect 1393 28290 7744 28346
rect 7800 28290 15123 28346
rect 15179 28338 16916 28346
rect 16972 28338 17826 28394
rect 17882 28338 18550 28394
rect 18606 28338 19460 28394
rect 19516 28338 20183 28394
rect 20239 28338 21093 28394
rect 21149 28338 21817 28394
rect 21873 28338 22727 28394
rect 22783 28347 23785 28394
rect 23841 28347 24224 28403
rect 24280 28347 28604 28403
rect 22783 28346 28604 28347
rect 22783 28338 25608 28346
rect 15179 28290 25608 28338
rect 25664 28290 28604 28346
rect 1393 28284 28604 28290
rect 1393 28228 1654 28284
rect 1710 28228 2094 28284
rect 2150 28228 3006 28284
rect 3062 28228 3446 28284
rect 3502 28228 3886 28284
rect 3942 28228 4798 28284
rect 4854 28228 5238 28284
rect 5294 28228 9033 28284
rect 9089 28228 9473 28284
rect 9529 28228 10385 28284
rect 10441 28228 10825 28284
rect 10881 28228 11265 28284
rect 11321 28228 12177 28284
rect 12233 28228 12617 28284
rect 12673 28228 28604 28284
rect 1393 28185 28604 28228
rect 1393 28129 5921 28185
rect 5977 28129 6360 28185
rect 6416 28129 13300 28185
rect 13356 28129 13739 28185
rect 13795 28176 23785 28185
rect 13795 28129 16916 28176
rect 1393 28128 16916 28129
rect 1393 28072 7744 28128
rect 7800 28072 15123 28128
rect 15179 28120 16916 28128
rect 16972 28120 17826 28176
rect 17882 28120 18550 28176
rect 18606 28120 19460 28176
rect 19516 28120 20183 28176
rect 20239 28120 21093 28176
rect 21149 28120 21817 28176
rect 21873 28120 22727 28176
rect 22783 28129 23785 28176
rect 23841 28129 24224 28185
rect 24280 28129 28604 28185
rect 22783 28128 28604 28129
rect 22783 28120 25608 28128
rect 15179 28072 25608 28120
rect 25664 28072 28604 28128
rect 1393 28066 28604 28072
rect 1393 28010 1654 28066
rect 1710 28010 2094 28066
rect 2150 28010 3006 28066
rect 3062 28010 3446 28066
rect 3502 28010 3886 28066
rect 3942 28010 4798 28066
rect 4854 28010 5238 28066
rect 5294 28010 9033 28066
rect 9089 28010 9473 28066
rect 9529 28010 10385 28066
rect 10441 28010 10825 28066
rect 10881 28010 11265 28066
rect 11321 28010 12177 28066
rect 12233 28010 12617 28066
rect 12673 28010 28604 28066
rect 1393 27967 28604 28010
rect 1393 27911 5921 27967
rect 5977 27911 6360 27967
rect 6416 27911 13300 27967
rect 13356 27911 13739 27967
rect 13795 27958 23785 27967
rect 13795 27911 16916 27958
rect 1393 27910 16916 27911
rect 1393 27854 7744 27910
rect 7800 27854 15123 27910
rect 15179 27902 16916 27910
rect 16972 27902 17826 27958
rect 17882 27902 18550 27958
rect 18606 27902 19460 27958
rect 19516 27902 20183 27958
rect 20239 27902 21093 27958
rect 21149 27902 21817 27958
rect 21873 27902 22727 27958
rect 22783 27911 23785 27958
rect 23841 27911 24224 27967
rect 24280 27911 28604 27967
rect 22783 27910 28604 27911
rect 22783 27902 25608 27910
rect 15179 27854 25608 27902
rect 25664 27854 28604 27910
rect 1393 27848 28604 27854
rect 1393 27792 1654 27848
rect 1710 27792 2094 27848
rect 2150 27792 3006 27848
rect 3062 27792 3446 27848
rect 3502 27792 3886 27848
rect 3942 27792 4798 27848
rect 4854 27792 5238 27848
rect 5294 27792 9033 27848
rect 9089 27792 9473 27848
rect 9529 27792 10385 27848
rect 10441 27792 10825 27848
rect 10881 27792 11265 27848
rect 11321 27792 12177 27848
rect 12233 27792 12617 27848
rect 12673 27792 28604 27848
rect 1393 27740 28604 27792
rect 1393 27684 16916 27740
rect 16972 27684 17826 27740
rect 17882 27684 18550 27740
rect 18606 27684 19460 27740
rect 19516 27684 20183 27740
rect 20239 27684 21093 27740
rect 21149 27684 21817 27740
rect 21873 27684 22727 27740
rect 22783 27684 28604 27740
rect 1393 27601 28604 27684
rect 1393 27600 16441 27601
rect 23230 27600 28604 27601
rect 1393 27439 28604 27488
rect 1393 27394 24971 27439
rect 1393 27380 8134 27394
rect 1393 27355 5645 27380
rect 1393 27299 1654 27355
rect 1710 27299 2102 27355
rect 2158 27299 2550 27355
rect 2606 27299 2998 27355
rect 3054 27299 3446 27355
rect 3502 27299 3894 27355
rect 3950 27299 4342 27355
rect 4398 27299 4790 27355
rect 4846 27299 5238 27355
rect 5294 27324 5645 27355
rect 5701 27324 5921 27380
rect 5977 27338 8134 27380
rect 8190 27380 15513 27394
rect 8190 27355 13024 27380
rect 8190 27338 9033 27355
rect 5977 27324 9033 27338
rect 5294 27299 9033 27324
rect 9089 27299 9481 27355
rect 9537 27299 9929 27355
rect 9985 27299 10377 27355
rect 10433 27299 10825 27355
rect 10881 27299 11273 27355
rect 11329 27299 11721 27355
rect 11777 27299 12169 27355
rect 12225 27299 12617 27355
rect 12673 27324 13024 27355
rect 13080 27324 13300 27380
rect 13356 27338 15513 27380
rect 15569 27383 24971 27394
rect 25027 27394 28604 27439
rect 25027 27383 25999 27394
rect 15569 27380 25999 27383
rect 15569 27338 23785 27380
rect 13356 27324 23785 27338
rect 23841 27338 25999 27380
rect 26055 27338 28604 27394
rect 23841 27324 28604 27338
rect 12673 27299 28604 27324
rect 1393 27221 28604 27299
rect 1393 27212 24971 27221
rect 1393 27162 7005 27212
rect 1393 27137 5645 27162
rect 1393 27081 1654 27137
rect 1710 27081 2102 27137
rect 2158 27081 2550 27137
rect 2606 27081 2998 27137
rect 3054 27081 3446 27137
rect 3502 27081 3894 27137
rect 3950 27081 4342 27137
rect 4398 27081 4790 27137
rect 4846 27081 5238 27137
rect 5294 27106 5645 27137
rect 5701 27106 5921 27162
rect 5977 27156 7005 27162
rect 7061 27156 7217 27212
rect 7273 27176 14384 27212
rect 7273 27156 8134 27176
rect 5977 27120 8134 27156
rect 8190 27162 14384 27176
rect 8190 27137 13024 27162
rect 8190 27120 9033 27137
rect 5977 27106 9033 27120
rect 5294 27081 9033 27106
rect 9089 27081 9481 27137
rect 9537 27081 9929 27137
rect 9985 27081 10377 27137
rect 10433 27081 10825 27137
rect 10881 27081 11273 27137
rect 11329 27081 11721 27137
rect 11777 27081 12169 27137
rect 12225 27081 12617 27137
rect 12673 27106 13024 27137
rect 13080 27106 13300 27162
rect 13356 27156 14384 27162
rect 14440 27156 14596 27212
rect 14652 27176 24971 27212
rect 14652 27156 15513 27176
rect 13356 27120 15513 27156
rect 15569 27165 24971 27176
rect 25027 27176 28604 27221
rect 25027 27165 25999 27176
rect 15569 27162 25999 27165
rect 15569 27120 23785 27162
rect 13356 27106 23785 27120
rect 23841 27120 25999 27162
rect 26055 27120 28604 27176
rect 23841 27106 28604 27120
rect 12673 27081 28604 27106
rect 1393 26958 28604 27081
rect 1393 26944 8134 26958
rect 1393 26919 5645 26944
rect 1393 26863 1654 26919
rect 1710 26863 2102 26919
rect 2158 26863 2550 26919
rect 2606 26863 2998 26919
rect 3054 26863 3446 26919
rect 3502 26863 3894 26919
rect 3950 26863 4342 26919
rect 4398 26863 4790 26919
rect 4846 26863 5238 26919
rect 5294 26888 5645 26919
rect 5701 26888 5921 26944
rect 5977 26902 8134 26944
rect 8190 26944 15513 26958
rect 8190 26919 13024 26944
rect 8190 26902 9033 26919
rect 5977 26888 9033 26902
rect 5294 26863 9033 26888
rect 9089 26863 9481 26919
rect 9537 26863 9929 26919
rect 9985 26863 10377 26919
rect 10433 26863 10825 26919
rect 10881 26863 11273 26919
rect 11329 26863 11721 26919
rect 11777 26863 12169 26919
rect 12225 26863 12617 26919
rect 12673 26888 13024 26919
rect 13080 26888 13300 26944
rect 13356 26902 15513 26944
rect 15569 26902 28604 26958
rect 13356 26888 28604 26902
rect 12673 26863 28604 26888
rect 1393 26775 28604 26863
rect 1393 26537 28654 26641
rect 1393 26516 23737 26537
rect 1393 26460 5872 26516
rect 5928 26460 6079 26516
rect 6135 26493 7563 26516
rect 6135 26460 6599 26493
rect 1393 26437 6599 26460
rect 6655 26460 7563 26493
rect 7619 26460 7770 26516
rect 7826 26493 13251 26516
rect 7826 26460 8290 26493
rect 6655 26437 8290 26460
rect 8346 26460 13251 26493
rect 13307 26460 13458 26516
rect 13514 26493 14942 26516
rect 13514 26460 13978 26493
rect 8346 26437 13978 26460
rect 14034 26460 14942 26493
rect 14998 26460 15149 26516
rect 15205 26493 23737 26516
rect 15205 26460 15669 26493
rect 14034 26437 15669 26460
rect 15725 26481 23737 26493
rect 23793 26481 23944 26537
rect 24000 26481 24464 26537
rect 24520 26481 25427 26537
rect 25483 26481 25634 26537
rect 25690 26481 26154 26537
rect 26210 26481 27118 26537
rect 27174 26481 27325 26537
rect 27381 26481 27845 26537
rect 27901 26481 28654 26537
rect 15725 26437 28654 26481
rect 1393 26319 28654 26437
rect 1393 26298 23737 26319
rect 1393 26242 5872 26298
rect 5928 26242 6079 26298
rect 6135 26275 7563 26298
rect 6135 26242 6599 26275
rect 1393 26219 6599 26242
rect 6655 26242 7563 26275
rect 7619 26242 7770 26298
rect 7826 26275 13251 26298
rect 7826 26242 8290 26275
rect 6655 26219 8290 26242
rect 8346 26242 13251 26275
rect 13307 26242 13458 26298
rect 13514 26275 14942 26298
rect 13514 26242 13978 26275
rect 8346 26219 13978 26242
rect 14034 26242 14942 26275
rect 14998 26242 15149 26298
rect 15205 26275 23737 26298
rect 15205 26242 15669 26275
rect 14034 26219 15669 26242
rect 15725 26263 23737 26275
rect 23793 26263 23944 26319
rect 24000 26263 24464 26319
rect 24520 26263 25427 26319
rect 25483 26263 25634 26319
rect 25690 26263 26154 26319
rect 26210 26263 27118 26319
rect 27174 26263 27325 26319
rect 27381 26263 27845 26319
rect 27901 26263 28654 26319
rect 15725 26219 28654 26263
rect 1393 26101 28654 26219
rect 1393 26080 23737 26101
rect 1393 26024 5872 26080
rect 5928 26024 6079 26080
rect 6135 26057 7563 26080
rect 6135 26024 6599 26057
rect 1393 26001 6599 26024
rect 6655 26024 7563 26057
rect 7619 26024 7770 26080
rect 7826 26057 13251 26080
rect 7826 26024 8290 26057
rect 6655 26001 8290 26024
rect 8346 26024 13251 26057
rect 13307 26024 13458 26080
rect 13514 26057 14942 26080
rect 13514 26024 13978 26057
rect 8346 26001 13978 26024
rect 14034 26024 14942 26057
rect 14998 26024 15149 26080
rect 15205 26057 23737 26080
rect 15205 26024 15669 26057
rect 14034 26001 15669 26024
rect 15725 26045 23737 26057
rect 23793 26045 23944 26101
rect 24000 26045 24464 26101
rect 24520 26045 25427 26101
rect 25483 26045 25634 26101
rect 25690 26045 26154 26101
rect 26210 26045 27118 26101
rect 27174 26045 27325 26101
rect 27381 26045 27845 26101
rect 27901 26045 28654 26101
rect 15725 26001 28654 26045
rect 1393 25883 28654 26001
rect 1393 25862 23737 25883
rect 1393 25806 5872 25862
rect 5928 25806 6079 25862
rect 6135 25839 7563 25862
rect 6135 25806 6599 25839
rect 1393 25783 6599 25806
rect 6655 25806 7563 25839
rect 7619 25806 7770 25862
rect 7826 25839 13251 25862
rect 7826 25806 8290 25839
rect 6655 25783 8290 25806
rect 8346 25806 13251 25839
rect 13307 25806 13458 25862
rect 13514 25839 14942 25862
rect 13514 25806 13978 25839
rect 8346 25783 13978 25806
rect 14034 25806 14942 25839
rect 14998 25806 15149 25862
rect 15205 25839 23737 25862
rect 15205 25806 15669 25839
rect 14034 25783 15669 25806
rect 15725 25827 23737 25839
rect 23793 25827 23944 25883
rect 24000 25827 24464 25883
rect 24520 25827 25427 25883
rect 25483 25827 25634 25883
rect 25690 25827 26154 25883
rect 26210 25827 27118 25883
rect 27174 25827 27325 25883
rect 27381 25827 27845 25883
rect 27901 25827 28654 25883
rect 15725 25783 28654 25827
rect 1393 25732 28654 25783
rect 1393 25302 28672 25394
rect 1393 25246 16923 25302
rect 16979 25246 17371 25302
rect 17427 25246 17819 25302
rect 17875 25246 18557 25302
rect 18613 25246 19005 25302
rect 19061 25246 19453 25302
rect 19509 25246 20190 25302
rect 20246 25246 20638 25302
rect 20694 25246 21086 25302
rect 21142 25246 21824 25302
rect 21880 25246 22272 25302
rect 22328 25246 22720 25302
rect 22776 25246 28672 25302
rect 1393 25084 28672 25246
rect 1393 25028 16923 25084
rect 16979 25028 17371 25084
rect 17427 25028 17819 25084
rect 17875 25028 18557 25084
rect 18613 25028 19005 25084
rect 19061 25028 19453 25084
rect 19509 25028 20190 25084
rect 20246 25028 20638 25084
rect 20694 25028 21086 25084
rect 21142 25028 21824 25084
rect 21880 25028 22272 25084
rect 22328 25028 22720 25084
rect 22776 25028 28672 25084
rect 1393 24999 28672 25028
rect 1393 24943 23957 24999
rect 24013 24943 24471 24999
rect 24527 24943 25647 24999
rect 25703 24943 26161 24999
rect 26217 24943 27338 24999
rect 27394 24943 27852 24999
rect 27908 24943 28672 24999
rect 1393 24866 28672 24943
rect 1393 24813 16923 24866
rect 1393 24804 6606 24813
rect 1393 24775 6092 24804
rect 1393 24719 1815 24775
rect 1871 24719 2267 24775
rect 2323 24719 2550 24775
rect 2606 24719 2833 24775
rect 2889 24719 3285 24775
rect 3341 24719 3607 24775
rect 3663 24719 4059 24775
rect 4115 24719 4342 24775
rect 4398 24719 4625 24775
rect 4681 24719 5077 24775
rect 5133 24748 6092 24775
rect 6148 24757 6606 24804
rect 6662 24804 8297 24813
rect 6662 24757 7783 24804
rect 6148 24748 7783 24757
rect 7839 24757 8297 24804
rect 8353 24804 13985 24813
rect 8353 24775 13471 24804
rect 8353 24757 9194 24775
rect 7839 24748 9194 24757
rect 5133 24719 9194 24748
rect 9250 24719 9646 24775
rect 9702 24719 9929 24775
rect 9985 24719 10212 24775
rect 10268 24719 10664 24775
rect 10720 24719 10986 24775
rect 11042 24719 11438 24775
rect 11494 24719 11721 24775
rect 11777 24719 12004 24775
rect 12060 24719 12456 24775
rect 12512 24748 13471 24775
rect 13527 24757 13985 24804
rect 14041 24804 15676 24813
rect 14041 24757 15162 24804
rect 13527 24748 15162 24757
rect 15218 24757 15676 24804
rect 15732 24810 16923 24813
rect 16979 24810 17371 24866
rect 17427 24810 17819 24866
rect 17875 24810 18557 24866
rect 18613 24810 19005 24866
rect 19061 24810 19453 24866
rect 19509 24810 20190 24866
rect 20246 24810 20638 24866
rect 20694 24810 21086 24866
rect 21142 24810 21824 24866
rect 21880 24810 22272 24866
rect 22328 24810 22720 24866
rect 22776 24810 28672 24866
rect 15732 24782 28672 24810
rect 15732 24757 23957 24782
rect 15218 24748 23957 24757
rect 12512 24726 23957 24748
rect 24013 24726 24471 24782
rect 24527 24726 25647 24782
rect 25703 24726 26161 24782
rect 26217 24726 27338 24782
rect 27394 24726 27852 24782
rect 27908 24726 28672 24782
rect 12512 24719 28672 24726
rect 1393 24595 28672 24719
rect 1393 24587 6606 24595
rect 1393 24558 6092 24587
rect 1393 24502 1815 24558
rect 1871 24502 2267 24558
rect 2323 24502 2550 24558
rect 2606 24502 2833 24558
rect 2889 24502 3285 24558
rect 3341 24502 3607 24558
rect 3663 24502 4059 24558
rect 4115 24502 4342 24558
rect 4398 24502 4625 24558
rect 4681 24502 5077 24558
rect 5133 24531 6092 24558
rect 6148 24539 6606 24587
rect 6662 24587 8297 24595
rect 6662 24539 7783 24587
rect 6148 24531 7783 24539
rect 7839 24539 8297 24587
rect 8353 24587 13985 24595
rect 8353 24558 13471 24587
rect 8353 24539 9194 24558
rect 7839 24531 9194 24539
rect 5133 24502 9194 24531
rect 9250 24502 9646 24558
rect 9702 24502 9929 24558
rect 9985 24502 10212 24558
rect 10268 24502 10664 24558
rect 10720 24502 10986 24558
rect 11042 24502 11438 24558
rect 11494 24502 11721 24558
rect 11777 24502 12004 24558
rect 12060 24502 12456 24558
rect 12512 24531 13471 24558
rect 13527 24539 13985 24587
rect 14041 24587 15676 24595
rect 14041 24539 15162 24587
rect 13527 24531 15162 24539
rect 15218 24539 15676 24587
rect 15732 24564 28672 24595
rect 15732 24539 23957 24564
rect 15218 24531 23957 24539
rect 12512 24508 23957 24531
rect 24013 24508 24471 24564
rect 24527 24508 25647 24564
rect 25703 24508 26161 24564
rect 26217 24508 27338 24564
rect 27394 24508 27852 24564
rect 27908 24508 28672 24564
rect 12512 24502 28672 24508
rect 1393 24378 28672 24502
rect 1393 24369 6606 24378
rect 1393 24340 6092 24369
rect 1393 24284 1815 24340
rect 1871 24284 2267 24340
rect 2323 24284 2550 24340
rect 2606 24284 2833 24340
rect 2889 24284 3285 24340
rect 3341 24284 3607 24340
rect 3663 24284 4059 24340
rect 4115 24284 4342 24340
rect 4398 24284 4625 24340
rect 4681 24284 5077 24340
rect 5133 24313 6092 24340
rect 6148 24322 6606 24369
rect 6662 24369 8297 24378
rect 6662 24322 7783 24369
rect 6148 24313 7783 24322
rect 7839 24322 8297 24369
rect 8353 24369 13985 24378
rect 8353 24340 13471 24369
rect 8353 24322 9194 24340
rect 7839 24313 9194 24322
rect 5133 24284 9194 24313
rect 9250 24284 9646 24340
rect 9702 24284 9929 24340
rect 9985 24284 10212 24340
rect 10268 24284 10664 24340
rect 10720 24284 10986 24340
rect 11042 24284 11438 24340
rect 11494 24284 11721 24340
rect 11777 24284 12004 24340
rect 12060 24284 12456 24340
rect 12512 24313 13471 24340
rect 13527 24322 13985 24369
rect 14041 24369 15676 24378
rect 14041 24322 15162 24369
rect 13527 24313 15162 24322
rect 15218 24322 15676 24369
rect 15732 24346 28672 24378
rect 15732 24322 23957 24346
rect 15218 24313 23957 24322
rect 12512 24290 23957 24313
rect 24013 24290 24471 24346
rect 24527 24290 25647 24346
rect 25703 24290 26161 24346
rect 26217 24290 27338 24346
rect 27394 24290 27852 24346
rect 27908 24290 28672 24346
rect 12512 24284 28672 24290
rect 1393 24182 28672 24284
rect 1393 24160 16927 24182
rect 1393 24152 6606 24160
rect 1393 24123 6092 24152
rect 1393 24067 1815 24123
rect 1871 24067 2267 24123
rect 2323 24067 2550 24123
rect 2606 24067 2833 24123
rect 2889 24067 3285 24123
rect 3341 24067 3607 24123
rect 3663 24067 4059 24123
rect 4115 24067 4342 24123
rect 4398 24067 4625 24123
rect 4681 24067 5077 24123
rect 5133 24096 6092 24123
rect 6148 24104 6606 24152
rect 6662 24152 8297 24160
rect 6662 24104 7783 24152
rect 6148 24096 7783 24104
rect 7839 24104 8297 24152
rect 8353 24152 13985 24160
rect 8353 24123 13471 24152
rect 8353 24104 9194 24123
rect 7839 24096 9194 24104
rect 5133 24067 9194 24096
rect 9250 24067 9646 24123
rect 9702 24067 9929 24123
rect 9985 24067 10212 24123
rect 10268 24067 10664 24123
rect 10720 24067 10986 24123
rect 11042 24067 11438 24123
rect 11494 24067 11721 24123
rect 11777 24067 12004 24123
rect 12060 24067 12456 24123
rect 12512 24096 13471 24123
rect 13527 24104 13985 24152
rect 14041 24152 15676 24160
rect 14041 24104 15162 24152
rect 13527 24096 15162 24104
rect 15218 24104 15676 24152
rect 15732 24126 16927 24160
rect 16983 24126 17371 24182
rect 17427 24126 17815 24182
rect 17871 24126 18561 24182
rect 18617 24126 19005 24182
rect 19061 24126 19449 24182
rect 19505 24126 20194 24182
rect 20250 24126 20638 24182
rect 20694 24126 21082 24182
rect 21138 24126 21828 24182
rect 21884 24126 22272 24182
rect 22328 24126 22716 24182
rect 22772 24128 28672 24182
rect 22772 24126 23957 24128
rect 15732 24104 23957 24126
rect 15218 24096 23957 24104
rect 12512 24072 23957 24096
rect 24013 24072 24471 24128
rect 24527 24072 25647 24128
rect 25703 24072 26161 24128
rect 26217 24072 27338 24128
rect 27394 24072 27852 24128
rect 27908 24072 28672 24128
rect 12512 24067 28672 24072
rect 1393 23964 28672 24067
rect 1393 23942 16927 23964
rect 1393 23934 6606 23942
rect 1393 23905 6092 23934
rect 1393 23849 1815 23905
rect 1871 23849 2267 23905
rect 2323 23849 2550 23905
rect 2606 23849 2833 23905
rect 2889 23849 3285 23905
rect 3341 23849 3607 23905
rect 3663 23849 4059 23905
rect 4115 23849 4342 23905
rect 4398 23849 4625 23905
rect 4681 23849 5077 23905
rect 5133 23878 6092 23905
rect 6148 23886 6606 23934
rect 6662 23934 8297 23942
rect 6662 23886 7783 23934
rect 6148 23878 7783 23886
rect 7839 23886 8297 23934
rect 8353 23934 13985 23942
rect 8353 23905 13471 23934
rect 8353 23886 9194 23905
rect 7839 23878 9194 23886
rect 5133 23849 9194 23878
rect 9250 23849 9646 23905
rect 9702 23849 9929 23905
rect 9985 23849 10212 23905
rect 10268 23849 10664 23905
rect 10720 23849 10986 23905
rect 11042 23849 11438 23905
rect 11494 23849 11721 23905
rect 11777 23849 12004 23905
rect 12060 23849 12456 23905
rect 12512 23878 13471 23905
rect 13527 23886 13985 23934
rect 14041 23934 15676 23942
rect 14041 23886 15162 23934
rect 13527 23878 15162 23886
rect 15218 23886 15676 23934
rect 15732 23908 16927 23942
rect 16983 23908 17371 23964
rect 17427 23908 17815 23964
rect 17871 23908 18561 23964
rect 18617 23908 19005 23964
rect 19061 23908 19449 23964
rect 19505 23908 20194 23964
rect 20250 23908 20638 23964
rect 20694 23908 21082 23964
rect 21138 23908 21828 23964
rect 21884 23908 22272 23964
rect 22328 23908 22716 23964
rect 22772 23911 28672 23964
rect 22772 23908 23957 23911
rect 15732 23886 23957 23908
rect 15218 23878 23957 23886
rect 12512 23855 23957 23878
rect 24013 23855 24471 23911
rect 24527 23855 25647 23911
rect 25703 23855 26161 23911
rect 26217 23855 27338 23911
rect 27394 23855 27852 23911
rect 27908 23855 28672 23911
rect 12512 23849 28672 23855
rect 1393 23747 28672 23849
rect 1393 23724 16927 23747
rect 1393 23716 6606 23724
rect 1393 23687 6092 23716
rect 1393 23631 1815 23687
rect 1871 23631 2267 23687
rect 2323 23631 2550 23687
rect 2606 23631 2833 23687
rect 2889 23631 3285 23687
rect 3341 23631 3607 23687
rect 3663 23631 4059 23687
rect 4115 23631 4342 23687
rect 4398 23631 4625 23687
rect 4681 23631 5077 23687
rect 5133 23660 6092 23687
rect 6148 23668 6606 23716
rect 6662 23716 8297 23724
rect 6662 23668 7783 23716
rect 6148 23660 7783 23668
rect 7839 23668 8297 23716
rect 8353 23716 13985 23724
rect 8353 23687 13471 23716
rect 8353 23668 9194 23687
rect 7839 23660 9194 23668
rect 5133 23631 9194 23660
rect 9250 23631 9646 23687
rect 9702 23631 9929 23687
rect 9985 23631 10212 23687
rect 10268 23631 10664 23687
rect 10720 23631 10986 23687
rect 11042 23631 11438 23687
rect 11494 23631 11721 23687
rect 11777 23631 12004 23687
rect 12060 23631 12456 23687
rect 12512 23660 13471 23687
rect 13527 23668 13985 23716
rect 14041 23716 15676 23724
rect 14041 23668 15162 23716
rect 13527 23660 15162 23668
rect 15218 23668 15676 23716
rect 15732 23691 16927 23724
rect 16983 23691 17371 23747
rect 17427 23691 17815 23747
rect 17871 23691 18561 23747
rect 18617 23691 19005 23747
rect 19061 23691 19449 23747
rect 19505 23691 20194 23747
rect 20250 23691 20638 23747
rect 20694 23691 21082 23747
rect 21138 23691 21828 23747
rect 21884 23691 22272 23747
rect 22328 23691 22716 23747
rect 22772 23691 28672 23747
rect 15732 23668 28672 23691
rect 15218 23660 28672 23668
rect 12512 23631 28672 23660
rect 1393 23529 28672 23631
rect 1393 23507 16927 23529
rect 1393 23498 6606 23507
rect 1393 23469 6092 23498
rect 1393 23413 1815 23469
rect 1871 23413 2267 23469
rect 2323 23413 2550 23469
rect 2606 23413 2833 23469
rect 2889 23413 3285 23469
rect 3341 23413 3607 23469
rect 3663 23413 4059 23469
rect 4115 23413 4342 23469
rect 4398 23413 4625 23469
rect 4681 23413 5077 23469
rect 5133 23442 6092 23469
rect 6148 23451 6606 23498
rect 6662 23498 8297 23507
rect 6662 23451 7783 23498
rect 6148 23442 7783 23451
rect 7839 23451 8297 23498
rect 8353 23498 13985 23507
rect 8353 23469 13471 23498
rect 8353 23451 9194 23469
rect 7839 23442 9194 23451
rect 5133 23413 9194 23442
rect 9250 23413 9646 23469
rect 9702 23413 9929 23469
rect 9985 23413 10212 23469
rect 10268 23413 10664 23469
rect 10720 23413 10986 23469
rect 11042 23413 11438 23469
rect 11494 23413 11721 23469
rect 11777 23413 12004 23469
rect 12060 23413 12456 23469
rect 12512 23442 13471 23469
rect 13527 23451 13985 23498
rect 14041 23498 15676 23507
rect 14041 23451 15162 23498
rect 13527 23442 15162 23451
rect 15218 23451 15676 23498
rect 15732 23473 16927 23507
rect 16983 23473 17371 23529
rect 17427 23473 17815 23529
rect 17871 23473 18561 23529
rect 18617 23473 19005 23529
rect 19061 23473 19449 23529
rect 19505 23473 20194 23529
rect 20250 23473 20638 23529
rect 20694 23473 21082 23529
rect 21138 23473 21828 23529
rect 21884 23473 22272 23529
rect 22328 23473 22716 23529
rect 22772 23473 28672 23529
rect 15732 23451 28672 23473
rect 15218 23442 28672 23451
rect 12512 23413 28672 23442
rect 1393 23311 28672 23413
rect 1393 23289 16927 23311
rect 1393 23281 6606 23289
rect 1393 23252 6092 23281
rect 1393 23196 1815 23252
rect 1871 23196 2267 23252
rect 2323 23196 2550 23252
rect 2606 23196 2833 23252
rect 2889 23196 3285 23252
rect 3341 23196 3607 23252
rect 3663 23196 4059 23252
rect 4115 23196 4342 23252
rect 4398 23196 4625 23252
rect 4681 23196 5077 23252
rect 5133 23225 6092 23252
rect 6148 23233 6606 23281
rect 6662 23281 8297 23289
rect 6662 23233 7783 23281
rect 6148 23225 7783 23233
rect 7839 23233 8297 23281
rect 8353 23281 13985 23289
rect 8353 23252 13471 23281
rect 8353 23233 9194 23252
rect 7839 23225 9194 23233
rect 5133 23196 9194 23225
rect 9250 23196 9646 23252
rect 9702 23196 9929 23252
rect 9985 23196 10212 23252
rect 10268 23196 10664 23252
rect 10720 23196 10986 23252
rect 11042 23196 11438 23252
rect 11494 23196 11721 23252
rect 11777 23196 12004 23252
rect 12060 23196 12456 23252
rect 12512 23225 13471 23252
rect 13527 23233 13985 23281
rect 14041 23281 15676 23289
rect 14041 23233 15162 23281
rect 13527 23225 15162 23233
rect 15218 23233 15676 23281
rect 15732 23255 16927 23289
rect 16983 23255 17371 23311
rect 17427 23255 17815 23311
rect 17871 23255 18561 23311
rect 18617 23255 19005 23311
rect 19061 23255 19449 23311
rect 19505 23255 20194 23311
rect 20250 23255 20638 23311
rect 20694 23255 21082 23311
rect 21138 23255 21828 23311
rect 21884 23255 22272 23311
rect 22328 23255 22716 23311
rect 22772 23255 28672 23311
rect 15732 23233 28672 23255
rect 15218 23225 28672 23233
rect 12512 23196 28672 23225
rect 1393 23094 28672 23196
rect 1393 23063 16927 23094
rect 1393 23034 6092 23063
rect 1393 22978 1815 23034
rect 1871 22978 2267 23034
rect 2323 22978 2550 23034
rect 2606 22978 2833 23034
rect 2889 22978 3285 23034
rect 3341 22978 3607 23034
rect 3663 22978 4059 23034
rect 4115 22978 4342 23034
rect 4398 22978 4625 23034
rect 4681 22978 5077 23034
rect 5133 23007 6092 23034
rect 6148 23007 7783 23063
rect 7839 23034 13471 23063
rect 7839 23007 9194 23034
rect 5133 22978 9194 23007
rect 9250 22978 9646 23034
rect 9702 22978 9929 23034
rect 9985 22978 10212 23034
rect 10268 22978 10664 23034
rect 10720 22978 10986 23034
rect 11042 22978 11438 23034
rect 11494 22978 11721 23034
rect 11777 22978 12004 23034
rect 12060 22978 12456 23034
rect 12512 23007 13471 23034
rect 13527 23007 15162 23063
rect 15218 23038 16927 23063
rect 16983 23038 17371 23094
rect 17427 23038 17815 23094
rect 17871 23038 18561 23094
rect 18617 23038 19005 23094
rect 19061 23038 19449 23094
rect 19505 23038 20194 23094
rect 20250 23038 20638 23094
rect 20694 23038 21082 23094
rect 21138 23038 21828 23094
rect 21884 23038 22272 23094
rect 22328 23038 22716 23094
rect 22772 23038 28672 23094
rect 15218 23007 28672 23038
rect 12512 22978 28672 23007
rect 1393 22876 28672 22978
rect 1393 22846 16927 22876
rect 1393 22817 6092 22846
rect 1393 22761 1815 22817
rect 1871 22761 2267 22817
rect 2323 22761 2550 22817
rect 2606 22761 2833 22817
rect 2889 22761 3285 22817
rect 3341 22761 3607 22817
rect 3663 22761 4059 22817
rect 4115 22761 4342 22817
rect 4398 22761 4625 22817
rect 4681 22761 5077 22817
rect 5133 22790 6092 22817
rect 6148 22790 7783 22846
rect 7839 22817 13471 22846
rect 7839 22790 9194 22817
rect 5133 22761 9194 22790
rect 9250 22761 9646 22817
rect 9702 22761 9929 22817
rect 9985 22761 10212 22817
rect 10268 22761 10664 22817
rect 10720 22761 10986 22817
rect 11042 22761 11438 22817
rect 11494 22761 11721 22817
rect 11777 22761 12004 22817
rect 12060 22761 12456 22817
rect 12512 22790 13471 22817
rect 13527 22790 15162 22846
rect 15218 22820 16927 22846
rect 16983 22820 17371 22876
rect 17427 22820 17815 22876
rect 17871 22820 18561 22876
rect 18617 22820 19005 22876
rect 19061 22820 19449 22876
rect 19505 22820 20194 22876
rect 20250 22820 20638 22876
rect 20694 22820 21082 22876
rect 21138 22820 21828 22876
rect 21884 22820 22272 22876
rect 22328 22820 22716 22876
rect 22772 22820 28672 22876
rect 15218 22790 28672 22820
rect 12512 22761 28672 22790
rect 1393 22671 28672 22761
rect 24915 22446 25041 22485
rect 24915 22390 24950 22446
rect 25006 22390 25041 22446
rect 24915 22376 25041 22390
rect 26605 22446 26731 22485
rect 26605 22390 26640 22446
rect 26696 22390 26731 22446
rect 26605 22376 26731 22390
rect 28296 22446 28422 22485
rect 28296 22390 28331 22446
rect 28387 22390 28422 22446
rect 28296 22376 28422 22390
rect 23286 22243 28423 22376
rect 24915 22228 25041 22243
rect 24915 22172 24950 22228
rect 25006 22172 25041 22228
rect 24915 22133 25041 22172
rect 26605 22228 26731 22243
rect 26605 22172 26640 22228
rect 26696 22172 26731 22228
rect 26605 22133 26731 22172
rect 28296 22228 28422 22243
rect 28296 22172 28331 22228
rect 28387 22172 28422 22228
rect 28296 22133 28422 22172
rect 7050 22043 7176 22082
rect 7050 21987 7085 22043
rect 7141 21987 7176 22043
rect 7050 21973 7176 21987
rect 8741 22043 8867 22082
rect 8741 21987 8776 22043
rect 8832 21987 8867 22043
rect 8741 21973 8867 21987
rect 14429 22043 14555 22082
rect 14429 21987 14464 22043
rect 14520 21987 14555 22043
rect 14429 21973 14555 21987
rect 16120 22043 16246 22082
rect 16120 21987 16155 22043
rect 16211 21987 16246 22043
rect 16120 21973 16246 21987
rect 5421 21839 8868 21973
rect 12800 21839 16247 21973
rect 23294 21970 28476 22009
rect 23294 21914 24460 21970
rect 24516 21914 26150 21970
rect 26206 21914 27841 21970
rect 27897 21914 28476 21970
rect 23294 21876 28476 21914
rect 24424 21875 24552 21876
rect 26114 21875 26242 21876
rect 27805 21875 27933 21876
rect 7050 21825 7176 21839
rect 7050 21769 7085 21825
rect 7141 21769 7176 21825
rect 7050 21730 7176 21769
rect 8741 21825 8867 21839
rect 8741 21769 8776 21825
rect 8832 21769 8867 21825
rect 8741 21730 8867 21769
rect 14429 21825 14555 21839
rect 14429 21769 14464 21825
rect 14520 21769 14555 21825
rect 14429 21730 14555 21769
rect 16120 21825 16246 21839
rect 16120 21769 16155 21825
rect 16211 21769 16246 21825
rect 16120 21730 16246 21769
rect 24425 21752 24551 21875
rect 24425 21696 24460 21752
rect 24516 21696 24551 21752
rect 24425 21657 24551 21696
rect 26115 21752 26241 21875
rect 26115 21696 26150 21752
rect 26206 21696 26241 21752
rect 26115 21657 26241 21696
rect 27806 21752 27932 21875
rect 27806 21696 27841 21752
rect 27897 21696 27932 21752
rect 27806 21657 27932 21696
rect 6560 21605 6686 21606
rect 8251 21605 8377 21606
rect 13939 21605 14065 21606
rect 15630 21605 15756 21606
rect 5430 21567 8921 21605
rect 5430 21511 6595 21567
rect 6651 21511 8286 21567
rect 8342 21511 8921 21567
rect 5430 21472 8921 21511
rect 12809 21567 16300 21605
rect 12809 21511 13974 21567
rect 14030 21511 15665 21567
rect 15721 21511 16300 21567
rect 12809 21472 16300 21511
rect 6560 21349 6686 21472
rect 6560 21293 6595 21349
rect 6651 21293 6686 21349
rect 6560 21254 6686 21293
rect 8251 21349 8377 21472
rect 8251 21293 8286 21349
rect 8342 21293 8377 21349
rect 8251 21254 8377 21293
rect 13939 21349 14065 21472
rect 13939 21293 13974 21349
rect 14030 21293 14065 21349
rect 13939 21254 14065 21293
rect 15630 21349 15756 21472
rect 15630 21293 15665 21349
rect 15721 21293 15756 21349
rect 15630 21254 15756 21293
rect 2096 20387 28424 20497
rect 2096 20366 17371 20387
rect 2096 20310 2267 20366
rect 2323 20310 2550 20366
rect 2606 20310 2833 20366
rect 2889 20310 4059 20366
rect 4115 20310 4342 20366
rect 4398 20310 4625 20366
rect 4681 20310 9646 20366
rect 9702 20310 9929 20366
rect 9985 20310 10212 20366
rect 10268 20310 11438 20366
rect 11494 20310 11721 20366
rect 11777 20310 12004 20366
rect 12060 20331 17371 20366
rect 17427 20331 19005 20387
rect 19061 20331 20638 20387
rect 20694 20331 22272 20387
rect 22328 20331 28424 20387
rect 12060 20310 28424 20331
rect 2096 20169 28424 20310
rect 2096 20148 17371 20169
rect 2096 20092 2267 20148
rect 2323 20092 2550 20148
rect 2606 20092 2833 20148
rect 2889 20092 4059 20148
rect 4115 20092 4342 20148
rect 4398 20092 4625 20148
rect 4681 20092 9646 20148
rect 9702 20092 9929 20148
rect 9985 20092 10212 20148
rect 10268 20092 11438 20148
rect 11494 20092 11721 20148
rect 11777 20092 12004 20148
rect 12060 20113 17371 20148
rect 17427 20113 19005 20169
rect 19061 20113 20638 20169
rect 20694 20113 22272 20169
rect 22328 20113 28424 20169
rect 12060 20092 28424 20113
rect 2096 19951 28424 20092
rect 2096 19930 17371 19951
rect 2096 19874 2267 19930
rect 2323 19874 2550 19930
rect 2606 19874 2833 19930
rect 2889 19874 4059 19930
rect 4115 19874 4342 19930
rect 4398 19874 4625 19930
rect 4681 19874 9646 19930
rect 9702 19874 9929 19930
rect 9985 19874 10212 19930
rect 10268 19874 11438 19930
rect 11494 19874 11721 19930
rect 11777 19874 12004 19930
rect 12060 19895 17371 19930
rect 17427 19895 19005 19951
rect 19061 19895 20638 19951
rect 20694 19895 22272 19951
rect 22328 19895 28424 19951
rect 12060 19874 28424 19895
rect 2096 19815 28424 19874
rect 2096 18659 28424 19567
rect 2096 18428 23261 18488
rect 2096 18408 17371 18428
rect 2096 18352 2267 18408
rect 2323 18352 2550 18408
rect 2606 18352 2833 18408
rect 2889 18352 4059 18408
rect 4115 18352 4342 18408
rect 4398 18352 4625 18408
rect 4681 18352 9646 18408
rect 9702 18352 9929 18408
rect 9985 18352 10212 18408
rect 10268 18352 11438 18408
rect 11494 18352 11721 18408
rect 11777 18352 12004 18408
rect 12060 18372 17371 18408
rect 17427 18372 19005 18428
rect 19061 18372 20638 18428
rect 20694 18372 22272 18428
rect 22328 18372 23261 18428
rect 12060 18352 23261 18372
rect 2096 18210 23261 18352
rect 2096 18190 17371 18210
rect 2096 18134 2267 18190
rect 2323 18134 2550 18190
rect 2606 18134 2833 18190
rect 2889 18134 4059 18190
rect 4115 18134 4342 18190
rect 4398 18134 4625 18190
rect 4681 18134 9646 18190
rect 9702 18134 9929 18190
rect 9985 18134 10212 18190
rect 10268 18134 11438 18190
rect 11494 18134 11721 18190
rect 11777 18134 12004 18190
rect 12060 18154 17371 18190
rect 17427 18154 19005 18210
rect 19061 18154 20638 18210
rect 20694 18154 22272 18210
rect 22328 18154 23261 18210
rect 12060 18134 23261 18154
rect 2096 17992 23261 18134
rect 28189 18104 28318 18237
rect 2096 17972 17371 17992
rect 2096 17916 2267 17972
rect 2323 17916 2550 17972
rect 2606 17916 2833 17972
rect 2889 17916 4059 17972
rect 4115 17916 4342 17972
rect 4398 17916 4625 17972
rect 4681 17916 9646 17972
rect 9702 17916 9929 17972
rect 9985 17916 10212 17972
rect 10268 17916 11438 17972
rect 11494 17916 11721 17972
rect 11777 17916 12004 17972
rect 12060 17936 17371 17972
rect 17427 17936 19005 17992
rect 19061 17936 20638 17992
rect 20694 17936 22272 17992
rect 22328 17936 23261 17992
rect 12060 17916 23261 17936
rect 2096 17774 23261 17916
rect 2096 17754 17371 17774
rect 2096 17698 2267 17754
rect 2323 17698 2550 17754
rect 2606 17698 2833 17754
rect 2889 17698 4059 17754
rect 4115 17698 4342 17754
rect 4398 17698 4625 17754
rect 4681 17698 9646 17754
rect 9702 17698 9929 17754
rect 9985 17698 10212 17754
rect 10268 17698 11438 17754
rect 11494 17698 11721 17754
rect 11777 17698 12004 17754
rect 12060 17718 17371 17754
rect 17427 17718 19005 17774
rect 19061 17718 20638 17774
rect 20694 17718 22272 17774
rect 22328 17718 23261 17774
rect 12060 17698 23261 17718
rect 2096 17580 23261 17698
rect 1988 16914 20547 16996
rect 1980 16904 20547 16914
rect 1980 16848 1990 16904
rect 2046 16848 2662 16904
rect 2718 16848 3110 16904
rect 3166 16848 3782 16904
rect 3838 16848 4230 16904
rect 4286 16848 4902 16904
rect 4958 16848 5350 16904
rect 5406 16848 6022 16904
rect 6078 16848 6470 16904
rect 6526 16848 7142 16904
rect 7198 16848 7590 16904
rect 7646 16848 8262 16904
rect 8318 16848 8710 16904
rect 8766 16848 9382 16904
rect 9438 16848 9830 16904
rect 9886 16848 10502 16904
rect 10558 16848 10950 16904
rect 11006 16848 11622 16904
rect 11678 16848 12070 16904
rect 12126 16848 12742 16904
rect 12798 16848 13190 16904
rect 13246 16848 13862 16904
rect 13918 16848 14310 16904
rect 14366 16848 14982 16904
rect 15038 16848 15430 16904
rect 15486 16848 16102 16904
rect 16158 16848 16550 16904
rect 16606 16848 17222 16904
rect 17278 16848 17670 16904
rect 17726 16848 18342 16904
rect 18398 16848 18790 16904
rect 18846 16848 19462 16904
rect 19518 16848 19910 16904
rect 19966 16848 20547 16904
rect 1980 16780 20547 16848
rect 1980 16724 1990 16780
rect 2046 16724 2662 16780
rect 2718 16724 3110 16780
rect 3166 16724 3782 16780
rect 3838 16724 4230 16780
rect 4286 16724 4902 16780
rect 4958 16724 5350 16780
rect 5406 16724 6022 16780
rect 6078 16724 6470 16780
rect 6526 16724 7142 16780
rect 7198 16724 7590 16780
rect 7646 16724 8262 16780
rect 8318 16724 8710 16780
rect 8766 16724 9382 16780
rect 9438 16724 9830 16780
rect 9886 16724 10502 16780
rect 10558 16724 10950 16780
rect 11006 16724 11622 16780
rect 11678 16724 12070 16780
rect 12126 16724 12742 16780
rect 12798 16724 13190 16780
rect 13246 16724 13862 16780
rect 13918 16724 14310 16780
rect 14366 16724 14982 16780
rect 15038 16724 15430 16780
rect 15486 16724 16102 16780
rect 16158 16724 16550 16780
rect 16606 16724 17222 16780
rect 17278 16724 17670 16780
rect 17726 16724 18342 16780
rect 18398 16724 18790 16780
rect 18846 16724 19462 16780
rect 19518 16724 19910 16780
rect 19966 16724 20547 16780
rect 1980 16656 20547 16724
rect 1980 16600 1990 16656
rect 2046 16600 2662 16656
rect 2718 16600 3110 16656
rect 3166 16600 3782 16656
rect 3838 16600 4230 16656
rect 4286 16600 4902 16656
rect 4958 16600 5350 16656
rect 5406 16600 6022 16656
rect 6078 16600 6470 16656
rect 6526 16600 7142 16656
rect 7198 16600 7590 16656
rect 7646 16600 8262 16656
rect 8318 16600 8710 16656
rect 8766 16600 9382 16656
rect 9438 16600 9830 16656
rect 9886 16600 10502 16656
rect 10558 16600 10950 16656
rect 11006 16600 11622 16656
rect 11678 16600 12070 16656
rect 12126 16600 12742 16656
rect 12798 16600 13190 16656
rect 13246 16600 13862 16656
rect 13918 16600 14310 16656
rect 14366 16600 14982 16656
rect 15038 16600 15430 16656
rect 15486 16600 16102 16656
rect 16158 16600 16550 16656
rect 16606 16600 17222 16656
rect 17278 16600 17670 16656
rect 17726 16600 18342 16656
rect 18398 16600 18790 16656
rect 18846 16600 19462 16656
rect 19518 16600 19910 16656
rect 19966 16600 20547 16656
rect 1980 16532 20547 16600
rect 1980 16476 1990 16532
rect 2046 16476 2662 16532
rect 2718 16476 3110 16532
rect 3166 16476 3782 16532
rect 3838 16476 4230 16532
rect 4286 16476 4902 16532
rect 4958 16476 5350 16532
rect 5406 16476 6022 16532
rect 6078 16476 6470 16532
rect 6526 16476 7142 16532
rect 7198 16476 7590 16532
rect 7646 16476 8262 16532
rect 8318 16476 8710 16532
rect 8766 16476 9382 16532
rect 9438 16476 9830 16532
rect 9886 16476 10502 16532
rect 10558 16476 10950 16532
rect 11006 16476 11622 16532
rect 11678 16476 12070 16532
rect 12126 16476 12742 16532
rect 12798 16476 13190 16532
rect 13246 16476 13862 16532
rect 13918 16476 14310 16532
rect 14366 16476 14982 16532
rect 15038 16476 15430 16532
rect 15486 16476 16102 16532
rect 16158 16476 16550 16532
rect 16606 16476 17222 16532
rect 17278 16476 17670 16532
rect 17726 16476 18342 16532
rect 18398 16476 18790 16532
rect 18846 16476 19462 16532
rect 19518 16476 19910 16532
rect 19966 16476 20547 16532
rect 1980 16408 20547 16476
rect 1980 16352 1990 16408
rect 2046 16352 2662 16408
rect 2718 16352 3110 16408
rect 3166 16352 3782 16408
rect 3838 16352 4230 16408
rect 4286 16352 4902 16408
rect 4958 16352 5350 16408
rect 5406 16352 6022 16408
rect 6078 16352 6470 16408
rect 6526 16352 7142 16408
rect 7198 16352 7590 16408
rect 7646 16352 8262 16408
rect 8318 16352 8710 16408
rect 8766 16352 9382 16408
rect 9438 16352 9830 16408
rect 9886 16352 10502 16408
rect 10558 16352 10950 16408
rect 11006 16352 11622 16408
rect 11678 16352 12070 16408
rect 12126 16352 12742 16408
rect 12798 16352 13190 16408
rect 13246 16352 13862 16408
rect 13918 16352 14310 16408
rect 14366 16352 14982 16408
rect 15038 16352 15430 16408
rect 15486 16352 16102 16408
rect 16158 16352 16550 16408
rect 16606 16352 17222 16408
rect 17278 16352 17670 16408
rect 17726 16352 18342 16408
rect 18398 16352 18790 16408
rect 18846 16352 19462 16408
rect 19518 16352 19910 16408
rect 19966 16352 20547 16408
rect 1980 16284 20547 16352
rect 1980 16228 1990 16284
rect 2046 16228 2662 16284
rect 2718 16228 3110 16284
rect 3166 16228 3782 16284
rect 3838 16228 4230 16284
rect 4286 16228 4902 16284
rect 4958 16228 5350 16284
rect 5406 16228 6022 16284
rect 6078 16228 6470 16284
rect 6526 16228 7142 16284
rect 7198 16228 7590 16284
rect 7646 16228 8262 16284
rect 8318 16228 8710 16284
rect 8766 16228 9382 16284
rect 9438 16228 9830 16284
rect 9886 16228 10502 16284
rect 10558 16228 10950 16284
rect 11006 16228 11622 16284
rect 11678 16228 12070 16284
rect 12126 16228 12742 16284
rect 12798 16228 13190 16284
rect 13246 16228 13862 16284
rect 13918 16228 14310 16284
rect 14366 16228 14982 16284
rect 15038 16228 15430 16284
rect 15486 16228 16102 16284
rect 16158 16228 16550 16284
rect 16606 16228 17222 16284
rect 17278 16228 17670 16284
rect 17726 16228 18342 16284
rect 18398 16228 18790 16284
rect 18846 16228 19462 16284
rect 19518 16228 19910 16284
rect 19966 16228 20547 16284
rect 1980 16160 20547 16228
rect 1980 16104 1990 16160
rect 2046 16104 2662 16160
rect 2718 16104 3110 16160
rect 3166 16104 3782 16160
rect 3838 16104 4230 16160
rect 4286 16104 4902 16160
rect 4958 16104 5350 16160
rect 5406 16104 6022 16160
rect 6078 16104 6470 16160
rect 6526 16104 7142 16160
rect 7198 16104 7590 16160
rect 7646 16104 8262 16160
rect 8318 16104 8710 16160
rect 8766 16104 9382 16160
rect 9438 16104 9830 16160
rect 9886 16104 10502 16160
rect 10558 16104 10950 16160
rect 11006 16104 11622 16160
rect 11678 16104 12070 16160
rect 12126 16104 12742 16160
rect 12798 16104 13190 16160
rect 13246 16104 13862 16160
rect 13918 16104 14310 16160
rect 14366 16104 14982 16160
rect 15038 16104 15430 16160
rect 15486 16104 16102 16160
rect 16158 16104 16550 16160
rect 16606 16104 17222 16160
rect 17278 16104 17670 16160
rect 17726 16104 18342 16160
rect 18398 16104 18790 16160
rect 18846 16104 19462 16160
rect 19518 16104 19910 16160
rect 19966 16104 20547 16160
rect 1980 16036 20547 16104
rect 1980 15980 1990 16036
rect 2046 15980 2662 16036
rect 2718 15980 3110 16036
rect 3166 15980 3782 16036
rect 3838 15980 4230 16036
rect 4286 15980 4902 16036
rect 4958 15980 5350 16036
rect 5406 15980 6022 16036
rect 6078 15980 6470 16036
rect 6526 15980 7142 16036
rect 7198 15980 7590 16036
rect 7646 15980 8262 16036
rect 8318 15980 8710 16036
rect 8766 15980 9382 16036
rect 9438 15980 9830 16036
rect 9886 15980 10502 16036
rect 10558 15980 10950 16036
rect 11006 15980 11622 16036
rect 11678 15980 12070 16036
rect 12126 15980 12742 16036
rect 12798 15980 13190 16036
rect 13246 15980 13862 16036
rect 13918 15980 14310 16036
rect 14366 15980 14982 16036
rect 15038 15980 15430 16036
rect 15486 15980 16102 16036
rect 16158 15980 16550 16036
rect 16606 15980 17222 16036
rect 17278 15980 17670 16036
rect 17726 15980 18342 16036
rect 18398 15980 18790 16036
rect 18846 15980 19462 16036
rect 19518 15980 19910 16036
rect 19966 15980 20547 16036
rect 1980 15912 20547 15980
rect 1980 15856 1990 15912
rect 2046 15856 2662 15912
rect 2718 15856 3110 15912
rect 3166 15856 3782 15912
rect 3838 15856 4230 15912
rect 4286 15856 4902 15912
rect 4958 15856 5350 15912
rect 5406 15856 6022 15912
rect 6078 15856 6470 15912
rect 6526 15856 7142 15912
rect 7198 15856 7590 15912
rect 7646 15856 8262 15912
rect 8318 15856 8710 15912
rect 8766 15856 9382 15912
rect 9438 15856 9830 15912
rect 9886 15856 10502 15912
rect 10558 15856 10950 15912
rect 11006 15856 11622 15912
rect 11678 15856 12070 15912
rect 12126 15856 12742 15912
rect 12798 15856 13190 15912
rect 13246 15856 13862 15912
rect 13918 15856 14310 15912
rect 14366 15856 14982 15912
rect 15038 15856 15430 15912
rect 15486 15856 16102 15912
rect 16158 15856 16550 15912
rect 16606 15856 17222 15912
rect 17278 15856 17670 15912
rect 17726 15856 18342 15912
rect 18398 15856 18790 15912
rect 18846 15856 19462 15912
rect 19518 15856 19910 15912
rect 19966 15856 20547 15912
rect 1980 15788 20547 15856
rect 1980 15732 1990 15788
rect 2046 15732 2662 15788
rect 2718 15732 3110 15788
rect 3166 15732 3782 15788
rect 3838 15732 4230 15788
rect 4286 15732 4902 15788
rect 4958 15732 5350 15788
rect 5406 15732 6022 15788
rect 6078 15732 6470 15788
rect 6526 15732 7142 15788
rect 7198 15732 7590 15788
rect 7646 15732 8262 15788
rect 8318 15732 8710 15788
rect 8766 15732 9382 15788
rect 9438 15732 9830 15788
rect 9886 15732 10502 15788
rect 10558 15732 10950 15788
rect 11006 15732 11622 15788
rect 11678 15732 12070 15788
rect 12126 15732 12742 15788
rect 12798 15732 13190 15788
rect 13246 15732 13862 15788
rect 13918 15732 14310 15788
rect 14366 15732 14982 15788
rect 15038 15732 15430 15788
rect 15486 15732 16102 15788
rect 16158 15732 16550 15788
rect 16606 15732 17222 15788
rect 17278 15732 17670 15788
rect 17726 15732 18342 15788
rect 18398 15732 18790 15788
rect 18846 15732 19462 15788
rect 19518 15732 19910 15788
rect 19966 15732 20547 15788
rect 1980 15664 20547 15732
rect 1980 15608 1990 15664
rect 2046 15608 2662 15664
rect 2718 15608 3110 15664
rect 3166 15608 3782 15664
rect 3838 15608 4230 15664
rect 4286 15608 4902 15664
rect 4958 15608 5350 15664
rect 5406 15608 6022 15664
rect 6078 15608 6470 15664
rect 6526 15608 7142 15664
rect 7198 15608 7590 15664
rect 7646 15608 8262 15664
rect 8318 15608 8710 15664
rect 8766 15608 9382 15664
rect 9438 15608 9830 15664
rect 9886 15608 10502 15664
rect 10558 15608 10950 15664
rect 11006 15608 11622 15664
rect 11678 15608 12070 15664
rect 12126 15608 12742 15664
rect 12798 15608 13190 15664
rect 13246 15608 13862 15664
rect 13918 15608 14310 15664
rect 14366 15608 14982 15664
rect 15038 15608 15430 15664
rect 15486 15608 16102 15664
rect 16158 15608 16550 15664
rect 16606 15608 17222 15664
rect 17278 15608 17670 15664
rect 17726 15608 18342 15664
rect 18398 15608 18790 15664
rect 18846 15608 19462 15664
rect 19518 15608 19910 15664
rect 19966 15608 20547 15664
rect 1980 15540 20547 15608
rect 1980 15484 1990 15540
rect 2046 15484 2662 15540
rect 2718 15484 3110 15540
rect 3166 15484 3782 15540
rect 3838 15484 4230 15540
rect 4286 15484 4902 15540
rect 4958 15484 5350 15540
rect 5406 15484 6022 15540
rect 6078 15484 6470 15540
rect 6526 15484 7142 15540
rect 7198 15484 7590 15540
rect 7646 15484 8262 15540
rect 8318 15484 8710 15540
rect 8766 15484 9382 15540
rect 9438 15484 9830 15540
rect 9886 15484 10502 15540
rect 10558 15484 10950 15540
rect 11006 15484 11622 15540
rect 11678 15484 12070 15540
rect 12126 15484 12742 15540
rect 12798 15484 13190 15540
rect 13246 15484 13862 15540
rect 13918 15484 14310 15540
rect 14366 15484 14982 15540
rect 15038 15484 15430 15540
rect 15486 15484 16102 15540
rect 16158 15484 16550 15540
rect 16606 15484 17222 15540
rect 17278 15484 17670 15540
rect 17726 15484 18342 15540
rect 18398 15484 18790 15540
rect 18846 15484 19462 15540
rect 19518 15484 19910 15540
rect 19966 15484 20547 15540
rect 1980 15474 20547 15484
rect 1988 15258 20547 15474
rect 1740 14934 10818 15020
rect 19201 14973 28239 15020
rect 1740 14878 10277 14934
rect 10333 14878 10725 14934
rect 10781 14878 10818 14934
rect 1740 14791 10818 14878
rect 19200 14934 28239 14973
rect 19200 14878 19237 14934
rect 19293 14878 19685 14934
rect 19741 14878 28239 14934
rect 19200 14839 28239 14878
rect 19201 14791 28239 14839
rect 1740 14594 9700 14680
rect 18081 14633 28239 14680
rect 1740 14538 9158 14594
rect 9214 14538 9605 14594
rect 9661 14538 9700 14594
rect 1740 14451 9700 14538
rect 18080 14594 28239 14633
rect 18080 14538 18117 14594
rect 18173 14538 18565 14594
rect 18621 14538 28239 14594
rect 18080 14499 28239 14538
rect 18081 14451 28239 14499
rect 1740 14292 8578 14340
rect 16961 14292 28239 14340
rect 1740 14253 8579 14292
rect 1740 14197 8038 14253
rect 8094 14197 8486 14253
rect 8542 14197 8579 14253
rect 1740 14158 8579 14197
rect 16960 14253 28239 14292
rect 16960 14197 16997 14253
rect 17053 14197 17445 14253
rect 17501 14197 28239 14253
rect 16960 14158 28239 14197
rect 1740 14111 8578 14158
rect 16961 14111 28239 14158
rect 1740 13952 7458 14000
rect 15841 13952 28239 14000
rect 1740 13913 7459 13952
rect 1740 13857 6918 13913
rect 6974 13857 7366 13913
rect 7422 13857 7459 13913
rect 1740 13818 7459 13857
rect 15840 13913 28239 13952
rect 15840 13857 15877 13913
rect 15933 13857 16325 13913
rect 16381 13857 28239 13913
rect 15840 13818 28239 13857
rect 1740 13771 7458 13818
rect 15841 13771 28239 13818
rect 1740 13612 6338 13660
rect 14721 13612 28239 13660
rect 1740 13573 6339 13612
rect 1740 13517 5798 13573
rect 5854 13517 6246 13573
rect 6302 13517 6339 13573
rect 1740 13478 6339 13517
rect 14720 13573 28239 13612
rect 14720 13517 14757 13573
rect 14813 13517 15205 13573
rect 15261 13517 28239 13573
rect 14720 13478 28239 13517
rect 1740 13431 6338 13478
rect 14721 13431 28239 13478
rect 1740 13272 5218 13320
rect 13601 13272 28239 13320
rect 1740 13233 5219 13272
rect 1740 13177 4678 13233
rect 4734 13177 5126 13233
rect 5182 13177 5219 13233
rect 1740 13138 5219 13177
rect 13600 13233 28239 13272
rect 13600 13177 13637 13233
rect 13693 13177 14085 13233
rect 14141 13177 28239 13233
rect 13600 13138 28239 13177
rect 1740 13091 5218 13138
rect 13601 13091 28239 13138
rect 1740 12932 4098 12980
rect 1740 12893 4099 12932
rect 1740 12837 3558 12893
rect 3614 12837 4006 12893
rect 4062 12837 4099 12893
rect 1740 12798 4099 12837
rect 12479 12893 28239 12980
rect 12479 12837 12517 12893
rect 12573 12837 12965 12893
rect 13021 12837 28239 12893
rect 1740 12751 4098 12798
rect 12479 12751 28239 12837
rect 1740 12592 2978 12640
rect 11361 12592 28239 12640
rect 1740 12553 2979 12592
rect 1740 12497 2438 12553
rect 2494 12497 2886 12553
rect 2942 12497 2979 12553
rect 1740 12458 2979 12497
rect 11360 12553 28239 12592
rect 11360 12497 11397 12553
rect 11453 12497 11845 12553
rect 11901 12497 28239 12553
rect 11360 12458 28239 12497
rect 1740 12411 2978 12458
rect 11361 12411 28239 12458
rect 1970 12152 2096 12191
rect 1970 12096 2005 12152
rect 2061 12096 2096 12152
rect 12706 12168 12832 12207
rect 12706 12112 12741 12168
rect 12797 12112 12832 12168
rect 1970 12077 2096 12096
rect 10928 12077 11268 12098
rect 12706 12077 12832 12112
rect 1970 12059 12834 12077
rect 1970 12003 10964 12059
rect 11020 12003 11176 12059
rect 11232 12003 12834 12059
rect 1970 11985 12834 12003
rect 1970 11934 2096 11985
rect 10928 11964 11268 11985
rect 1970 11878 2005 11934
rect 2061 11878 2096 11934
rect 12706 11950 12832 11985
rect 12706 11894 12741 11950
rect 12797 11894 12832 11950
rect 1970 11839 2096 11878
rect 3089 11869 3429 11889
rect 12048 11869 12388 11889
rect 3089 11850 12388 11869
rect 12706 11855 12832 11894
rect 3089 11794 3125 11850
rect 3181 11794 3337 11850
rect 3393 11794 12084 11850
rect 12140 11794 12296 11850
rect 12352 11794 12388 11850
rect 3089 11776 12388 11794
rect 3089 11755 3429 11776
rect 12048 11755 12388 11776
rect 4210 11660 4336 11661
rect 11582 11660 11712 11681
rect 13168 11660 13508 11687
rect 4209 11649 13508 11660
rect 4209 11642 13204 11649
rect 4209 11622 11619 11642
rect 4209 11568 4245 11622
rect 4210 11566 4245 11568
rect 4301 11586 11619 11622
rect 11675 11593 13204 11642
rect 13260 11593 13416 11649
rect 13472 11593 13508 11649
rect 11675 11586 13508 11593
rect 4301 11568 13508 11586
rect 4301 11566 4336 11568
rect 4210 11404 4336 11566
rect 11582 11547 11712 11568
rect 13168 11554 13508 11568
rect 14290 11672 14416 11711
rect 14290 11616 14325 11672
rect 14381 11616 14416 11672
rect 4210 11348 4245 11404
rect 4301 11348 4336 11404
rect 4210 11309 4336 11348
rect 5328 11452 5668 11472
rect 10915 11452 11255 11472
rect 14290 11454 14416 11616
rect 14290 11452 14325 11454
rect 5328 11433 14325 11452
rect 5328 11377 5364 11433
rect 5420 11377 5576 11433
rect 5632 11377 10951 11433
rect 11007 11377 11163 11433
rect 11219 11398 14325 11433
rect 14381 11452 14416 11454
rect 15410 11463 15536 11502
rect 14381 11398 14417 11452
rect 11219 11377 14417 11398
rect 5328 11359 14417 11377
rect 15410 11407 15445 11463
rect 15501 11407 15536 11463
rect 5328 11338 5668 11359
rect 10915 11338 11255 11359
rect 6343 11243 6683 11264
rect 10232 11243 10572 11264
rect 15410 11245 15536 11407
rect 15410 11243 15445 11245
rect 6343 11225 15445 11243
rect 6343 11169 6379 11225
rect 6435 11169 6591 11225
rect 6647 11169 10268 11225
rect 10324 11169 10480 11225
rect 10536 11189 15445 11225
rect 15501 11243 15536 11245
rect 16530 11254 16656 11293
rect 15501 11189 15537 11243
rect 10536 11169 15537 11189
rect 6343 11150 15537 11169
rect 16530 11198 16565 11254
rect 16621 11198 16656 11254
rect 6343 11130 6683 11150
rect 10232 11130 10572 11150
rect 7463 11035 7803 11055
rect 9281 11035 9621 11055
rect 16530 11036 16656 11198
rect 16530 11035 16565 11036
rect 7463 11016 16565 11035
rect 7463 10960 7499 11016
rect 7555 10960 7711 11016
rect 7767 10960 9317 11016
rect 9373 10960 9529 11016
rect 9585 10980 16565 11016
rect 16621 11035 16656 11036
rect 17650 11046 17776 11085
rect 16621 10980 16657 11035
rect 9585 10960 16657 10980
rect 7463 10942 16657 10960
rect 17650 10990 17685 11046
rect 17741 10990 17776 11046
rect 7463 10921 7803 10942
rect 9281 10921 9621 10942
rect 16530 10941 16656 10942
rect 8390 10826 8730 10847
rect 17650 10828 17776 10990
rect 17650 10826 17685 10828
rect 8390 10808 17685 10826
rect 8390 10752 8426 10808
rect 8482 10752 8638 10808
rect 8694 10772 17685 10808
rect 17741 10826 17776 10828
rect 18770 10837 18896 10876
rect 17741 10772 17777 10826
rect 8694 10752 17777 10772
rect 8390 10733 17777 10752
rect 18770 10781 18805 10837
rect 18861 10781 18896 10837
rect 8390 10713 8730 10733
rect 7753 10617 8093 10638
rect 9808 10617 10148 10638
rect 18770 10619 18896 10781
rect 18770 10617 18805 10619
rect 7753 10599 18805 10617
rect 7753 10543 7789 10599
rect 7845 10543 8001 10599
rect 8057 10543 9844 10599
rect 9900 10543 10056 10599
rect 10112 10563 18805 10599
rect 18861 10617 18896 10619
rect 18861 10563 18897 10617
rect 10112 10543 18897 10563
rect 7753 10525 18897 10543
rect 7753 10504 8093 10525
rect 9808 10504 10148 10525
rect 18770 10524 18896 10525
rect 28591 10044 29353 10082
rect 28591 9988 28627 10044
rect 28683 9988 28838 10044
rect 28894 9988 29050 10044
rect 29106 9988 29261 10044
rect 29317 9988 29353 10044
rect 28591 9826 29353 9988
rect 1945 9366 14007 9792
rect 1945 9310 2402 9366
rect 2458 9310 2609 9366
rect 2665 9310 3129 9366
rect 3185 9310 4093 9366
rect 4149 9310 4300 9366
rect 4356 9310 4820 9366
rect 4876 9310 5784 9366
rect 5840 9310 5991 9366
rect 6047 9310 6511 9366
rect 6567 9326 14007 9366
rect 6567 9310 7669 9326
rect 1945 9270 7669 9310
rect 7725 9270 8117 9326
rect 8173 9270 8565 9326
rect 8621 9270 9302 9326
rect 9358 9270 9750 9326
rect 9806 9270 10198 9326
rect 10254 9270 10936 9326
rect 10992 9270 11384 9326
rect 11440 9270 11832 9326
rect 11888 9270 12570 9326
rect 12626 9270 13018 9326
rect 13074 9270 13466 9326
rect 13522 9270 14007 9326
rect 28591 9770 28627 9826
rect 28683 9770 28838 9826
rect 28894 9770 29050 9826
rect 29106 9770 29261 9826
rect 29317 9770 29353 9826
rect 28591 9608 29353 9770
rect 28591 9552 28627 9608
rect 28683 9552 28838 9608
rect 28894 9552 29050 9608
rect 29106 9552 29261 9608
rect 29317 9552 29353 9608
rect 28591 9390 29353 9552
rect 28591 9334 28627 9390
rect 28683 9334 28838 9390
rect 28894 9334 29050 9390
rect 29106 9334 29261 9390
rect 29317 9334 29353 9390
rect 28591 9296 29353 9334
rect 1945 9148 14007 9270
rect 1945 9092 2402 9148
rect 2458 9092 2609 9148
rect 2665 9092 3129 9148
rect 3185 9092 4093 9148
rect 4149 9092 4300 9148
rect 4356 9092 4820 9148
rect 4876 9092 5784 9148
rect 5840 9092 5991 9148
rect 6047 9092 6511 9148
rect 6567 9108 14007 9148
rect 6567 9092 7669 9108
rect 1945 9052 7669 9092
rect 7725 9052 8117 9108
rect 8173 9052 8565 9108
rect 8621 9052 9302 9108
rect 9358 9052 9750 9108
rect 9806 9052 10198 9108
rect 10254 9052 10936 9108
rect 10992 9052 11384 9108
rect 11440 9052 11832 9108
rect 11888 9052 12570 9108
rect 12626 9052 13018 9108
rect 13074 9052 13466 9108
rect 13522 9052 14007 9108
rect 1945 8930 14007 9052
rect 1945 8874 2402 8930
rect 2458 8874 2609 8930
rect 2665 8874 3129 8930
rect 3185 8874 4093 8930
rect 4149 8874 4300 8930
rect 4356 8874 4820 8930
rect 4876 8874 5784 8930
rect 5840 8874 5991 8930
rect 6047 8874 6511 8930
rect 6567 8890 14007 8930
rect 6567 8874 7669 8890
rect 1945 8834 7669 8874
rect 7725 8834 8117 8890
rect 8173 8834 8565 8890
rect 8621 8834 9302 8890
rect 9358 8834 9750 8890
rect 9806 8834 10198 8890
rect 10254 8834 10936 8890
rect 10992 8834 11384 8890
rect 11440 8834 11832 8890
rect 11888 8834 12570 8890
rect 12626 8834 13018 8890
rect 13074 8834 13466 8890
rect 13522 8834 14007 8890
rect 1945 8712 14007 8834
rect 1945 8656 2402 8712
rect 2458 8656 2609 8712
rect 2665 8656 3129 8712
rect 3185 8656 4093 8712
rect 4149 8656 4300 8712
rect 4356 8656 4820 8712
rect 4876 8656 5784 8712
rect 5840 8656 5991 8712
rect 6047 8656 6511 8712
rect 6567 8672 14007 8712
rect 6567 8656 7669 8672
rect 1945 8616 7669 8656
rect 7725 8616 8117 8672
rect 8173 8616 8565 8672
rect 8621 8616 9302 8672
rect 9358 8616 9750 8672
rect 9806 8616 10198 8672
rect 10254 8616 10936 8672
rect 10992 8616 11384 8672
rect 11440 8616 11832 8672
rect 11888 8616 12570 8672
rect 12626 8616 13018 8672
rect 13074 8616 13466 8672
rect 13522 8616 14007 8672
rect 1945 8532 14007 8616
rect 1945 7881 7228 8223
rect 1945 7825 2622 7881
rect 2678 7825 3136 7881
rect 3192 7825 4313 7881
rect 4369 7825 4827 7881
rect 4883 7825 6004 7881
rect 6060 7825 6518 7881
rect 6574 7863 7228 7881
rect 6574 7825 14239 7863
rect 1945 7821 14239 7825
rect 1945 7765 7669 7821
rect 7725 7765 8117 7821
rect 8173 7765 8565 7821
rect 8621 7765 9302 7821
rect 9358 7765 9750 7821
rect 9806 7765 10198 7821
rect 10254 7765 10936 7821
rect 10992 7765 11384 7821
rect 11440 7765 11832 7821
rect 11888 7765 12570 7821
rect 12626 7765 13018 7821
rect 13074 7765 13466 7821
rect 13522 7765 14239 7821
rect 1945 7664 14239 7765
rect 1945 7608 2622 7664
rect 2678 7608 3136 7664
rect 3192 7608 4313 7664
rect 4369 7608 4827 7664
rect 4883 7608 6004 7664
rect 6060 7608 6518 7664
rect 6574 7608 14239 7664
rect 1945 7603 14239 7608
rect 1945 7547 7669 7603
rect 7725 7547 8117 7603
rect 8173 7547 8565 7603
rect 8621 7547 9302 7603
rect 9358 7547 9750 7603
rect 9806 7547 10198 7603
rect 10254 7547 10936 7603
rect 10992 7547 11384 7603
rect 11440 7547 11832 7603
rect 11888 7547 12570 7603
rect 12626 7547 13018 7603
rect 13074 7547 13466 7603
rect 13522 7547 14239 7603
rect 1945 7446 14239 7547
rect 1945 7390 2622 7446
rect 2678 7390 3136 7446
rect 3192 7390 4313 7446
rect 4369 7390 4827 7446
rect 4883 7390 6004 7446
rect 6060 7390 6518 7446
rect 6574 7390 14239 7446
rect 1945 7385 14239 7390
rect 1945 7329 7669 7385
rect 7725 7329 8117 7385
rect 8173 7329 8565 7385
rect 8621 7329 9302 7385
rect 9358 7329 9750 7385
rect 9806 7329 10198 7385
rect 10254 7329 10936 7385
rect 10992 7329 11384 7385
rect 11440 7329 11832 7385
rect 11888 7329 12570 7385
rect 12626 7329 13018 7385
rect 13074 7329 13466 7385
rect 13522 7329 14239 7385
rect 1945 7228 14239 7329
rect 1945 7172 2622 7228
rect 2678 7172 3136 7228
rect 3192 7172 4313 7228
rect 4369 7172 4827 7228
rect 4883 7172 6004 7228
rect 6060 7172 6518 7228
rect 6574 7172 14239 7228
rect 1945 7010 14239 7172
rect 1945 6954 2622 7010
rect 2678 6954 3136 7010
rect 3192 6954 4313 7010
rect 4369 6954 4827 7010
rect 4883 6954 6004 7010
rect 6060 6954 6518 7010
rect 6574 6986 14239 7010
rect 6574 6954 13983 6986
rect 1945 6793 13983 6954
rect 1945 6737 2622 6793
rect 2678 6737 3136 6793
rect 3192 6737 4313 6793
rect 4369 6737 4827 6793
rect 4883 6737 6004 6793
rect 6060 6737 6518 6793
rect 6574 6737 13983 6793
rect 1945 6712 13983 6737
rect 1945 6711 8117 6712
rect 1945 6655 7673 6711
rect 7729 6656 8117 6711
rect 8173 6711 9750 6712
rect 8173 6656 8561 6711
rect 7729 6655 8561 6656
rect 8617 6655 9306 6711
rect 9362 6656 9750 6711
rect 9806 6711 11384 6712
rect 9806 6656 10194 6711
rect 9362 6655 10194 6656
rect 10250 6655 10940 6711
rect 10996 6656 11384 6711
rect 11440 6711 13018 6712
rect 11440 6656 11828 6711
rect 10996 6655 11828 6656
rect 11884 6655 12574 6711
rect 12630 6656 13018 6711
rect 13074 6711 13983 6712
rect 13074 6656 13462 6711
rect 12630 6655 13462 6656
rect 13518 6655 13983 6711
rect 1945 6494 13983 6655
rect 1945 6438 7673 6494
rect 7729 6438 8117 6494
rect 8173 6438 8561 6494
rect 8617 6438 9306 6494
rect 9362 6438 9750 6494
rect 9806 6438 10194 6494
rect 10250 6438 10940 6494
rect 10996 6438 11384 6494
rect 11440 6438 11828 6494
rect 11884 6438 12574 6494
rect 12630 6438 13018 6494
rect 13074 6438 13462 6494
rect 13518 6438 13983 6494
rect 1945 6277 13983 6438
rect 1945 6276 8117 6277
rect 1945 6220 7673 6276
rect 7729 6221 8117 6276
rect 8173 6276 9750 6277
rect 8173 6221 8561 6276
rect 7729 6220 8561 6221
rect 8617 6220 9306 6276
rect 9362 6221 9750 6276
rect 9806 6276 11384 6277
rect 9806 6221 10194 6276
rect 9362 6220 10194 6221
rect 10250 6220 10940 6276
rect 10996 6221 11384 6276
rect 11440 6276 13018 6277
rect 11440 6221 11828 6276
rect 10996 6220 11828 6221
rect 11884 6220 12574 6276
rect 12630 6221 13018 6276
rect 13074 6276 13983 6277
rect 13074 6221 13462 6276
rect 12630 6220 13462 6221
rect 13518 6220 13983 6276
rect 1945 6059 13983 6220
rect 1945 6058 8117 6059
rect 1945 6045 7673 6058
rect 7208 6002 7673 6045
rect 7729 6003 8117 6058
rect 8173 6058 9750 6059
rect 8173 6003 8561 6058
rect 7729 6002 8561 6003
rect 8617 6002 9306 6058
rect 9362 6003 9750 6058
rect 9806 6058 11384 6059
rect 9806 6003 10194 6058
rect 9362 6002 10194 6003
rect 10250 6002 10940 6058
rect 10996 6003 11384 6058
rect 11440 6058 13018 6059
rect 11440 6003 11828 6058
rect 10996 6002 11828 6003
rect 11884 6002 12574 6058
rect 12630 6003 13018 6058
rect 13074 6058 13983 6059
rect 13074 6003 13462 6058
rect 12630 6002 13462 6003
rect 13518 6002 13983 6058
rect 3580 5820 3706 5859
rect 3580 5764 3615 5820
rect 3671 5764 3706 5820
rect 3580 5750 3706 5764
rect 5271 5820 5397 5859
rect 5271 5764 5306 5820
rect 5362 5764 5397 5820
rect 5271 5750 5397 5764
rect 6962 5820 7088 5859
rect 6962 5764 6997 5820
rect 7053 5764 7088 5820
rect 6962 5750 7088 5764
rect 1951 5617 7088 5750
rect 3580 5602 3706 5617
rect 3580 5546 3615 5602
rect 3671 5546 3706 5602
rect 3580 5507 3706 5546
rect 5271 5602 5397 5617
rect 5271 5546 5306 5602
rect 5362 5546 5397 5602
rect 5271 5507 5397 5546
rect 6962 5602 7088 5617
rect 6962 5546 6997 5602
rect 7053 5546 7088 5602
rect 6962 5507 7088 5546
rect 7208 5841 13983 6002
rect 7208 5785 7673 5841
rect 7729 5785 8117 5841
rect 8173 5785 8561 5841
rect 8617 5785 9306 5841
rect 9362 5785 9750 5841
rect 9806 5785 10194 5841
rect 10250 5785 10940 5841
rect 10996 5785 11384 5841
rect 11440 5785 11828 5841
rect 11884 5785 12574 5841
rect 12630 5785 13018 5841
rect 13074 5785 13462 5841
rect 13518 5785 13983 5841
rect 7208 5624 13983 5785
rect 7208 5568 8117 5624
rect 8173 5568 9750 5624
rect 9806 5568 11384 5624
rect 11440 5568 13018 5624
rect 13074 5568 13983 5624
rect 7208 5406 13983 5568
rect 1960 5344 7087 5383
rect 1960 5288 3125 5344
rect 3181 5288 4816 5344
rect 4872 5288 6507 5344
rect 6563 5288 7087 5344
rect 1960 5249 7087 5288
rect 7208 5350 8117 5406
rect 8173 5350 9750 5406
rect 9806 5350 11384 5406
rect 11440 5350 13018 5406
rect 13074 5350 13983 5406
rect 7208 5261 13983 5350
rect 3090 5126 3216 5249
rect 3090 5070 3125 5126
rect 3181 5070 3216 5126
rect 3090 5031 3216 5070
rect 4781 5126 4907 5249
rect 4781 5070 4816 5126
rect 4872 5070 4907 5126
rect 4781 5031 4907 5070
rect 6472 5126 6598 5249
rect 6472 5070 6507 5126
rect 6563 5070 6598 5126
rect 6472 5031 6598 5070
rect 1980 3586 13864 3871
rect 1980 3189 8117 3586
rect 2004 2033 7032 2941
rect 7327 2594 8117 3189
rect 8173 2594 9751 3586
rect 9807 2594 11384 3586
rect 11440 2594 13018 3586
rect 13074 2594 13864 3586
rect 7327 2010 13864 2594
rect 7327 1954 9898 2010
rect 9954 1954 10109 2010
rect 10165 1954 10319 2010
rect 10375 1954 10530 2010
rect 10586 1954 10741 2010
rect 10797 1954 10952 2010
rect 11008 1954 11163 2010
rect 11219 1954 11373 2010
rect 11429 1954 11584 2010
rect 11640 1954 11796 2010
rect 11852 1954 12007 2010
rect 12063 1954 12217 2010
rect 12273 1954 12428 2010
rect 12484 1954 12639 2010
rect 12695 1954 12850 2010
rect 12906 1954 13061 2010
rect 13117 1954 13271 2010
rect 13327 1954 13482 2010
rect 13538 1954 13864 2010
rect 7327 1878 13864 1954
rect 7327 1862 7836 1878
rect 6338 1822 7836 1862
rect 7892 1822 13864 1878
rect 6338 1792 13864 1822
rect 6338 1736 9898 1792
rect 9954 1736 10109 1792
rect 10165 1736 10319 1792
rect 10375 1736 10530 1792
rect 10586 1736 10741 1792
rect 10797 1736 10952 1792
rect 11008 1736 11163 1792
rect 11219 1736 11373 1792
rect 11429 1736 11584 1792
rect 11640 1736 11796 1792
rect 11852 1736 12007 1792
rect 12063 1736 12217 1792
rect 12273 1736 12428 1792
rect 12484 1736 12639 1792
rect 12695 1736 12850 1792
rect 12906 1736 13061 1792
rect 13117 1736 13271 1792
rect 13327 1736 13482 1792
rect 13538 1736 13864 1792
rect 6338 1660 13864 1736
rect 6338 1604 7836 1660
rect 7892 1604 13864 1660
rect 6338 1466 13864 1604
rect 16097 1580 16589 1668
rect 7255 1180 13860 1250
rect 7255 1162 8472 1180
rect 7255 1106 7445 1162
rect 7501 1124 8472 1162
rect 8528 1175 13860 1180
rect 8528 1124 9658 1175
rect 7501 1119 9658 1124
rect 9714 1119 9869 1175
rect 9925 1119 10080 1175
rect 10136 1119 10291 1175
rect 10347 1119 10502 1175
rect 10558 1119 10712 1175
rect 10768 1119 10923 1175
rect 10979 1119 11134 1175
rect 11190 1119 11345 1175
rect 11401 1119 11556 1175
rect 11612 1119 11767 1175
rect 11823 1119 11978 1175
rect 12034 1119 12189 1175
rect 12245 1119 12400 1175
rect 12456 1119 12610 1175
rect 12666 1119 12821 1175
rect 12877 1119 13032 1175
rect 13088 1119 13243 1175
rect 13299 1119 13454 1175
rect 13510 1119 13860 1175
rect 7501 1106 13860 1119
rect 7255 962 13860 1106
rect 7255 944 8472 962
rect 7255 888 7445 944
rect 7501 906 8472 944
rect 8528 957 13860 962
rect 8528 906 9658 957
rect 7501 901 9658 906
rect 9714 901 9869 957
rect 9925 901 10080 957
rect 10136 901 10291 957
rect 10347 901 10502 957
rect 10558 901 10712 957
rect 10768 901 10923 957
rect 10979 901 11134 957
rect 11190 901 11345 957
rect 11401 901 11556 957
rect 11612 901 11767 957
rect 11823 901 11978 957
rect 12034 901 12189 957
rect 12245 901 12400 957
rect 12456 901 12610 957
rect 12666 901 12821 957
rect 12877 901 13032 957
rect 13088 901 13243 957
rect 13299 901 13454 957
rect 13510 901 13860 957
rect 7501 888 13860 901
rect 7255 786 13860 888
rect 21650 879 21934 889
rect 21650 615 21660 879
rect 21924 615 21934 879
rect 21650 605 21934 615
rect 21650 -189 21934 -179
rect 21650 -453 21660 -189
rect 21924 -453 21934 -189
rect 21650 -463 21934 -453
rect 300 -1332 640 -1293
rect 300 -1388 336 -1332
rect 392 -1388 548 -1332
rect 604 -1388 640 -1332
rect 300 -1426 640 -1388
rect 8028 -1332 8368 -1293
rect 8028 -1388 8064 -1332
rect 8120 -1388 8276 -1332
rect 8332 -1388 8368 -1332
rect 8028 -1426 8368 -1388
rect 29417 -1332 29757 -1293
rect 29417 -1388 29453 -1332
rect 29509 -1388 29665 -1332
rect 29721 -1388 29757 -1332
rect 29417 -1426 29757 -1388
use gen_512x8_128x8m81  gen_512x8_128x8m81_0
timestamp 1698431365
transform 1 0 14166 0 1 714
box -17790 -2370 17624 16428
use M1_NACTIVE4310590548746_128x8m81  M1_NACTIVE4310590548746_128x8m81_0
timestamp 1698431365
transform 0 -1 26031 1 0 27258
box 0 0 1 1
use M1_NACTIVE4310590548746_128x8m81  M1_NACTIVE4310590548746_128x8m81_1
timestamp 1698431365
transform 0 -1 25001 1 0 27314
box 0 0 1 1
use M1_PACTIVE4310590548747_128x8m81  M1_PACTIVE4310590548747_128x8m81_0
timestamp 1698431365
transform 1 0 3487 0 1 28973
box 0 0 1 1
use M1_PACTIVE4310590548747_128x8m81  M1_PACTIVE4310590548747_128x8m81_1
timestamp 1698431365
transform 1 0 10847 0 1 28973
box 0 0 1 1
use M1_PACTIVE4310590548748_128x8m81  M1_PACTIVE4310590548748_128x8m81_0
timestamp 1698431365
transform 1 0 23865 0 1 28384
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1698431365
transform -1 0 29587 0 1 28861
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1698431365
transform -1 0 29587 0 1 982
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1698431365
transform 1 0 470 0 1 28861
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_3
timestamp 1698431365
transform 1 0 470 0 1 982
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_0
timestamp 1698431365
transform 1 0 865 0 1 102
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_1
timestamp 1698431365
transform 1 0 29191 0 1 102
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_2
timestamp 1698431365
transform 1 0 9050 0 1 154
box 0 0 1 1
use M2_M1$$201262124_128x8m81  M2_M1$$201262124_128x8m81_0
timestamp 1698431365
transform 1 0 9050 0 1 263
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_0
timestamp 1698431365
transform 1 0 28796 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_1
timestamp 1698431365
transform 1 0 28555 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_2
timestamp 1698431365
transform 1 0 28313 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_3
timestamp 1698431365
transform 1 0 28071 0 1 886
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_0
timestamp 1698431365
transform 1 0 1779 0 1 982
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_1
timestamp 1698431365
transform 1 0 1537 0 1 982
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_2
timestamp 1698431365
transform 1 0 1296 0 1 982
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_0
timestamp 1698431365
transform -1 0 29587 0 1 28861
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_1
timestamp 1698431365
transform 1 0 470 0 1 28861
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_0
timestamp 1698431365
transform -1 0 29587 0 1 -1360
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_1
timestamp 1698431365
transform 1 0 470 0 1 -1360
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_2
timestamp 1698431365
transform 1 0 8198 0 1 -1360
box 0 0 1 1
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_0
timestamp 1698431365
transform 1 0 28972 0 1 29671
box 0 0 1 1
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_1
timestamp 1698431365
transform 1 0 1085 0 1 29671
box 0 0 1 1
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_2
timestamp 1698431365
transform 1 0 28972 0 1 9689
box 0 0 1 1
use M3_M24310590548749_128x8m81  M3_M24310590548749_128x8m81_0
timestamp 1698431365
transform 1 0 21792 0 1 -321
box 0 0 1 1
use M3_M24310590548749_128x8m81  M3_M24310590548749_128x8m81_1
timestamp 1698431365
transform 1 0 21792 0 1 747
box 0 0 1 1
use prexdec_top_128x8m81  prexdec_top_128x8m81_0
timestamp 1698431365
transform 1 0 1357 0 1 17581
box 325 -1 27066 12091
use ypredec1_128x8m81  ypredec1_128x8m81_0
timestamp 1698431365
transform 1 0 1561 0 1 560
box 364 179 18378 16305
<< labels >>
flabel metal3 s 8281 -1000 8281 -1000 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 8281 -352 8281 -352 0 FreeSans 448 0 0 0 VDD
port 2 nsew
rlabel metal3 s 28175 14906 28175 14906 4 RYS[7]
port 3 nsew
rlabel metal3 s 28175 14565 28175 14565 4 RYS[6]
port 4 nsew
rlabel metal3 s 28175 14225 28175 14225 4 RYS[5]
port 5 nsew
rlabel metal3 s 28175 13885 28175 13885 4 RYS[4]
port 6 nsew
rlabel metal3 s 28175 13545 28175 13545 4 RYS[3]
port 7 nsew
rlabel metal3 s 28175 13205 28175 13205 4 RYS[2]
port 8 nsew
rlabel metal3 s 28175 12865 28175 12865 4 RYS[1]
port 9 nsew
rlabel metal3 s 28175 12525 28175 12525 4 RYS[0]
port 10 nsew
rlabel metal3 s 1805 12525 1805 12525 4 LYS[0]
port 11 nsew
rlabel metal3 s 1805 12865 1805 12865 4 LYS[1]
port 12 nsew
rlabel metal3 s 1805 13205 1805 13205 4 LYS[2]
port 13 nsew
rlabel metal3 s 1805 13545 1805 13545 4 LYS[3]
port 14 nsew
rlabel metal3 s 1805 14565 1805 14565 4 LYS[6]
port 15 nsew
rlabel metal3 s 1805 14225 1805 14225 4 LYS[5]
port 16 nsew
rlabel metal3 s 1805 13885 1805 13885 4 LYS[4]
port 17 nsew
rlabel metal3 s 26861 29671 26861 29671 4 men
port 18 nsew
rlabel metal3 s 1805 14906 1805 14906 4 LYS[7]
port 19 nsew
rlabel metal3 s 27957 5019 27957 5019 4 tblhl
port 20 nsew
flabel metal3 s 6236 9021 6236 9021 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 18161 6236 18161 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 3499 6236 3499 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 1395 6236 1395 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 8281 1059 8281 1059 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 18981 6236 18981 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 24007 6236 24007 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 2448 6236 2448 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 28103 6236 28103 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 26066 6236 26066 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 6539 6236 6539 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 15970 6236 15970 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 27112 6236 27112 0 FreeSans 448 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 20288 6236 20288 0 FreeSans 448 0 0 0 VSS
port 1 nsew
flabel metal2 s 16356 -1340 16356 -1340 0 FreeSans 1000 0 0 0 IGWEN
port 21 nsew
rlabel metal2 s 9726 28748 9726 28748 4 xb[3]
port 22 nsew
rlabel metal2 s 10163 28755 10163 28755 4 xb[2]
port 23 nsew
rlabel metal2 s 11966 28730 11966 28730 4 xb[0]
port 24 nsew
rlabel metal2 s 17221 28931 17221 28931 4 xa[7]
port 25 nsew
rlabel metal2 s 17572 28931 17572 28931 4 xa[6]
port 26 nsew
rlabel metal2 s 18855 28931 18855 28931 4 xa[5]
port 27 nsew
rlabel metal2 s 19211 28931 19211 28931 4 xa[4]
port 28 nsew
rlabel metal2 s 20491 28931 20491 28931 4 xa[3]
port 29 nsew
rlabel metal2 s 20833 28931 20833 28931 4 xa[2]
port 30 nsew
rlabel metal2 s 6821 -1360 6821 -1360 4 A[0]
port 31 nsew
rlabel metal2 s 22924 -1360 22924 -1360 4 CEN
port 32 nsew
rlabel metal2 s 11527 28712 11527 28712 4 xb[1]
port 33 nsew
rlabel metal2 s 10135 28705 10135 28705 4 xb[2]
port 23 nsew
rlabel metal2 s 11931 28700 11931 28700 4 xb[0]
port 24 nsew
rlabel metal2 s 2400 28705 2400 28705 4 xc[3]
port 34 nsew
rlabel metal2 s 4190 28700 4190 28700 4 xc[1]
port 35 nsew
rlabel metal2 s 2756 28705 2756 28705 4 xc[2]
port 36 nsew
rlabel metal2 s 4552 28700 4552 28700 4 xc[0]
port 37 nsew
rlabel metal2 s 22480 28931 22480 28931 4 xa[0]
port 38 nsew
rlabel metal2 s 22120 28931 22120 28931 4 xa[1]
port 39 nsew
rlabel metal2 s 1296 -1360 1296 -1360 4 A[9]
port 40 nsew
rlabel metal2 s 1779 -1360 1779 -1360 4 A[7]
port 41 nsew
rlabel metal2 s 470 -1360 470 -1360 4 CLK
port 42 nsew
rlabel metal2 s 11569 28700 11569 28700 4 xb[1]
port 33 nsew
rlabel metal2 s 9779 28705 9779 28705 4 xb[3]
port 22 nsew
rlabel metal2 s 3437 -1360 3437 -1360 4 A[2]
port 43 nsew
rlabel metal2 s 5128 -1360 5128 -1360 4 A[1]
port 44 nsew
rlabel metal2 s 28071 -1360 28071 -1360 4 A[6]
port 45 nsew
rlabel metal2 s 28796 -1360 28796 -1360 4 A[3]
port 46 nsew
rlabel metal2 s 28555 -1360 28555 -1360 4 A[4]
port 47 nsew
rlabel metal2 s 28313 -1360 28313 -1360 4 A[5]
port 48 nsew
rlabel metal2 s 1537 -1360 1537 -1360 4 A[8]
port 49 nsew
flabel metal1 s 22454 1053 22454 1053 0 FreeSans 1000 0 0 0 GWE
port 50 nsew
<< properties >>
string GDS_END 2297908
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2287334
string path 80.485 8.120 82.945 8.120 
<< end >>
