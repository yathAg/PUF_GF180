magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< pwell >>
rect 5431 6633 7607 11633
rect 7867 6633 10043 11633
rect 5431 621 7607 5621
rect 7867 621 10043 5621
<< mvndiff >>
rect 5431 11596 5519 11633
rect 5431 6670 5444 11596
rect 5490 6670 5519 11596
rect 5431 6633 5519 6670
rect 7519 11596 7607 11633
rect 7519 6670 7548 11596
rect 7594 6670 7607 11596
rect 7519 6633 7607 6670
rect 7867 11596 7955 11633
rect 7867 6670 7880 11596
rect 7926 6670 7955 11596
rect 7867 6633 7955 6670
rect 9955 11596 10043 11633
rect 9955 6670 9984 11596
rect 10030 6670 10043 11596
rect 9955 6633 10043 6670
rect 5431 5584 5519 5621
rect 5431 658 5444 5584
rect 5490 658 5519 5584
rect 5431 621 5519 658
rect 7519 5584 7607 5621
rect 7519 658 7548 5584
rect 7594 658 7607 5584
rect 7519 621 7607 658
rect 7867 5584 7955 5621
rect 7867 658 7880 5584
rect 7926 658 7955 5584
rect 7867 621 7955 658
rect 9955 5584 10043 5621
rect 9955 658 9984 5584
rect 10030 658 10043 5584
rect 9955 621 10043 658
<< mvndiffc >>
rect 5444 6670 5490 11596
rect 7548 6670 7594 11596
rect 7880 6670 7926 11596
rect 9984 6670 10030 11596
rect 5444 658 5490 5584
rect 7548 658 7594 5584
rect 7880 658 7926 5584
rect 9984 658 10030 5584
<< psubdiff >>
rect 4904 12298 10576 12320
rect 4904 12252 4926 12298
rect 4972 12252 5040 12298
rect 5086 12252 5217 12298
rect 5263 12252 5331 12298
rect 5377 12252 5445 12298
rect 5491 12252 5559 12298
rect 5605 12252 5673 12298
rect 5719 12252 5787 12298
rect 5833 12252 5901 12298
rect 5947 12252 6015 12298
rect 6061 12252 6129 12298
rect 6175 12252 6243 12298
rect 6289 12252 6357 12298
rect 6403 12252 6471 12298
rect 6517 12252 6585 12298
rect 6631 12252 6699 12298
rect 6745 12252 6813 12298
rect 6859 12252 6927 12298
rect 6973 12252 7041 12298
rect 7087 12252 7155 12298
rect 7201 12252 7269 12298
rect 7315 12252 7383 12298
rect 7429 12252 7497 12298
rect 7543 12252 7611 12298
rect 7657 12252 7725 12298
rect 7771 12252 7839 12298
rect 7885 12252 7953 12298
rect 7999 12252 8067 12298
rect 8113 12252 8181 12298
rect 8227 12252 8295 12298
rect 8341 12252 8409 12298
rect 8455 12252 8523 12298
rect 8569 12252 8637 12298
rect 8683 12252 8751 12298
rect 8797 12252 8865 12298
rect 8911 12252 8979 12298
rect 9025 12252 9093 12298
rect 9139 12252 9207 12298
rect 9253 12252 9321 12298
rect 9367 12252 9435 12298
rect 9481 12252 9549 12298
rect 9595 12252 9663 12298
rect 9709 12252 9777 12298
rect 9823 12252 9891 12298
rect 9937 12252 10005 12298
rect 10051 12252 10119 12298
rect 10165 12252 10233 12298
rect 10279 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10576 12298
rect 4904 12184 10576 12252
rect 4904 12138 4926 12184
rect 4972 12138 5040 12184
rect 5086 12138 5217 12184
rect 5263 12138 5331 12184
rect 5377 12138 5445 12184
rect 5491 12138 5559 12184
rect 5605 12138 5673 12184
rect 5719 12138 5787 12184
rect 5833 12138 5901 12184
rect 5947 12138 6015 12184
rect 6061 12138 6129 12184
rect 6175 12138 6243 12184
rect 6289 12138 6357 12184
rect 6403 12138 6471 12184
rect 6517 12138 6585 12184
rect 6631 12138 6699 12184
rect 6745 12138 6813 12184
rect 6859 12138 6927 12184
rect 6973 12138 7041 12184
rect 7087 12138 7155 12184
rect 7201 12138 7269 12184
rect 7315 12138 7383 12184
rect 7429 12138 7497 12184
rect 7543 12138 7611 12184
rect 7657 12138 7725 12184
rect 7771 12138 7839 12184
rect 7885 12138 7953 12184
rect 7999 12138 8067 12184
rect 8113 12138 8181 12184
rect 8227 12138 8295 12184
rect 8341 12138 8409 12184
rect 8455 12138 8523 12184
rect 8569 12138 8637 12184
rect 8683 12138 8751 12184
rect 8797 12138 8865 12184
rect 8911 12138 8979 12184
rect 9025 12138 9093 12184
rect 9139 12138 9207 12184
rect 9253 12138 9321 12184
rect 9367 12138 9435 12184
rect 9481 12138 9549 12184
rect 9595 12138 9663 12184
rect 9709 12138 9777 12184
rect 9823 12138 9891 12184
rect 9937 12138 10005 12184
rect 10051 12138 10119 12184
rect 10165 12138 10233 12184
rect 10279 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10576 12184
rect 4904 12116 10576 12138
rect 4904 12070 5108 12116
rect 4904 12024 4926 12070
rect 4972 12024 5040 12070
rect 5086 12024 5108 12070
rect 4904 11500 5108 12024
rect 10372 12070 10576 12116
rect 10372 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10576 12070
rect 10372 11956 10576 12024
rect 10372 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10576 11956
rect 10372 11842 10576 11910
rect 10372 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10576 11842
rect 10372 11728 10576 11796
rect 10372 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10576 11728
rect 4904 11454 4926 11500
rect 4972 11454 5040 11500
rect 5086 11454 5108 11500
rect 4904 11386 5108 11454
rect 4904 11340 4926 11386
rect 4972 11340 5040 11386
rect 5086 11340 5108 11386
rect 4904 11272 5108 11340
rect 4904 11226 4926 11272
rect 4972 11226 5040 11272
rect 5086 11226 5108 11272
rect 4904 11158 5108 11226
rect 4904 11112 4926 11158
rect 4972 11112 5040 11158
rect 5086 11112 5108 11158
rect 4904 11044 5108 11112
rect 4904 10998 4926 11044
rect 4972 10998 5040 11044
rect 5086 10998 5108 11044
rect 4904 10930 5108 10998
rect 4904 10884 4926 10930
rect 4972 10884 5040 10930
rect 5086 10884 5108 10930
rect 4904 10816 5108 10884
rect 4904 10770 4926 10816
rect 4972 10770 5040 10816
rect 5086 10770 5108 10816
rect 4904 10702 5108 10770
rect 4904 10656 4926 10702
rect 4972 10656 5040 10702
rect 5086 10656 5108 10702
rect 4904 10588 5108 10656
rect 4904 10542 4926 10588
rect 4972 10542 5040 10588
rect 5086 10542 5108 10588
rect 4904 10474 5108 10542
rect 4904 10428 4926 10474
rect 4972 10428 5040 10474
rect 5086 10428 5108 10474
rect 4904 10360 5108 10428
rect 4904 10314 4926 10360
rect 4972 10314 5040 10360
rect 5086 10314 5108 10360
rect 4904 10246 5108 10314
rect 4904 10200 4926 10246
rect 4972 10200 5040 10246
rect 5086 10200 5108 10246
rect 4904 10132 5108 10200
rect 4904 10086 4926 10132
rect 4972 10086 5040 10132
rect 5086 10086 5108 10132
rect 4904 10018 5108 10086
rect 4904 9972 4926 10018
rect 4972 9972 5040 10018
rect 5086 9972 5108 10018
rect 4904 9904 5108 9972
rect 4904 9858 4926 9904
rect 4972 9858 5040 9904
rect 5086 9858 5108 9904
rect 4904 9790 5108 9858
rect 4904 9744 4926 9790
rect 4972 9744 5040 9790
rect 5086 9744 5108 9790
rect 4904 9676 5108 9744
rect 4904 9630 4926 9676
rect 4972 9630 5040 9676
rect 5086 9630 5108 9676
rect 4904 9562 5108 9630
rect 4904 9516 4926 9562
rect 4972 9516 5040 9562
rect 5086 9516 5108 9562
rect 4904 9448 5108 9516
rect 4904 9402 4926 9448
rect 4972 9402 5040 9448
rect 5086 9402 5108 9448
rect 4904 9334 5108 9402
rect 4904 9288 4926 9334
rect 4972 9288 5040 9334
rect 5086 9288 5108 9334
rect 4904 9220 5108 9288
rect 4904 9174 4926 9220
rect 4972 9174 5040 9220
rect 5086 9174 5108 9220
rect 4904 9106 5108 9174
rect 4904 9060 4926 9106
rect 4972 9060 5040 9106
rect 5086 9060 5108 9106
rect 4904 8992 5108 9060
rect 4904 8946 4926 8992
rect 4972 8946 5040 8992
rect 5086 8946 5108 8992
rect 4904 8878 5108 8946
rect 4904 8832 4926 8878
rect 4972 8832 5040 8878
rect 5086 8832 5108 8878
rect 4904 8764 5108 8832
rect 4904 8718 4926 8764
rect 4972 8718 5040 8764
rect 5086 8718 5108 8764
rect 4904 8650 5108 8718
rect 4904 8604 4926 8650
rect 4972 8604 5040 8650
rect 5086 8604 5108 8650
rect 4904 8536 5108 8604
rect 4904 8490 4926 8536
rect 4972 8490 5040 8536
rect 5086 8490 5108 8536
rect 4904 8422 5108 8490
rect 4904 8376 4926 8422
rect 4972 8376 5040 8422
rect 5086 8376 5108 8422
rect 4904 8308 5108 8376
rect 4904 8262 4926 8308
rect 4972 8262 5040 8308
rect 5086 8262 5108 8308
rect 4904 8194 5108 8262
rect 4904 8148 4926 8194
rect 4972 8148 5040 8194
rect 5086 8148 5108 8194
rect 4904 8080 5108 8148
rect 4904 8034 4926 8080
rect 4972 8034 5040 8080
rect 5086 8034 5108 8080
rect 4904 7966 5108 8034
rect 4904 7920 4926 7966
rect 4972 7920 5040 7966
rect 5086 7920 5108 7966
rect 4904 7852 5108 7920
rect 4904 7806 4926 7852
rect 4972 7806 5040 7852
rect 5086 7806 5108 7852
rect 4904 7738 5108 7806
rect 4904 7692 4926 7738
rect 4972 7692 5040 7738
rect 5086 7692 5108 7738
rect 4904 7624 5108 7692
rect 4904 7578 4926 7624
rect 4972 7578 5040 7624
rect 5086 7578 5108 7624
rect 4904 7510 5108 7578
rect 4904 7464 4926 7510
rect 4972 7464 5040 7510
rect 5086 7464 5108 7510
rect 4904 7396 5108 7464
rect 4904 7350 4926 7396
rect 4972 7350 5040 7396
rect 5086 7350 5108 7396
rect 4904 7282 5108 7350
rect 4904 7236 4926 7282
rect 4972 7236 5040 7282
rect 5086 7236 5108 7282
rect 4904 7168 5108 7236
rect 4904 7122 4926 7168
rect 4972 7122 5040 7168
rect 5086 7122 5108 7168
rect 4904 7054 5108 7122
rect 4904 7008 4926 7054
rect 4972 7008 5040 7054
rect 5086 7008 5108 7054
rect 4904 6940 5108 7008
rect 4904 6894 4926 6940
rect 4972 6894 5040 6940
rect 5086 6894 5108 6940
rect 4904 6826 5108 6894
rect 4904 6780 4926 6826
rect 4972 6780 5040 6826
rect 5086 6780 5108 6826
rect 4904 6712 5108 6780
rect 4904 6666 4926 6712
rect 4972 6666 5040 6712
rect 5086 6666 5108 6712
rect 4904 6598 5108 6666
rect 10372 11614 10576 11682
rect 10372 11568 10394 11614
rect 10440 11568 10508 11614
rect 10554 11568 10576 11614
rect 10372 11500 10576 11568
rect 10372 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10576 11500
rect 10372 11386 10576 11454
rect 10372 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10576 11386
rect 10372 11272 10576 11340
rect 10372 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10576 11272
rect 10372 11158 10576 11226
rect 10372 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10576 11158
rect 10372 11044 10576 11112
rect 10372 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10576 11044
rect 10372 10930 10576 10998
rect 10372 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10576 10930
rect 10372 10816 10576 10884
rect 10372 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10576 10816
rect 10372 10702 10576 10770
rect 10372 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10576 10702
rect 10372 10588 10576 10656
rect 10372 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10576 10588
rect 10372 10474 10576 10542
rect 10372 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10576 10474
rect 10372 10360 10576 10428
rect 10372 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10576 10360
rect 10372 10246 10576 10314
rect 10372 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10576 10246
rect 10372 10132 10576 10200
rect 10372 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10576 10132
rect 10372 10018 10576 10086
rect 10372 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10576 10018
rect 10372 9904 10576 9972
rect 10372 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10576 9904
rect 10372 9790 10576 9858
rect 10372 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10576 9790
rect 10372 9676 10576 9744
rect 10372 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10576 9676
rect 10372 9562 10576 9630
rect 10372 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10576 9562
rect 10372 9448 10576 9516
rect 10372 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10576 9448
rect 10372 9334 10576 9402
rect 10372 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10576 9334
rect 10372 9220 10576 9288
rect 10372 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10576 9220
rect 10372 9106 10576 9174
rect 10372 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10576 9106
rect 10372 8992 10576 9060
rect 10372 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10576 8992
rect 10372 8878 10576 8946
rect 10372 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10576 8878
rect 10372 8764 10576 8832
rect 10372 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10576 8764
rect 10372 8650 10576 8718
rect 10372 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10576 8650
rect 10372 8536 10576 8604
rect 10372 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10576 8536
rect 10372 8422 10576 8490
rect 10372 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10576 8422
rect 10372 8308 10576 8376
rect 10372 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10576 8308
rect 10372 8194 10576 8262
rect 10372 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10576 8194
rect 10372 8080 10576 8148
rect 10372 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10576 8080
rect 10372 7966 10576 8034
rect 10372 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10576 7966
rect 10372 7852 10576 7920
rect 10372 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10576 7852
rect 10372 7738 10576 7806
rect 10372 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10576 7738
rect 10372 7624 10576 7692
rect 10372 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10576 7624
rect 10372 7510 10576 7578
rect 10372 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10576 7510
rect 10372 7396 10576 7464
rect 10372 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10576 7396
rect 10372 7282 10576 7350
rect 10372 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10576 7282
rect 10372 7168 10576 7236
rect 10372 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10576 7168
rect 10372 7054 10576 7122
rect 10372 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10576 7054
rect 10372 6940 10576 7008
rect 10372 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10576 6940
rect 10372 6826 10576 6894
rect 10372 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10576 6826
rect 10372 6712 10576 6780
rect 10372 6666 10394 6712
rect 10440 6666 10508 6712
rect 10554 6666 10576 6712
rect 4904 6552 4926 6598
rect 4972 6552 5040 6598
rect 5086 6552 5108 6598
rect 4904 6484 5108 6552
rect 10372 6598 10576 6666
rect 10372 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10576 6598
rect 4904 6438 4926 6484
rect 4972 6438 5040 6484
rect 5086 6438 5108 6484
rect 4904 6370 5108 6438
rect 4904 6324 4926 6370
rect 4972 6324 5040 6370
rect 5086 6324 5108 6370
rect 4904 6256 5108 6324
rect 4904 6210 4926 6256
rect 4972 6210 5040 6256
rect 5086 6229 5108 6256
rect 10372 6484 10576 6552
rect 10372 6438 10394 6484
rect 10440 6438 10508 6484
rect 10554 6438 10576 6484
rect 10372 6370 10576 6438
rect 10372 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10576 6370
rect 10372 6256 10576 6324
rect 10372 6229 10394 6256
rect 5086 6210 10394 6229
rect 10440 6210 10508 6256
rect 10554 6210 10576 6256
rect 4904 6207 10576 6210
rect 4904 6161 5214 6207
rect 5260 6161 5328 6207
rect 5374 6161 5442 6207
rect 5488 6161 5556 6207
rect 5602 6161 5670 6207
rect 5716 6161 5784 6207
rect 5830 6161 5898 6207
rect 5944 6161 6012 6207
rect 6058 6161 6126 6207
rect 6172 6161 6240 6207
rect 6286 6161 6354 6207
rect 6400 6161 6468 6207
rect 6514 6161 6582 6207
rect 6628 6161 6696 6207
rect 6742 6161 6810 6207
rect 6856 6161 6924 6207
rect 6970 6161 7038 6207
rect 7084 6161 7152 6207
rect 7198 6161 7266 6207
rect 7312 6161 7380 6207
rect 7426 6161 7494 6207
rect 7540 6161 7608 6207
rect 7654 6161 7722 6207
rect 7768 6161 7836 6207
rect 7882 6161 7950 6207
rect 7996 6161 8064 6207
rect 8110 6161 8178 6207
rect 8224 6161 8292 6207
rect 8338 6161 8406 6207
rect 8452 6161 8520 6207
rect 8566 6161 8634 6207
rect 8680 6161 8748 6207
rect 8794 6161 8862 6207
rect 8908 6161 8976 6207
rect 9022 6161 9090 6207
rect 9136 6161 9204 6207
rect 9250 6161 9318 6207
rect 9364 6161 9432 6207
rect 9478 6161 9546 6207
rect 9592 6161 9660 6207
rect 9706 6161 9774 6207
rect 9820 6161 9888 6207
rect 9934 6161 10002 6207
rect 10048 6161 10116 6207
rect 10162 6161 10230 6207
rect 10276 6161 10576 6207
rect 4904 6142 10576 6161
rect 4904 6096 4926 6142
rect 4972 6096 5040 6142
rect 5086 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10576 6142
rect 4904 6093 10576 6096
rect 4904 6047 5214 6093
rect 5260 6047 5328 6093
rect 5374 6047 5442 6093
rect 5488 6047 5556 6093
rect 5602 6047 5670 6093
rect 5716 6047 5784 6093
rect 5830 6047 5898 6093
rect 5944 6047 6012 6093
rect 6058 6047 6126 6093
rect 6172 6047 6240 6093
rect 6286 6047 6354 6093
rect 6400 6047 6468 6093
rect 6514 6047 6582 6093
rect 6628 6047 6696 6093
rect 6742 6047 6810 6093
rect 6856 6047 6924 6093
rect 6970 6047 7038 6093
rect 7084 6047 7152 6093
rect 7198 6047 7266 6093
rect 7312 6047 7380 6093
rect 7426 6047 7494 6093
rect 7540 6047 7608 6093
rect 7654 6047 7722 6093
rect 7768 6047 7836 6093
rect 7882 6047 7950 6093
rect 7996 6047 8064 6093
rect 8110 6047 8178 6093
rect 8224 6047 8292 6093
rect 8338 6047 8406 6093
rect 8452 6047 8520 6093
rect 8566 6047 8634 6093
rect 8680 6047 8748 6093
rect 8794 6047 8862 6093
rect 8908 6047 8976 6093
rect 9022 6047 9090 6093
rect 9136 6047 9204 6093
rect 9250 6047 9318 6093
rect 9364 6047 9432 6093
rect 9478 6047 9546 6093
rect 9592 6047 9660 6093
rect 9706 6047 9774 6093
rect 9820 6047 9888 6093
rect 9934 6047 10002 6093
rect 10048 6047 10116 6093
rect 10162 6047 10230 6093
rect 10276 6047 10576 6093
rect 4904 6028 10576 6047
rect 4904 5982 4926 6028
rect 4972 5982 5040 6028
rect 5086 6025 10394 6028
rect 5086 5982 5108 6025
rect 4904 5914 5108 5982
rect 4904 5868 4926 5914
rect 4972 5868 5040 5914
rect 5086 5868 5108 5914
rect 4904 5800 5108 5868
rect 4904 5754 4926 5800
rect 4972 5754 5040 5800
rect 5086 5754 5108 5800
rect 4904 5686 5108 5754
rect 10372 5982 10394 6025
rect 10440 5982 10508 6028
rect 10554 5982 10576 6028
rect 10372 5914 10576 5982
rect 10372 5868 10394 5914
rect 10440 5868 10508 5914
rect 10554 5868 10576 5914
rect 10372 5800 10576 5868
rect 10372 5754 10394 5800
rect 10440 5754 10508 5800
rect 10554 5754 10576 5800
rect 4904 5640 4926 5686
rect 4972 5640 5040 5686
rect 5086 5640 5108 5686
rect 4904 5572 5108 5640
rect 10372 5686 10576 5754
rect 10372 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10576 5686
rect 4904 5526 4926 5572
rect 4972 5526 5040 5572
rect 5086 5526 5108 5572
rect 4904 5458 5108 5526
rect 4904 5412 4926 5458
rect 4972 5412 5040 5458
rect 5086 5412 5108 5458
rect 4904 5344 5108 5412
rect 4904 5298 4926 5344
rect 4972 5298 5040 5344
rect 5086 5298 5108 5344
rect 4904 5230 5108 5298
rect 4904 5184 4926 5230
rect 4972 5184 5040 5230
rect 5086 5184 5108 5230
rect 4904 5116 5108 5184
rect 4904 5070 4926 5116
rect 4972 5070 5040 5116
rect 5086 5070 5108 5116
rect 4904 5002 5108 5070
rect 4904 4956 4926 5002
rect 4972 4956 5040 5002
rect 5086 4956 5108 5002
rect 4904 4888 5108 4956
rect 4904 4842 4926 4888
rect 4972 4842 5040 4888
rect 5086 4842 5108 4888
rect 4904 4774 5108 4842
rect 4904 4728 4926 4774
rect 4972 4728 5040 4774
rect 5086 4728 5108 4774
rect 4904 4660 5108 4728
rect 4904 4614 4926 4660
rect 4972 4614 5040 4660
rect 5086 4614 5108 4660
rect 4904 4546 5108 4614
rect 4904 4500 4926 4546
rect 4972 4500 5040 4546
rect 5086 4500 5108 4546
rect 4904 4432 5108 4500
rect 4904 4386 4926 4432
rect 4972 4386 5040 4432
rect 5086 4386 5108 4432
rect 4904 4318 5108 4386
rect 4904 4272 4926 4318
rect 4972 4272 5040 4318
rect 5086 4272 5108 4318
rect 4904 4204 5108 4272
rect 4904 4158 4926 4204
rect 4972 4158 5040 4204
rect 5086 4158 5108 4204
rect 4904 4090 5108 4158
rect 4904 4044 4926 4090
rect 4972 4044 5040 4090
rect 5086 4044 5108 4090
rect 4904 3976 5108 4044
rect 4904 3930 4926 3976
rect 4972 3930 5040 3976
rect 5086 3930 5108 3976
rect 4904 3862 5108 3930
rect 4904 3816 4926 3862
rect 4972 3816 5040 3862
rect 5086 3816 5108 3862
rect 4904 3748 5108 3816
rect 4904 3702 4926 3748
rect 4972 3702 5040 3748
rect 5086 3702 5108 3748
rect 4904 3634 5108 3702
rect 4904 3588 4926 3634
rect 4972 3588 5040 3634
rect 5086 3588 5108 3634
rect 4904 3520 5108 3588
rect 4904 3474 4926 3520
rect 4972 3474 5040 3520
rect 5086 3474 5108 3520
rect 4904 3406 5108 3474
rect 4904 3360 4926 3406
rect 4972 3360 5040 3406
rect 5086 3360 5108 3406
rect 4904 3292 5108 3360
rect 4904 3246 4926 3292
rect 4972 3246 5040 3292
rect 5086 3246 5108 3292
rect 4904 3178 5108 3246
rect 4904 3132 4926 3178
rect 4972 3132 5040 3178
rect 5086 3132 5108 3178
rect 4904 3064 5108 3132
rect 4904 3018 4926 3064
rect 4972 3018 5040 3064
rect 5086 3018 5108 3064
rect 4904 2950 5108 3018
rect 4904 2904 4926 2950
rect 4972 2904 5040 2950
rect 5086 2904 5108 2950
rect 4904 2836 5108 2904
rect 4904 2790 4926 2836
rect 4972 2790 5040 2836
rect 5086 2790 5108 2836
rect 4904 2722 5108 2790
rect 4904 2676 4926 2722
rect 4972 2676 5040 2722
rect 5086 2676 5108 2722
rect 4904 2608 5108 2676
rect 4904 2562 4926 2608
rect 4972 2562 5040 2608
rect 5086 2562 5108 2608
rect 4904 2494 5108 2562
rect 4904 2448 4926 2494
rect 4972 2448 5040 2494
rect 5086 2448 5108 2494
rect 4904 2380 5108 2448
rect 4904 2334 4926 2380
rect 4972 2334 5040 2380
rect 5086 2334 5108 2380
rect 4904 2266 5108 2334
rect 4904 2220 4926 2266
rect 4972 2220 5040 2266
rect 5086 2220 5108 2266
rect 4904 2152 5108 2220
rect 4904 2106 4926 2152
rect 4972 2106 5040 2152
rect 5086 2106 5108 2152
rect 4904 2038 5108 2106
rect 4904 1992 4926 2038
rect 4972 1992 5040 2038
rect 5086 1992 5108 2038
rect 4904 1924 5108 1992
rect 4904 1878 4926 1924
rect 4972 1878 5040 1924
rect 5086 1878 5108 1924
rect 4904 1810 5108 1878
rect 4904 1764 4926 1810
rect 4972 1764 5040 1810
rect 5086 1764 5108 1810
rect 4904 1696 5108 1764
rect 4904 1650 4926 1696
rect 4972 1650 5040 1696
rect 5086 1650 5108 1696
rect 4904 1582 5108 1650
rect 4904 1536 4926 1582
rect 4972 1536 5040 1582
rect 5086 1536 5108 1582
rect 4904 1468 5108 1536
rect 4904 1422 4926 1468
rect 4972 1422 5040 1468
rect 5086 1422 5108 1468
rect 4904 1354 5108 1422
rect 4904 1308 4926 1354
rect 4972 1308 5040 1354
rect 5086 1308 5108 1354
rect 4904 1240 5108 1308
rect 4904 1194 4926 1240
rect 4972 1194 5040 1240
rect 5086 1194 5108 1240
rect 4904 1126 5108 1194
rect 4904 1080 4926 1126
rect 4972 1080 5040 1126
rect 5086 1080 5108 1126
rect 4904 1012 5108 1080
rect 4904 966 4926 1012
rect 4972 966 5040 1012
rect 5086 966 5108 1012
rect 4904 898 5108 966
rect 4904 852 4926 898
rect 4972 852 5040 898
rect 5086 852 5108 898
rect 4904 784 5108 852
rect 4904 738 4926 784
rect 4972 738 5040 784
rect 5086 738 5108 784
rect 4904 328 5108 738
rect 10372 5572 10576 5640
rect 10372 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10576 5572
rect 10372 5458 10576 5526
rect 10372 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10576 5458
rect 10372 5344 10576 5412
rect 10372 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10576 5344
rect 10372 5230 10576 5298
rect 10372 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10576 5230
rect 10372 5116 10576 5184
rect 10372 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10576 5116
rect 10372 5002 10576 5070
rect 10372 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10576 5002
rect 10372 4888 10576 4956
rect 10372 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10576 4888
rect 10372 4774 10576 4842
rect 10372 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10576 4774
rect 10372 4660 10576 4728
rect 10372 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10576 4660
rect 10372 4546 10576 4614
rect 10372 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10576 4546
rect 10372 4432 10576 4500
rect 10372 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10576 4432
rect 10372 4318 10576 4386
rect 10372 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10576 4318
rect 10372 4204 10576 4272
rect 10372 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10576 4204
rect 10372 4090 10576 4158
rect 10372 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10576 4090
rect 10372 3976 10576 4044
rect 10372 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10576 3976
rect 10372 3862 10576 3930
rect 10372 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10576 3862
rect 10372 3748 10576 3816
rect 10372 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10576 3748
rect 10372 3634 10576 3702
rect 10372 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10576 3634
rect 10372 3520 10576 3588
rect 10372 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10576 3520
rect 10372 3406 10576 3474
rect 10372 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10576 3406
rect 10372 3292 10576 3360
rect 10372 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10576 3292
rect 10372 3178 10576 3246
rect 10372 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10576 3178
rect 10372 3064 10576 3132
rect 10372 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10576 3064
rect 10372 2950 10576 3018
rect 10372 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10576 2950
rect 10372 2836 10576 2904
rect 10372 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10576 2836
rect 10372 2722 10576 2790
rect 10372 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10576 2722
rect 10372 2608 10576 2676
rect 10372 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10576 2608
rect 10372 2494 10576 2562
rect 10372 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10576 2494
rect 10372 2380 10576 2448
rect 10372 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10576 2380
rect 10372 2266 10576 2334
rect 10372 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10576 2266
rect 10372 2152 10576 2220
rect 10372 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10576 2152
rect 10372 2038 10576 2106
rect 10372 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10576 2038
rect 10372 1924 10576 1992
rect 10372 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10576 1924
rect 10372 1810 10576 1878
rect 10372 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10576 1810
rect 10372 1696 10576 1764
rect 10372 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10576 1696
rect 10372 1582 10576 1650
rect 10372 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10576 1582
rect 10372 1468 10576 1536
rect 10372 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10576 1468
rect 10372 1354 10576 1422
rect 10372 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10576 1354
rect 10372 1240 10576 1308
rect 10372 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10576 1240
rect 10372 1126 10576 1194
rect 10372 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10576 1126
rect 10372 1012 10576 1080
rect 10372 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10576 1012
rect 10372 898 10576 966
rect 10372 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10576 898
rect 10372 784 10576 852
rect 10372 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10576 784
rect 10372 670 10576 738
rect 10372 624 10394 670
rect 10440 624 10508 670
rect 10554 624 10576 670
rect 10372 556 10576 624
rect 4904 282 4926 328
rect 4972 282 5040 328
rect 5086 282 5108 328
rect 4904 236 5108 282
rect 10372 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10576 556
rect 10372 442 10576 510
rect 10372 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10576 442
rect 10372 328 10576 396
rect 10372 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10576 328
rect 10372 236 10576 282
rect 4904 214 10576 236
rect 4904 168 4926 214
rect 4972 168 5040 214
rect 5086 168 5222 214
rect 5268 168 5336 214
rect 5382 168 5450 214
rect 5496 168 5564 214
rect 5610 168 5678 214
rect 5724 168 5792 214
rect 5838 168 5906 214
rect 5952 168 6020 214
rect 6066 168 6134 214
rect 6180 168 6248 214
rect 6294 168 6362 214
rect 6408 168 6476 214
rect 6522 168 6590 214
rect 6636 168 6704 214
rect 6750 168 6818 214
rect 6864 168 6932 214
rect 6978 168 7046 214
rect 7092 168 7160 214
rect 7206 168 7274 214
rect 7320 168 7388 214
rect 7434 168 7502 214
rect 7548 168 7616 214
rect 7662 168 7730 214
rect 7776 168 7844 214
rect 7890 168 7958 214
rect 8004 168 8072 214
rect 8118 168 8186 214
rect 8232 168 8300 214
rect 8346 168 8414 214
rect 8460 168 8528 214
rect 8574 168 8642 214
rect 8688 168 8756 214
rect 8802 168 8870 214
rect 8916 168 8984 214
rect 9030 168 9098 214
rect 9144 168 9212 214
rect 9258 168 9326 214
rect 9372 168 9440 214
rect 9486 168 9554 214
rect 9600 168 9668 214
rect 9714 168 9782 214
rect 9828 168 9896 214
rect 9942 168 10010 214
rect 10056 168 10124 214
rect 10170 168 10238 214
rect 10284 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10576 214
rect 4904 100 10576 168
rect 4904 54 4926 100
rect 4972 54 5040 100
rect 5086 54 5222 100
rect 5268 54 5336 100
rect 5382 54 5450 100
rect 5496 54 5564 100
rect 5610 54 5678 100
rect 5724 54 5792 100
rect 5838 54 5906 100
rect 5952 54 6020 100
rect 6066 54 6134 100
rect 6180 54 6248 100
rect 6294 54 6362 100
rect 6408 54 6476 100
rect 6522 54 6590 100
rect 6636 54 6704 100
rect 6750 54 6818 100
rect 6864 54 6932 100
rect 6978 54 7046 100
rect 7092 54 7160 100
rect 7206 54 7274 100
rect 7320 54 7388 100
rect 7434 54 7502 100
rect 7548 54 7616 100
rect 7662 54 7730 100
rect 7776 54 7844 100
rect 7890 54 7958 100
rect 8004 54 8072 100
rect 8118 54 8186 100
rect 8232 54 8300 100
rect 8346 54 8414 100
rect 8460 54 8528 100
rect 8574 54 8642 100
rect 8688 54 8756 100
rect 8802 54 8870 100
rect 8916 54 8984 100
rect 9030 54 9098 100
rect 9144 54 9212 100
rect 9258 54 9326 100
rect 9372 54 9440 100
rect 9486 54 9554 100
rect 9600 54 9668 100
rect 9714 54 9782 100
rect 9828 54 9896 100
rect 9942 54 10010 100
rect 10056 54 10124 100
rect 10170 54 10238 100
rect 10284 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10576 100
rect 4904 32 10576 54
<< psubdiffcont >>
rect 4926 12252 4972 12298
rect 5040 12252 5086 12298
rect 5217 12252 5263 12298
rect 5331 12252 5377 12298
rect 5445 12252 5491 12298
rect 5559 12252 5605 12298
rect 5673 12252 5719 12298
rect 5787 12252 5833 12298
rect 5901 12252 5947 12298
rect 6015 12252 6061 12298
rect 6129 12252 6175 12298
rect 6243 12252 6289 12298
rect 6357 12252 6403 12298
rect 6471 12252 6517 12298
rect 6585 12252 6631 12298
rect 6699 12252 6745 12298
rect 6813 12252 6859 12298
rect 6927 12252 6973 12298
rect 7041 12252 7087 12298
rect 7155 12252 7201 12298
rect 7269 12252 7315 12298
rect 7383 12252 7429 12298
rect 7497 12252 7543 12298
rect 7611 12252 7657 12298
rect 7725 12252 7771 12298
rect 7839 12252 7885 12298
rect 7953 12252 7999 12298
rect 8067 12252 8113 12298
rect 8181 12252 8227 12298
rect 8295 12252 8341 12298
rect 8409 12252 8455 12298
rect 8523 12252 8569 12298
rect 8637 12252 8683 12298
rect 8751 12252 8797 12298
rect 8865 12252 8911 12298
rect 8979 12252 9025 12298
rect 9093 12252 9139 12298
rect 9207 12252 9253 12298
rect 9321 12252 9367 12298
rect 9435 12252 9481 12298
rect 9549 12252 9595 12298
rect 9663 12252 9709 12298
rect 9777 12252 9823 12298
rect 9891 12252 9937 12298
rect 10005 12252 10051 12298
rect 10119 12252 10165 12298
rect 10233 12252 10279 12298
rect 10394 12252 10440 12298
rect 10508 12252 10554 12298
rect 4926 12138 4972 12184
rect 5040 12138 5086 12184
rect 5217 12138 5263 12184
rect 5331 12138 5377 12184
rect 5445 12138 5491 12184
rect 5559 12138 5605 12184
rect 5673 12138 5719 12184
rect 5787 12138 5833 12184
rect 5901 12138 5947 12184
rect 6015 12138 6061 12184
rect 6129 12138 6175 12184
rect 6243 12138 6289 12184
rect 6357 12138 6403 12184
rect 6471 12138 6517 12184
rect 6585 12138 6631 12184
rect 6699 12138 6745 12184
rect 6813 12138 6859 12184
rect 6927 12138 6973 12184
rect 7041 12138 7087 12184
rect 7155 12138 7201 12184
rect 7269 12138 7315 12184
rect 7383 12138 7429 12184
rect 7497 12138 7543 12184
rect 7611 12138 7657 12184
rect 7725 12138 7771 12184
rect 7839 12138 7885 12184
rect 7953 12138 7999 12184
rect 8067 12138 8113 12184
rect 8181 12138 8227 12184
rect 8295 12138 8341 12184
rect 8409 12138 8455 12184
rect 8523 12138 8569 12184
rect 8637 12138 8683 12184
rect 8751 12138 8797 12184
rect 8865 12138 8911 12184
rect 8979 12138 9025 12184
rect 9093 12138 9139 12184
rect 9207 12138 9253 12184
rect 9321 12138 9367 12184
rect 9435 12138 9481 12184
rect 9549 12138 9595 12184
rect 9663 12138 9709 12184
rect 9777 12138 9823 12184
rect 9891 12138 9937 12184
rect 10005 12138 10051 12184
rect 10119 12138 10165 12184
rect 10233 12138 10279 12184
rect 10394 12138 10440 12184
rect 10508 12138 10554 12184
rect 4926 12024 4972 12070
rect 5040 12024 5086 12070
rect 10394 12024 10440 12070
rect 10508 12024 10554 12070
rect 10394 11910 10440 11956
rect 10508 11910 10554 11956
rect 10394 11796 10440 11842
rect 10508 11796 10554 11842
rect 10394 11682 10440 11728
rect 10508 11682 10554 11728
rect 4926 11454 4972 11500
rect 5040 11454 5086 11500
rect 4926 11340 4972 11386
rect 5040 11340 5086 11386
rect 4926 11226 4972 11272
rect 5040 11226 5086 11272
rect 4926 11112 4972 11158
rect 5040 11112 5086 11158
rect 4926 10998 4972 11044
rect 5040 10998 5086 11044
rect 4926 10884 4972 10930
rect 5040 10884 5086 10930
rect 4926 10770 4972 10816
rect 5040 10770 5086 10816
rect 4926 10656 4972 10702
rect 5040 10656 5086 10702
rect 4926 10542 4972 10588
rect 5040 10542 5086 10588
rect 4926 10428 4972 10474
rect 5040 10428 5086 10474
rect 4926 10314 4972 10360
rect 5040 10314 5086 10360
rect 4926 10200 4972 10246
rect 5040 10200 5086 10246
rect 4926 10086 4972 10132
rect 5040 10086 5086 10132
rect 4926 9972 4972 10018
rect 5040 9972 5086 10018
rect 4926 9858 4972 9904
rect 5040 9858 5086 9904
rect 4926 9744 4972 9790
rect 5040 9744 5086 9790
rect 4926 9630 4972 9676
rect 5040 9630 5086 9676
rect 4926 9516 4972 9562
rect 5040 9516 5086 9562
rect 4926 9402 4972 9448
rect 5040 9402 5086 9448
rect 4926 9288 4972 9334
rect 5040 9288 5086 9334
rect 4926 9174 4972 9220
rect 5040 9174 5086 9220
rect 4926 9060 4972 9106
rect 5040 9060 5086 9106
rect 4926 8946 4972 8992
rect 5040 8946 5086 8992
rect 4926 8832 4972 8878
rect 5040 8832 5086 8878
rect 4926 8718 4972 8764
rect 5040 8718 5086 8764
rect 4926 8604 4972 8650
rect 5040 8604 5086 8650
rect 4926 8490 4972 8536
rect 5040 8490 5086 8536
rect 4926 8376 4972 8422
rect 5040 8376 5086 8422
rect 4926 8262 4972 8308
rect 5040 8262 5086 8308
rect 4926 8148 4972 8194
rect 5040 8148 5086 8194
rect 4926 8034 4972 8080
rect 5040 8034 5086 8080
rect 4926 7920 4972 7966
rect 5040 7920 5086 7966
rect 4926 7806 4972 7852
rect 5040 7806 5086 7852
rect 4926 7692 4972 7738
rect 5040 7692 5086 7738
rect 4926 7578 4972 7624
rect 5040 7578 5086 7624
rect 4926 7464 4972 7510
rect 5040 7464 5086 7510
rect 4926 7350 4972 7396
rect 5040 7350 5086 7396
rect 4926 7236 4972 7282
rect 5040 7236 5086 7282
rect 4926 7122 4972 7168
rect 5040 7122 5086 7168
rect 4926 7008 4972 7054
rect 5040 7008 5086 7054
rect 4926 6894 4972 6940
rect 5040 6894 5086 6940
rect 4926 6780 4972 6826
rect 5040 6780 5086 6826
rect 4926 6666 4972 6712
rect 5040 6666 5086 6712
rect 10394 11568 10440 11614
rect 10508 11568 10554 11614
rect 10394 11454 10440 11500
rect 10508 11454 10554 11500
rect 10394 11340 10440 11386
rect 10508 11340 10554 11386
rect 10394 11226 10440 11272
rect 10508 11226 10554 11272
rect 10394 11112 10440 11158
rect 10508 11112 10554 11158
rect 10394 10998 10440 11044
rect 10508 10998 10554 11044
rect 10394 10884 10440 10930
rect 10508 10884 10554 10930
rect 10394 10770 10440 10816
rect 10508 10770 10554 10816
rect 10394 10656 10440 10702
rect 10508 10656 10554 10702
rect 10394 10542 10440 10588
rect 10508 10542 10554 10588
rect 10394 10428 10440 10474
rect 10508 10428 10554 10474
rect 10394 10314 10440 10360
rect 10508 10314 10554 10360
rect 10394 10200 10440 10246
rect 10508 10200 10554 10246
rect 10394 10086 10440 10132
rect 10508 10086 10554 10132
rect 10394 9972 10440 10018
rect 10508 9972 10554 10018
rect 10394 9858 10440 9904
rect 10508 9858 10554 9904
rect 10394 9744 10440 9790
rect 10508 9744 10554 9790
rect 10394 9630 10440 9676
rect 10508 9630 10554 9676
rect 10394 9516 10440 9562
rect 10508 9516 10554 9562
rect 10394 9402 10440 9448
rect 10508 9402 10554 9448
rect 10394 9288 10440 9334
rect 10508 9288 10554 9334
rect 10394 9174 10440 9220
rect 10508 9174 10554 9220
rect 10394 9060 10440 9106
rect 10508 9060 10554 9106
rect 10394 8946 10440 8992
rect 10508 8946 10554 8992
rect 10394 8832 10440 8878
rect 10508 8832 10554 8878
rect 10394 8718 10440 8764
rect 10508 8718 10554 8764
rect 10394 8604 10440 8650
rect 10508 8604 10554 8650
rect 10394 8490 10440 8536
rect 10508 8490 10554 8536
rect 10394 8376 10440 8422
rect 10508 8376 10554 8422
rect 10394 8262 10440 8308
rect 10508 8262 10554 8308
rect 10394 8148 10440 8194
rect 10508 8148 10554 8194
rect 10394 8034 10440 8080
rect 10508 8034 10554 8080
rect 10394 7920 10440 7966
rect 10508 7920 10554 7966
rect 10394 7806 10440 7852
rect 10508 7806 10554 7852
rect 10394 7692 10440 7738
rect 10508 7692 10554 7738
rect 10394 7578 10440 7624
rect 10508 7578 10554 7624
rect 10394 7464 10440 7510
rect 10508 7464 10554 7510
rect 10394 7350 10440 7396
rect 10508 7350 10554 7396
rect 10394 7236 10440 7282
rect 10508 7236 10554 7282
rect 10394 7122 10440 7168
rect 10508 7122 10554 7168
rect 10394 7008 10440 7054
rect 10508 7008 10554 7054
rect 10394 6894 10440 6940
rect 10508 6894 10554 6940
rect 10394 6780 10440 6826
rect 10508 6780 10554 6826
rect 10394 6666 10440 6712
rect 10508 6666 10554 6712
rect 4926 6552 4972 6598
rect 5040 6552 5086 6598
rect 10394 6552 10440 6598
rect 10508 6552 10554 6598
rect 4926 6438 4972 6484
rect 5040 6438 5086 6484
rect 4926 6324 4972 6370
rect 5040 6324 5086 6370
rect 4926 6210 4972 6256
rect 5040 6210 5086 6256
rect 10394 6438 10440 6484
rect 10508 6438 10554 6484
rect 10394 6324 10440 6370
rect 10508 6324 10554 6370
rect 10394 6210 10440 6256
rect 10508 6210 10554 6256
rect 5214 6161 5260 6207
rect 5328 6161 5374 6207
rect 5442 6161 5488 6207
rect 5556 6161 5602 6207
rect 5670 6161 5716 6207
rect 5784 6161 5830 6207
rect 5898 6161 5944 6207
rect 6012 6161 6058 6207
rect 6126 6161 6172 6207
rect 6240 6161 6286 6207
rect 6354 6161 6400 6207
rect 6468 6161 6514 6207
rect 6582 6161 6628 6207
rect 6696 6161 6742 6207
rect 6810 6161 6856 6207
rect 6924 6161 6970 6207
rect 7038 6161 7084 6207
rect 7152 6161 7198 6207
rect 7266 6161 7312 6207
rect 7380 6161 7426 6207
rect 7494 6161 7540 6207
rect 7608 6161 7654 6207
rect 7722 6161 7768 6207
rect 7836 6161 7882 6207
rect 7950 6161 7996 6207
rect 8064 6161 8110 6207
rect 8178 6161 8224 6207
rect 8292 6161 8338 6207
rect 8406 6161 8452 6207
rect 8520 6161 8566 6207
rect 8634 6161 8680 6207
rect 8748 6161 8794 6207
rect 8862 6161 8908 6207
rect 8976 6161 9022 6207
rect 9090 6161 9136 6207
rect 9204 6161 9250 6207
rect 9318 6161 9364 6207
rect 9432 6161 9478 6207
rect 9546 6161 9592 6207
rect 9660 6161 9706 6207
rect 9774 6161 9820 6207
rect 9888 6161 9934 6207
rect 10002 6161 10048 6207
rect 10116 6161 10162 6207
rect 10230 6161 10276 6207
rect 4926 6096 4972 6142
rect 5040 6096 5086 6142
rect 10394 6096 10440 6142
rect 10508 6096 10554 6142
rect 5214 6047 5260 6093
rect 5328 6047 5374 6093
rect 5442 6047 5488 6093
rect 5556 6047 5602 6093
rect 5670 6047 5716 6093
rect 5784 6047 5830 6093
rect 5898 6047 5944 6093
rect 6012 6047 6058 6093
rect 6126 6047 6172 6093
rect 6240 6047 6286 6093
rect 6354 6047 6400 6093
rect 6468 6047 6514 6093
rect 6582 6047 6628 6093
rect 6696 6047 6742 6093
rect 6810 6047 6856 6093
rect 6924 6047 6970 6093
rect 7038 6047 7084 6093
rect 7152 6047 7198 6093
rect 7266 6047 7312 6093
rect 7380 6047 7426 6093
rect 7494 6047 7540 6093
rect 7608 6047 7654 6093
rect 7722 6047 7768 6093
rect 7836 6047 7882 6093
rect 7950 6047 7996 6093
rect 8064 6047 8110 6093
rect 8178 6047 8224 6093
rect 8292 6047 8338 6093
rect 8406 6047 8452 6093
rect 8520 6047 8566 6093
rect 8634 6047 8680 6093
rect 8748 6047 8794 6093
rect 8862 6047 8908 6093
rect 8976 6047 9022 6093
rect 9090 6047 9136 6093
rect 9204 6047 9250 6093
rect 9318 6047 9364 6093
rect 9432 6047 9478 6093
rect 9546 6047 9592 6093
rect 9660 6047 9706 6093
rect 9774 6047 9820 6093
rect 9888 6047 9934 6093
rect 10002 6047 10048 6093
rect 10116 6047 10162 6093
rect 10230 6047 10276 6093
rect 4926 5982 4972 6028
rect 5040 5982 5086 6028
rect 4926 5868 4972 5914
rect 5040 5868 5086 5914
rect 4926 5754 4972 5800
rect 5040 5754 5086 5800
rect 10394 5982 10440 6028
rect 10508 5982 10554 6028
rect 10394 5868 10440 5914
rect 10508 5868 10554 5914
rect 10394 5754 10440 5800
rect 10508 5754 10554 5800
rect 4926 5640 4972 5686
rect 5040 5640 5086 5686
rect 10394 5640 10440 5686
rect 10508 5640 10554 5686
rect 4926 5526 4972 5572
rect 5040 5526 5086 5572
rect 4926 5412 4972 5458
rect 5040 5412 5086 5458
rect 4926 5298 4972 5344
rect 5040 5298 5086 5344
rect 4926 5184 4972 5230
rect 5040 5184 5086 5230
rect 4926 5070 4972 5116
rect 5040 5070 5086 5116
rect 4926 4956 4972 5002
rect 5040 4956 5086 5002
rect 4926 4842 4972 4888
rect 5040 4842 5086 4888
rect 4926 4728 4972 4774
rect 5040 4728 5086 4774
rect 4926 4614 4972 4660
rect 5040 4614 5086 4660
rect 4926 4500 4972 4546
rect 5040 4500 5086 4546
rect 4926 4386 4972 4432
rect 5040 4386 5086 4432
rect 4926 4272 4972 4318
rect 5040 4272 5086 4318
rect 4926 4158 4972 4204
rect 5040 4158 5086 4204
rect 4926 4044 4972 4090
rect 5040 4044 5086 4090
rect 4926 3930 4972 3976
rect 5040 3930 5086 3976
rect 4926 3816 4972 3862
rect 5040 3816 5086 3862
rect 4926 3702 4972 3748
rect 5040 3702 5086 3748
rect 4926 3588 4972 3634
rect 5040 3588 5086 3634
rect 4926 3474 4972 3520
rect 5040 3474 5086 3520
rect 4926 3360 4972 3406
rect 5040 3360 5086 3406
rect 4926 3246 4972 3292
rect 5040 3246 5086 3292
rect 4926 3132 4972 3178
rect 5040 3132 5086 3178
rect 4926 3018 4972 3064
rect 5040 3018 5086 3064
rect 4926 2904 4972 2950
rect 5040 2904 5086 2950
rect 4926 2790 4972 2836
rect 5040 2790 5086 2836
rect 4926 2676 4972 2722
rect 5040 2676 5086 2722
rect 4926 2562 4972 2608
rect 5040 2562 5086 2608
rect 4926 2448 4972 2494
rect 5040 2448 5086 2494
rect 4926 2334 4972 2380
rect 5040 2334 5086 2380
rect 4926 2220 4972 2266
rect 5040 2220 5086 2266
rect 4926 2106 4972 2152
rect 5040 2106 5086 2152
rect 4926 1992 4972 2038
rect 5040 1992 5086 2038
rect 4926 1878 4972 1924
rect 5040 1878 5086 1924
rect 4926 1764 4972 1810
rect 5040 1764 5086 1810
rect 4926 1650 4972 1696
rect 5040 1650 5086 1696
rect 4926 1536 4972 1582
rect 5040 1536 5086 1582
rect 4926 1422 4972 1468
rect 5040 1422 5086 1468
rect 4926 1308 4972 1354
rect 5040 1308 5086 1354
rect 4926 1194 4972 1240
rect 5040 1194 5086 1240
rect 4926 1080 4972 1126
rect 5040 1080 5086 1126
rect 4926 966 4972 1012
rect 5040 966 5086 1012
rect 4926 852 4972 898
rect 5040 852 5086 898
rect 4926 738 4972 784
rect 5040 738 5086 784
rect 10394 5526 10440 5572
rect 10508 5526 10554 5572
rect 10394 5412 10440 5458
rect 10508 5412 10554 5458
rect 10394 5298 10440 5344
rect 10508 5298 10554 5344
rect 10394 5184 10440 5230
rect 10508 5184 10554 5230
rect 10394 5070 10440 5116
rect 10508 5070 10554 5116
rect 10394 4956 10440 5002
rect 10508 4956 10554 5002
rect 10394 4842 10440 4888
rect 10508 4842 10554 4888
rect 10394 4728 10440 4774
rect 10508 4728 10554 4774
rect 10394 4614 10440 4660
rect 10508 4614 10554 4660
rect 10394 4500 10440 4546
rect 10508 4500 10554 4546
rect 10394 4386 10440 4432
rect 10508 4386 10554 4432
rect 10394 4272 10440 4318
rect 10508 4272 10554 4318
rect 10394 4158 10440 4204
rect 10508 4158 10554 4204
rect 10394 4044 10440 4090
rect 10508 4044 10554 4090
rect 10394 3930 10440 3976
rect 10508 3930 10554 3976
rect 10394 3816 10440 3862
rect 10508 3816 10554 3862
rect 10394 3702 10440 3748
rect 10508 3702 10554 3748
rect 10394 3588 10440 3634
rect 10508 3588 10554 3634
rect 10394 3474 10440 3520
rect 10508 3474 10554 3520
rect 10394 3360 10440 3406
rect 10508 3360 10554 3406
rect 10394 3246 10440 3292
rect 10508 3246 10554 3292
rect 10394 3132 10440 3178
rect 10508 3132 10554 3178
rect 10394 3018 10440 3064
rect 10508 3018 10554 3064
rect 10394 2904 10440 2950
rect 10508 2904 10554 2950
rect 10394 2790 10440 2836
rect 10508 2790 10554 2836
rect 10394 2676 10440 2722
rect 10508 2676 10554 2722
rect 10394 2562 10440 2608
rect 10508 2562 10554 2608
rect 10394 2448 10440 2494
rect 10508 2448 10554 2494
rect 10394 2334 10440 2380
rect 10508 2334 10554 2380
rect 10394 2220 10440 2266
rect 10508 2220 10554 2266
rect 10394 2106 10440 2152
rect 10508 2106 10554 2152
rect 10394 1992 10440 2038
rect 10508 1992 10554 2038
rect 10394 1878 10440 1924
rect 10508 1878 10554 1924
rect 10394 1764 10440 1810
rect 10508 1764 10554 1810
rect 10394 1650 10440 1696
rect 10508 1650 10554 1696
rect 10394 1536 10440 1582
rect 10508 1536 10554 1582
rect 10394 1422 10440 1468
rect 10508 1422 10554 1468
rect 10394 1308 10440 1354
rect 10508 1308 10554 1354
rect 10394 1194 10440 1240
rect 10508 1194 10554 1240
rect 10394 1080 10440 1126
rect 10508 1080 10554 1126
rect 10394 966 10440 1012
rect 10508 966 10554 1012
rect 10394 852 10440 898
rect 10508 852 10554 898
rect 10394 738 10440 784
rect 10508 738 10554 784
rect 10394 624 10440 670
rect 10508 624 10554 670
rect 4926 282 4972 328
rect 5040 282 5086 328
rect 10394 510 10440 556
rect 10508 510 10554 556
rect 10394 396 10440 442
rect 10508 396 10554 442
rect 10394 282 10440 328
rect 10508 282 10554 328
rect 4926 168 4972 214
rect 5040 168 5086 214
rect 5222 168 5268 214
rect 5336 168 5382 214
rect 5450 168 5496 214
rect 5564 168 5610 214
rect 5678 168 5724 214
rect 5792 168 5838 214
rect 5906 168 5952 214
rect 6020 168 6066 214
rect 6134 168 6180 214
rect 6248 168 6294 214
rect 6362 168 6408 214
rect 6476 168 6522 214
rect 6590 168 6636 214
rect 6704 168 6750 214
rect 6818 168 6864 214
rect 6932 168 6978 214
rect 7046 168 7092 214
rect 7160 168 7206 214
rect 7274 168 7320 214
rect 7388 168 7434 214
rect 7502 168 7548 214
rect 7616 168 7662 214
rect 7730 168 7776 214
rect 7844 168 7890 214
rect 7958 168 8004 214
rect 8072 168 8118 214
rect 8186 168 8232 214
rect 8300 168 8346 214
rect 8414 168 8460 214
rect 8528 168 8574 214
rect 8642 168 8688 214
rect 8756 168 8802 214
rect 8870 168 8916 214
rect 8984 168 9030 214
rect 9098 168 9144 214
rect 9212 168 9258 214
rect 9326 168 9372 214
rect 9440 168 9486 214
rect 9554 168 9600 214
rect 9668 168 9714 214
rect 9782 168 9828 214
rect 9896 168 9942 214
rect 10010 168 10056 214
rect 10124 168 10170 214
rect 10238 168 10284 214
rect 10394 168 10440 214
rect 10508 168 10554 214
rect 4926 54 4972 100
rect 5040 54 5086 100
rect 5222 54 5268 100
rect 5336 54 5382 100
rect 5450 54 5496 100
rect 5564 54 5610 100
rect 5678 54 5724 100
rect 5792 54 5838 100
rect 5906 54 5952 100
rect 6020 54 6066 100
rect 6134 54 6180 100
rect 6248 54 6294 100
rect 6362 54 6408 100
rect 6476 54 6522 100
rect 6590 54 6636 100
rect 6704 54 6750 100
rect 6818 54 6864 100
rect 6932 54 6978 100
rect 7046 54 7092 100
rect 7160 54 7206 100
rect 7274 54 7320 100
rect 7388 54 7434 100
rect 7502 54 7548 100
rect 7616 54 7662 100
rect 7730 54 7776 100
rect 7844 54 7890 100
rect 7958 54 8004 100
rect 8072 54 8118 100
rect 8186 54 8232 100
rect 8300 54 8346 100
rect 8414 54 8460 100
rect 8528 54 8574 100
rect 8642 54 8688 100
rect 8756 54 8802 100
rect 8870 54 8916 100
rect 8984 54 9030 100
rect 9098 54 9144 100
rect 9212 54 9258 100
rect 9326 54 9372 100
rect 9440 54 9486 100
rect 9554 54 9600 100
rect 9668 54 9714 100
rect 9782 54 9828 100
rect 9896 54 9942 100
rect 10010 54 10056 100
rect 10124 54 10170 100
rect 10238 54 10284 100
rect 10394 54 10440 100
rect 10508 54 10554 100
<< mvnmoscap >>
rect 5519 6633 7519 11633
rect 7955 6633 9955 11633
rect 5519 621 7519 5621
rect 7955 621 9955 5621
<< polysilicon >>
rect 5519 11712 7519 11725
rect 5519 11666 5572 11712
rect 7466 11666 7519 11712
rect 5519 11633 7519 11666
rect 7955 11712 9955 11725
rect 7955 11666 8008 11712
rect 9902 11666 9955 11712
rect 7955 11633 9955 11666
rect 5519 6600 7519 6633
rect 5519 6554 5572 6600
rect 7466 6554 7519 6600
rect 5519 6541 7519 6554
rect 7955 6600 9955 6633
rect 7955 6554 8008 6600
rect 9902 6554 9955 6600
rect 7955 6541 9955 6554
rect 5519 5700 7519 5713
rect 5519 5654 5572 5700
rect 7466 5654 7519 5700
rect 5519 5621 7519 5654
rect 7955 5700 9955 5713
rect 7955 5654 8008 5700
rect 9902 5654 9955 5700
rect 7955 5621 9955 5654
rect 5519 588 7519 621
rect 5519 542 5572 588
rect 7466 542 7519 588
rect 5519 529 7519 542
rect 7955 588 9955 621
rect 7955 542 8008 588
rect 9902 542 9955 588
rect 7955 529 9955 542
<< polycontact >>
rect 5572 11666 7466 11712
rect 8008 11666 9902 11712
rect 5572 6554 7466 6600
rect 8008 6554 9902 6600
rect 5572 5654 7466 5700
rect 8008 5654 9902 5700
rect 5572 542 7466 588
rect 8008 542 9902 588
<< metal1 >>
rect 4915 12298 10565 12310
rect 4915 12252 4926 12298
rect 4972 12252 5040 12298
rect 5086 12252 5217 12298
rect 5263 12252 5331 12298
rect 5377 12252 5445 12298
rect 5491 12252 5559 12298
rect 5605 12252 5673 12298
rect 5719 12252 5787 12298
rect 5833 12252 5901 12298
rect 5947 12252 6015 12298
rect 6061 12252 6129 12298
rect 6175 12252 6243 12298
rect 6289 12252 6357 12298
rect 6403 12252 6471 12298
rect 6517 12252 6585 12298
rect 6631 12252 6699 12298
rect 6745 12252 6813 12298
rect 6859 12252 6927 12298
rect 6973 12252 7041 12298
rect 7087 12252 7155 12298
rect 7201 12252 7269 12298
rect 7315 12252 7383 12298
rect 7429 12252 7497 12298
rect 7543 12252 7611 12298
rect 7657 12252 7725 12298
rect 7771 12252 7839 12298
rect 7885 12252 7953 12298
rect 7999 12252 8067 12298
rect 8113 12252 8181 12298
rect 8227 12252 8295 12298
rect 8341 12252 8409 12298
rect 8455 12252 8523 12298
rect 8569 12252 8637 12298
rect 8683 12252 8751 12298
rect 8797 12252 8865 12298
rect 8911 12252 8979 12298
rect 9025 12252 9093 12298
rect 9139 12252 9207 12298
rect 9253 12252 9321 12298
rect 9367 12252 9435 12298
rect 9481 12252 9549 12298
rect 9595 12252 9663 12298
rect 9709 12252 9777 12298
rect 9823 12252 9891 12298
rect 9937 12252 10005 12298
rect 10051 12252 10119 12298
rect 10165 12252 10233 12298
rect 10279 12252 10394 12298
rect 10440 12252 10508 12298
rect 10554 12252 10565 12298
rect 4915 12184 10565 12252
rect 4915 12138 4926 12184
rect 4972 12138 5040 12184
rect 5086 12138 5217 12184
rect 5263 12138 5331 12184
rect 5377 12138 5445 12184
rect 5491 12138 5559 12184
rect 5605 12138 5673 12184
rect 5719 12138 5787 12184
rect 5833 12138 5901 12184
rect 5947 12138 6015 12184
rect 6061 12138 6129 12184
rect 6175 12138 6243 12184
rect 6289 12138 6357 12184
rect 6403 12138 6471 12184
rect 6517 12138 6585 12184
rect 6631 12138 6699 12184
rect 6745 12138 6813 12184
rect 6859 12138 6927 12184
rect 6973 12138 7041 12184
rect 7087 12138 7155 12184
rect 7201 12138 7269 12184
rect 7315 12138 7383 12184
rect 7429 12138 7497 12184
rect 7543 12138 7611 12184
rect 7657 12138 7725 12184
rect 7771 12138 7839 12184
rect 7885 12138 7953 12184
rect 7999 12138 8067 12184
rect 8113 12138 8181 12184
rect 8227 12138 8295 12184
rect 8341 12138 8409 12184
rect 8455 12138 8523 12184
rect 8569 12138 8637 12184
rect 8683 12138 8751 12184
rect 8797 12138 8865 12184
rect 8911 12138 8979 12184
rect 9025 12138 9093 12184
rect 9139 12138 9207 12184
rect 9253 12138 9321 12184
rect 9367 12138 9435 12184
rect 9481 12138 9549 12184
rect 9595 12138 9663 12184
rect 9709 12138 9777 12184
rect 9823 12138 9891 12184
rect 9937 12138 10005 12184
rect 10051 12138 10119 12184
rect 10165 12138 10233 12184
rect 10279 12138 10394 12184
rect 10440 12138 10508 12184
rect 10554 12138 10565 12184
rect 4915 12126 10565 12138
rect 4915 12070 5097 12126
rect 4915 12024 4926 12070
rect 4972 12024 5040 12070
rect 5086 12024 5097 12070
rect 4915 11633 5097 12024
rect 10383 12070 10565 12126
rect 10383 12024 10394 12070
rect 10440 12024 10508 12070
rect 10554 12024 10565 12070
rect 10383 11956 10565 12024
rect 10383 11910 10394 11956
rect 10440 11910 10508 11956
rect 10554 11910 10565 11956
rect 5561 11723 9913 11855
rect 5561 11712 7477 11723
rect 5561 11666 5572 11712
rect 7466 11666 7477 11712
rect 5561 11655 7477 11666
rect 7997 11712 9913 11723
rect 7997 11666 8008 11712
rect 9902 11666 9913 11712
rect 7997 11655 9913 11666
rect 10383 11842 10565 11910
rect 10383 11796 10394 11842
rect 10440 11796 10508 11842
rect 10554 11796 10565 11842
rect 10383 11728 10565 11796
rect 10383 11682 10394 11728
rect 10440 11682 10508 11728
rect 10554 11682 10565 11728
rect 4915 11596 5501 11633
rect 4915 11500 5444 11596
rect 4915 11454 4926 11500
rect 4972 11454 5040 11500
rect 5086 11454 5444 11500
rect 4915 11386 5444 11454
rect 4915 11340 4926 11386
rect 4972 11340 5040 11386
rect 5086 11340 5444 11386
rect 4915 11272 5444 11340
rect 4915 11226 4926 11272
rect 4972 11226 5040 11272
rect 5086 11226 5444 11272
rect 4915 11158 5444 11226
rect 4915 11112 4926 11158
rect 4972 11112 5040 11158
rect 5086 11112 5444 11158
rect 4915 11044 5444 11112
rect 4915 10998 4926 11044
rect 4972 10998 5040 11044
rect 5086 10998 5444 11044
rect 4915 10930 5444 10998
rect 4915 10884 4926 10930
rect 4972 10884 5040 10930
rect 5086 10884 5444 10930
rect 4915 10816 5444 10884
rect 4915 10770 4926 10816
rect 4972 10770 5040 10816
rect 5086 10770 5444 10816
rect 4915 10702 5444 10770
rect 4915 10656 4926 10702
rect 4972 10656 5040 10702
rect 5086 10656 5444 10702
rect 4915 10588 5444 10656
rect 4915 10542 4926 10588
rect 4972 10542 5040 10588
rect 5086 10542 5444 10588
rect 4915 10474 5444 10542
rect 4915 10428 4926 10474
rect 4972 10428 5040 10474
rect 5086 10428 5444 10474
rect 4915 10360 5444 10428
rect 4915 10314 4926 10360
rect 4972 10314 5040 10360
rect 5086 10314 5444 10360
rect 4915 10246 5444 10314
rect 4915 10200 4926 10246
rect 4972 10200 5040 10246
rect 5086 10200 5444 10246
rect 4915 10132 5444 10200
rect 4915 10086 4926 10132
rect 4972 10086 5040 10132
rect 5086 10086 5444 10132
rect 4915 10018 5444 10086
rect 4915 9972 4926 10018
rect 4972 9972 5040 10018
rect 5086 9972 5444 10018
rect 4915 9904 5444 9972
rect 4915 9858 4926 9904
rect 4972 9858 5040 9904
rect 5086 9858 5444 9904
rect 4915 9790 5444 9858
rect 4915 9744 4926 9790
rect 4972 9744 5040 9790
rect 5086 9744 5444 9790
rect 4915 9676 5444 9744
rect 4915 9630 4926 9676
rect 4972 9630 5040 9676
rect 5086 9630 5444 9676
rect 4915 9562 5444 9630
rect 4915 9516 4926 9562
rect 4972 9516 5040 9562
rect 5086 9516 5444 9562
rect 4915 9448 5444 9516
rect 4915 9402 4926 9448
rect 4972 9402 5040 9448
rect 5086 9402 5444 9448
rect 4915 9334 5444 9402
rect 4915 9288 4926 9334
rect 4972 9288 5040 9334
rect 5086 9288 5444 9334
rect 4915 9220 5444 9288
rect 4915 9174 4926 9220
rect 4972 9174 5040 9220
rect 5086 9174 5444 9220
rect 4915 9106 5444 9174
rect 4915 9060 4926 9106
rect 4972 9060 5040 9106
rect 5086 9060 5444 9106
rect 4915 8992 5444 9060
rect 4915 8946 4926 8992
rect 4972 8946 5040 8992
rect 5086 8946 5444 8992
rect 4915 8878 5444 8946
rect 4915 8832 4926 8878
rect 4972 8832 5040 8878
rect 5086 8832 5444 8878
rect 4915 8764 5444 8832
rect 4915 8718 4926 8764
rect 4972 8718 5040 8764
rect 5086 8718 5444 8764
rect 4915 8650 5444 8718
rect 4915 8604 4926 8650
rect 4972 8604 5040 8650
rect 5086 8604 5444 8650
rect 4915 8536 5444 8604
rect 4915 8490 4926 8536
rect 4972 8490 5040 8536
rect 5086 8490 5444 8536
rect 4915 8422 5444 8490
rect 4915 8376 4926 8422
rect 4972 8376 5040 8422
rect 5086 8376 5444 8422
rect 4915 8308 5444 8376
rect 4915 8262 4926 8308
rect 4972 8262 5040 8308
rect 5086 8262 5444 8308
rect 4915 8194 5444 8262
rect 4915 8148 4926 8194
rect 4972 8148 5040 8194
rect 5086 8148 5444 8194
rect 4915 8080 5444 8148
rect 4915 8034 4926 8080
rect 4972 8034 5040 8080
rect 5086 8034 5444 8080
rect 4915 7966 5444 8034
rect 4915 7920 4926 7966
rect 4972 7920 5040 7966
rect 5086 7920 5444 7966
rect 4915 7852 5444 7920
rect 4915 7806 4926 7852
rect 4972 7806 5040 7852
rect 5086 7806 5444 7852
rect 4915 7738 5444 7806
rect 4915 7692 4926 7738
rect 4972 7692 5040 7738
rect 5086 7692 5444 7738
rect 4915 7624 5444 7692
rect 4915 7578 4926 7624
rect 4972 7578 5040 7624
rect 5086 7578 5444 7624
rect 4915 7510 5444 7578
rect 4915 7464 4926 7510
rect 4972 7464 5040 7510
rect 5086 7464 5444 7510
rect 4915 7396 5444 7464
rect 4915 7350 4926 7396
rect 4972 7350 5040 7396
rect 5086 7350 5444 7396
rect 4915 7282 5444 7350
rect 4915 7236 4926 7282
rect 4972 7236 5040 7282
rect 5086 7236 5444 7282
rect 4915 7168 5444 7236
rect 4915 7122 4926 7168
rect 4972 7122 5040 7168
rect 5086 7122 5444 7168
rect 4915 7054 5444 7122
rect 4915 7008 4926 7054
rect 4972 7008 5040 7054
rect 5086 7008 5444 7054
rect 4915 6940 5444 7008
rect 4915 6894 4926 6940
rect 4972 6894 5040 6940
rect 5086 6894 5444 6940
rect 4915 6826 5444 6894
rect 4915 6780 4926 6826
rect 4972 6780 5040 6826
rect 5086 6780 5444 6826
rect 4915 6712 5444 6780
rect 4915 6666 4926 6712
rect 4972 6666 5040 6712
rect 5086 6670 5444 6712
rect 5490 6670 5501 11596
rect 5086 6666 5501 6670
rect 4915 6598 5501 6666
rect 6019 6611 7019 11655
rect 7537 11596 7937 11633
rect 7537 6670 7548 11596
rect 7594 6670 7880 11596
rect 7926 6670 7937 11596
rect 4915 6552 4926 6598
rect 4972 6552 5040 6598
rect 5086 6552 5501 6598
rect 4915 6484 5501 6552
rect 5561 6600 7477 6611
rect 5561 6554 5572 6600
rect 7466 6554 7477 6600
rect 5561 6543 7477 6554
rect 4915 6438 4926 6484
rect 4972 6438 5040 6484
rect 5086 6483 5501 6484
rect 7537 6483 7937 6670
rect 8455 6611 9455 11655
rect 10383 11633 10565 11682
rect 9973 11614 10565 11633
rect 9973 11596 10394 11614
rect 9973 6670 9984 11596
rect 10030 11568 10394 11596
rect 10440 11568 10508 11614
rect 10554 11568 10565 11614
rect 10030 11500 10565 11568
rect 10030 11454 10394 11500
rect 10440 11454 10508 11500
rect 10554 11454 10565 11500
rect 10030 11386 10565 11454
rect 10030 11340 10394 11386
rect 10440 11340 10508 11386
rect 10554 11340 10565 11386
rect 10030 11272 10565 11340
rect 10030 11226 10394 11272
rect 10440 11226 10508 11272
rect 10554 11226 10565 11272
rect 10030 11158 10565 11226
rect 10030 11112 10394 11158
rect 10440 11112 10508 11158
rect 10554 11112 10565 11158
rect 10030 11044 10565 11112
rect 10030 10998 10394 11044
rect 10440 10998 10508 11044
rect 10554 10998 10565 11044
rect 10030 10930 10565 10998
rect 10030 10884 10394 10930
rect 10440 10884 10508 10930
rect 10554 10884 10565 10930
rect 10030 10816 10565 10884
rect 10030 10770 10394 10816
rect 10440 10770 10508 10816
rect 10554 10770 10565 10816
rect 10030 10702 10565 10770
rect 10030 10656 10394 10702
rect 10440 10656 10508 10702
rect 10554 10656 10565 10702
rect 10030 10588 10565 10656
rect 10030 10542 10394 10588
rect 10440 10542 10508 10588
rect 10554 10542 10565 10588
rect 10030 10474 10565 10542
rect 10030 10428 10394 10474
rect 10440 10428 10508 10474
rect 10554 10428 10565 10474
rect 10030 10360 10565 10428
rect 10030 10314 10394 10360
rect 10440 10314 10508 10360
rect 10554 10314 10565 10360
rect 10030 10246 10565 10314
rect 10030 10200 10394 10246
rect 10440 10200 10508 10246
rect 10554 10200 10565 10246
rect 10030 10132 10565 10200
rect 10030 10086 10394 10132
rect 10440 10086 10508 10132
rect 10554 10086 10565 10132
rect 10030 10018 10565 10086
rect 10030 9972 10394 10018
rect 10440 9972 10508 10018
rect 10554 9972 10565 10018
rect 10030 9904 10565 9972
rect 10030 9858 10394 9904
rect 10440 9858 10508 9904
rect 10554 9858 10565 9904
rect 10030 9790 10565 9858
rect 10030 9744 10394 9790
rect 10440 9744 10508 9790
rect 10554 9744 10565 9790
rect 10030 9676 10565 9744
rect 10030 9630 10394 9676
rect 10440 9630 10508 9676
rect 10554 9630 10565 9676
rect 10030 9562 10565 9630
rect 10030 9516 10394 9562
rect 10440 9516 10508 9562
rect 10554 9516 10565 9562
rect 10030 9448 10565 9516
rect 10030 9402 10394 9448
rect 10440 9402 10508 9448
rect 10554 9402 10565 9448
rect 10030 9334 10565 9402
rect 10030 9288 10394 9334
rect 10440 9288 10508 9334
rect 10554 9288 10565 9334
rect 10030 9220 10565 9288
rect 10030 9174 10394 9220
rect 10440 9174 10508 9220
rect 10554 9174 10565 9220
rect 10030 9106 10565 9174
rect 10030 9060 10394 9106
rect 10440 9060 10508 9106
rect 10554 9060 10565 9106
rect 10030 8992 10565 9060
rect 10030 8946 10394 8992
rect 10440 8946 10508 8992
rect 10554 8946 10565 8992
rect 10030 8878 10565 8946
rect 10030 8832 10394 8878
rect 10440 8832 10508 8878
rect 10554 8832 10565 8878
rect 10030 8764 10565 8832
rect 10030 8718 10394 8764
rect 10440 8718 10508 8764
rect 10554 8718 10565 8764
rect 10030 8650 10565 8718
rect 10030 8604 10394 8650
rect 10440 8604 10508 8650
rect 10554 8604 10565 8650
rect 10030 8536 10565 8604
rect 10030 8490 10394 8536
rect 10440 8490 10508 8536
rect 10554 8490 10565 8536
rect 10030 8422 10565 8490
rect 10030 8376 10394 8422
rect 10440 8376 10508 8422
rect 10554 8376 10565 8422
rect 10030 8308 10565 8376
rect 10030 8262 10394 8308
rect 10440 8262 10508 8308
rect 10554 8262 10565 8308
rect 10030 8194 10565 8262
rect 10030 8148 10394 8194
rect 10440 8148 10508 8194
rect 10554 8148 10565 8194
rect 10030 8080 10565 8148
rect 10030 8034 10394 8080
rect 10440 8034 10508 8080
rect 10554 8034 10565 8080
rect 10030 7966 10565 8034
rect 10030 7920 10394 7966
rect 10440 7920 10508 7966
rect 10554 7920 10565 7966
rect 10030 7852 10565 7920
rect 10030 7806 10394 7852
rect 10440 7806 10508 7852
rect 10554 7806 10565 7852
rect 10030 7738 10565 7806
rect 10030 7692 10394 7738
rect 10440 7692 10508 7738
rect 10554 7692 10565 7738
rect 10030 7624 10565 7692
rect 10030 7578 10394 7624
rect 10440 7578 10508 7624
rect 10554 7578 10565 7624
rect 10030 7510 10565 7578
rect 10030 7464 10394 7510
rect 10440 7464 10508 7510
rect 10554 7464 10565 7510
rect 10030 7396 10565 7464
rect 10030 7350 10394 7396
rect 10440 7350 10508 7396
rect 10554 7350 10565 7396
rect 10030 7282 10565 7350
rect 10030 7236 10394 7282
rect 10440 7236 10508 7282
rect 10554 7236 10565 7282
rect 10030 7168 10565 7236
rect 10030 7122 10394 7168
rect 10440 7122 10508 7168
rect 10554 7122 10565 7168
rect 10030 7054 10565 7122
rect 10030 7008 10394 7054
rect 10440 7008 10508 7054
rect 10554 7008 10565 7054
rect 10030 6940 10565 7008
rect 10030 6894 10394 6940
rect 10440 6894 10508 6940
rect 10554 6894 10565 6940
rect 10030 6826 10565 6894
rect 10030 6780 10394 6826
rect 10440 6780 10508 6826
rect 10554 6780 10565 6826
rect 10030 6712 10565 6780
rect 10030 6670 10394 6712
rect 9973 6666 10394 6670
rect 10440 6666 10508 6712
rect 10554 6666 10565 6712
rect 7997 6600 9913 6611
rect 7997 6554 8008 6600
rect 9902 6554 9913 6600
rect 7997 6543 9913 6554
rect 9973 6598 10565 6666
rect 9973 6552 10394 6598
rect 10440 6552 10508 6598
rect 10554 6552 10565 6598
rect 9973 6484 10565 6552
rect 9973 6483 10394 6484
rect 5086 6438 10394 6483
rect 10440 6438 10508 6484
rect 10554 6438 10565 6484
rect 4915 6370 10565 6438
rect 4915 6324 4926 6370
rect 4972 6324 5040 6370
rect 5086 6324 10394 6370
rect 10440 6324 10508 6370
rect 10554 6324 10565 6370
rect 4915 6256 10565 6324
rect 4915 6210 4926 6256
rect 4972 6210 5040 6256
rect 5086 6210 10394 6256
rect 10440 6210 10508 6256
rect 10554 6210 10565 6256
rect 4915 6207 10565 6210
rect 4915 6161 5214 6207
rect 5260 6161 5328 6207
rect 5374 6161 5442 6207
rect 5488 6161 5556 6207
rect 5602 6161 5670 6207
rect 5716 6161 5784 6207
rect 5830 6161 5898 6207
rect 5944 6161 6012 6207
rect 6058 6161 6126 6207
rect 6172 6161 6240 6207
rect 6286 6161 6354 6207
rect 6400 6161 6468 6207
rect 6514 6161 6582 6207
rect 6628 6161 6696 6207
rect 6742 6161 6810 6207
rect 6856 6161 6924 6207
rect 6970 6161 7038 6207
rect 7084 6161 7152 6207
rect 7198 6161 7266 6207
rect 7312 6161 7380 6207
rect 7426 6161 7494 6207
rect 7540 6161 7608 6207
rect 7654 6161 7722 6207
rect 7768 6161 7836 6207
rect 7882 6161 7950 6207
rect 7996 6161 8064 6207
rect 8110 6161 8178 6207
rect 8224 6161 8292 6207
rect 8338 6161 8406 6207
rect 8452 6161 8520 6207
rect 8566 6161 8634 6207
rect 8680 6161 8748 6207
rect 8794 6161 8862 6207
rect 8908 6161 8976 6207
rect 9022 6161 9090 6207
rect 9136 6161 9204 6207
rect 9250 6161 9318 6207
rect 9364 6161 9432 6207
rect 9478 6161 9546 6207
rect 9592 6161 9660 6207
rect 9706 6161 9774 6207
rect 9820 6161 9888 6207
rect 9934 6161 10002 6207
rect 10048 6161 10116 6207
rect 10162 6161 10230 6207
rect 10276 6161 10565 6207
rect 4915 6142 10565 6161
rect 4915 6096 4926 6142
rect 4972 6096 5040 6142
rect 5086 6096 10394 6142
rect 10440 6096 10508 6142
rect 10554 6096 10565 6142
rect 4915 6093 10565 6096
rect 4915 6047 5214 6093
rect 5260 6047 5328 6093
rect 5374 6047 5442 6093
rect 5488 6047 5556 6093
rect 5602 6047 5670 6093
rect 5716 6047 5784 6093
rect 5830 6047 5898 6093
rect 5944 6047 6012 6093
rect 6058 6047 6126 6093
rect 6172 6047 6240 6093
rect 6286 6047 6354 6093
rect 6400 6047 6468 6093
rect 6514 6047 6582 6093
rect 6628 6047 6696 6093
rect 6742 6047 6810 6093
rect 6856 6047 6924 6093
rect 6970 6047 7038 6093
rect 7084 6047 7152 6093
rect 7198 6047 7266 6093
rect 7312 6047 7380 6093
rect 7426 6047 7494 6093
rect 7540 6047 7608 6093
rect 7654 6047 7722 6093
rect 7768 6047 7836 6093
rect 7882 6047 7950 6093
rect 7996 6047 8064 6093
rect 8110 6047 8178 6093
rect 8224 6047 8292 6093
rect 8338 6047 8406 6093
rect 8452 6047 8520 6093
rect 8566 6047 8634 6093
rect 8680 6047 8748 6093
rect 8794 6047 8862 6093
rect 8908 6047 8976 6093
rect 9022 6047 9090 6093
rect 9136 6047 9204 6093
rect 9250 6047 9318 6093
rect 9364 6047 9432 6093
rect 9478 6047 9546 6093
rect 9592 6047 9660 6093
rect 9706 6047 9774 6093
rect 9820 6047 9888 6093
rect 9934 6047 10002 6093
rect 10048 6047 10116 6093
rect 10162 6047 10230 6093
rect 10276 6047 10565 6093
rect 4915 6028 10565 6047
rect 4915 5982 4926 6028
rect 4972 5982 5040 6028
rect 5086 5982 10394 6028
rect 10440 5982 10508 6028
rect 10554 5982 10565 6028
rect 4915 5914 10565 5982
rect 4915 5868 4926 5914
rect 4972 5868 5040 5914
rect 5086 5868 10394 5914
rect 10440 5868 10508 5914
rect 10554 5868 10565 5914
rect 4915 5800 10565 5868
rect 4915 5754 4926 5800
rect 4972 5754 5040 5800
rect 5086 5771 10394 5800
rect 5086 5754 5501 5771
rect 4915 5686 5501 5754
rect 4915 5640 4926 5686
rect 4972 5640 5040 5686
rect 5086 5640 5501 5686
rect 5561 5700 7477 5711
rect 5561 5654 5572 5700
rect 7466 5654 7477 5700
rect 5561 5643 7477 5654
rect 4915 5584 5501 5640
rect 4915 5572 5444 5584
rect 4915 5526 4926 5572
rect 4972 5526 5040 5572
rect 5086 5526 5444 5572
rect 4915 5458 5444 5526
rect 4915 5412 4926 5458
rect 4972 5412 5040 5458
rect 5086 5412 5444 5458
rect 4915 5344 5444 5412
rect 4915 5298 4926 5344
rect 4972 5298 5040 5344
rect 5086 5298 5444 5344
rect 4915 5230 5444 5298
rect 4915 5184 4926 5230
rect 4972 5184 5040 5230
rect 5086 5184 5444 5230
rect 4915 5116 5444 5184
rect 4915 5070 4926 5116
rect 4972 5070 5040 5116
rect 5086 5070 5444 5116
rect 4915 5002 5444 5070
rect 4915 4956 4926 5002
rect 4972 4956 5040 5002
rect 5086 4956 5444 5002
rect 4915 4888 5444 4956
rect 4915 4842 4926 4888
rect 4972 4842 5040 4888
rect 5086 4842 5444 4888
rect 4915 4774 5444 4842
rect 4915 4728 4926 4774
rect 4972 4728 5040 4774
rect 5086 4728 5444 4774
rect 4915 4660 5444 4728
rect 4915 4614 4926 4660
rect 4972 4614 5040 4660
rect 5086 4614 5444 4660
rect 4915 4546 5444 4614
rect 4915 4500 4926 4546
rect 4972 4500 5040 4546
rect 5086 4500 5444 4546
rect 4915 4432 5444 4500
rect 4915 4386 4926 4432
rect 4972 4386 5040 4432
rect 5086 4386 5444 4432
rect 4915 4318 5444 4386
rect 4915 4272 4926 4318
rect 4972 4272 5040 4318
rect 5086 4272 5444 4318
rect 4915 4204 5444 4272
rect 4915 4158 4926 4204
rect 4972 4158 5040 4204
rect 5086 4158 5444 4204
rect 4915 4090 5444 4158
rect 4915 4044 4926 4090
rect 4972 4044 5040 4090
rect 5086 4044 5444 4090
rect 4915 3976 5444 4044
rect 4915 3930 4926 3976
rect 4972 3930 5040 3976
rect 5086 3930 5444 3976
rect 4915 3862 5444 3930
rect 4915 3816 4926 3862
rect 4972 3816 5040 3862
rect 5086 3816 5444 3862
rect 4915 3748 5444 3816
rect 4915 3702 4926 3748
rect 4972 3702 5040 3748
rect 5086 3702 5444 3748
rect 4915 3634 5444 3702
rect 4915 3588 4926 3634
rect 4972 3588 5040 3634
rect 5086 3588 5444 3634
rect 4915 3520 5444 3588
rect 4915 3474 4926 3520
rect 4972 3474 5040 3520
rect 5086 3474 5444 3520
rect 4915 3406 5444 3474
rect 4915 3360 4926 3406
rect 4972 3360 5040 3406
rect 5086 3360 5444 3406
rect 4915 3292 5444 3360
rect 4915 3246 4926 3292
rect 4972 3246 5040 3292
rect 5086 3246 5444 3292
rect 4915 3178 5444 3246
rect 4915 3132 4926 3178
rect 4972 3132 5040 3178
rect 5086 3132 5444 3178
rect 4915 3064 5444 3132
rect 4915 3018 4926 3064
rect 4972 3018 5040 3064
rect 5086 3018 5444 3064
rect 4915 2950 5444 3018
rect 4915 2904 4926 2950
rect 4972 2904 5040 2950
rect 5086 2904 5444 2950
rect 4915 2836 5444 2904
rect 4915 2790 4926 2836
rect 4972 2790 5040 2836
rect 5086 2790 5444 2836
rect 4915 2722 5444 2790
rect 4915 2676 4926 2722
rect 4972 2676 5040 2722
rect 5086 2676 5444 2722
rect 4915 2608 5444 2676
rect 4915 2562 4926 2608
rect 4972 2562 5040 2608
rect 5086 2562 5444 2608
rect 4915 2494 5444 2562
rect 4915 2448 4926 2494
rect 4972 2448 5040 2494
rect 5086 2448 5444 2494
rect 4915 2380 5444 2448
rect 4915 2334 4926 2380
rect 4972 2334 5040 2380
rect 5086 2334 5444 2380
rect 4915 2266 5444 2334
rect 4915 2220 4926 2266
rect 4972 2220 5040 2266
rect 5086 2220 5444 2266
rect 4915 2152 5444 2220
rect 4915 2106 4926 2152
rect 4972 2106 5040 2152
rect 5086 2106 5444 2152
rect 4915 2038 5444 2106
rect 4915 1992 4926 2038
rect 4972 1992 5040 2038
rect 5086 1992 5444 2038
rect 4915 1924 5444 1992
rect 4915 1878 4926 1924
rect 4972 1878 5040 1924
rect 5086 1878 5444 1924
rect 4915 1810 5444 1878
rect 4915 1764 4926 1810
rect 4972 1764 5040 1810
rect 5086 1764 5444 1810
rect 4915 1696 5444 1764
rect 4915 1650 4926 1696
rect 4972 1650 5040 1696
rect 5086 1650 5444 1696
rect 4915 1582 5444 1650
rect 4915 1536 4926 1582
rect 4972 1536 5040 1582
rect 5086 1536 5444 1582
rect 4915 1468 5444 1536
rect 4915 1422 4926 1468
rect 4972 1422 5040 1468
rect 5086 1422 5444 1468
rect 4915 1354 5444 1422
rect 4915 1308 4926 1354
rect 4972 1308 5040 1354
rect 5086 1308 5444 1354
rect 4915 1240 5444 1308
rect 4915 1194 4926 1240
rect 4972 1194 5040 1240
rect 5086 1194 5444 1240
rect 4915 1126 5444 1194
rect 4915 1080 4926 1126
rect 4972 1080 5040 1126
rect 5086 1080 5444 1126
rect 4915 1012 5444 1080
rect 4915 966 4926 1012
rect 4972 966 5040 1012
rect 5086 966 5444 1012
rect 4915 898 5444 966
rect 4915 852 4926 898
rect 4972 852 5040 898
rect 5086 852 5444 898
rect 4915 784 5444 852
rect 4915 738 4926 784
rect 4972 738 5040 784
rect 5086 738 5444 784
rect 4915 658 5444 738
rect 5490 658 5501 5584
rect 4915 621 5501 658
rect 4915 328 5097 621
rect 6019 599 7019 5643
rect 7537 5584 7937 5771
rect 9973 5754 10394 5771
rect 10440 5754 10508 5800
rect 10554 5754 10565 5800
rect 7997 5700 9913 5711
rect 7997 5654 8008 5700
rect 9902 5654 9913 5700
rect 7997 5643 9913 5654
rect 9973 5686 10565 5754
rect 7537 658 7548 5584
rect 7594 658 7880 5584
rect 7926 658 7937 5584
rect 7537 621 7937 658
rect 8455 599 9455 5643
rect 9973 5640 10394 5686
rect 10440 5640 10508 5686
rect 10554 5640 10565 5686
rect 9973 5584 10565 5640
rect 9973 658 9984 5584
rect 10030 5572 10565 5584
rect 10030 5526 10394 5572
rect 10440 5526 10508 5572
rect 10554 5526 10565 5572
rect 10030 5458 10565 5526
rect 10030 5412 10394 5458
rect 10440 5412 10508 5458
rect 10554 5412 10565 5458
rect 10030 5344 10565 5412
rect 10030 5298 10394 5344
rect 10440 5298 10508 5344
rect 10554 5298 10565 5344
rect 10030 5230 10565 5298
rect 10030 5184 10394 5230
rect 10440 5184 10508 5230
rect 10554 5184 10565 5230
rect 10030 5116 10565 5184
rect 10030 5070 10394 5116
rect 10440 5070 10508 5116
rect 10554 5070 10565 5116
rect 10030 5002 10565 5070
rect 10030 4956 10394 5002
rect 10440 4956 10508 5002
rect 10554 4956 10565 5002
rect 10030 4888 10565 4956
rect 10030 4842 10394 4888
rect 10440 4842 10508 4888
rect 10554 4842 10565 4888
rect 10030 4774 10565 4842
rect 10030 4728 10394 4774
rect 10440 4728 10508 4774
rect 10554 4728 10565 4774
rect 10030 4660 10565 4728
rect 10030 4614 10394 4660
rect 10440 4614 10508 4660
rect 10554 4614 10565 4660
rect 10030 4546 10565 4614
rect 10030 4500 10394 4546
rect 10440 4500 10508 4546
rect 10554 4500 10565 4546
rect 10030 4432 10565 4500
rect 10030 4386 10394 4432
rect 10440 4386 10508 4432
rect 10554 4386 10565 4432
rect 10030 4318 10565 4386
rect 10030 4272 10394 4318
rect 10440 4272 10508 4318
rect 10554 4272 10565 4318
rect 10030 4204 10565 4272
rect 10030 4158 10394 4204
rect 10440 4158 10508 4204
rect 10554 4158 10565 4204
rect 10030 4090 10565 4158
rect 10030 4044 10394 4090
rect 10440 4044 10508 4090
rect 10554 4044 10565 4090
rect 10030 3976 10565 4044
rect 10030 3930 10394 3976
rect 10440 3930 10508 3976
rect 10554 3930 10565 3976
rect 10030 3862 10565 3930
rect 10030 3816 10394 3862
rect 10440 3816 10508 3862
rect 10554 3816 10565 3862
rect 10030 3748 10565 3816
rect 10030 3702 10394 3748
rect 10440 3702 10508 3748
rect 10554 3702 10565 3748
rect 10030 3634 10565 3702
rect 10030 3588 10394 3634
rect 10440 3588 10508 3634
rect 10554 3588 10565 3634
rect 10030 3520 10565 3588
rect 10030 3474 10394 3520
rect 10440 3474 10508 3520
rect 10554 3474 10565 3520
rect 10030 3406 10565 3474
rect 10030 3360 10394 3406
rect 10440 3360 10508 3406
rect 10554 3360 10565 3406
rect 10030 3292 10565 3360
rect 10030 3246 10394 3292
rect 10440 3246 10508 3292
rect 10554 3246 10565 3292
rect 10030 3178 10565 3246
rect 10030 3132 10394 3178
rect 10440 3132 10508 3178
rect 10554 3132 10565 3178
rect 10030 3064 10565 3132
rect 10030 3018 10394 3064
rect 10440 3018 10508 3064
rect 10554 3018 10565 3064
rect 10030 2950 10565 3018
rect 10030 2904 10394 2950
rect 10440 2904 10508 2950
rect 10554 2904 10565 2950
rect 10030 2836 10565 2904
rect 10030 2790 10394 2836
rect 10440 2790 10508 2836
rect 10554 2790 10565 2836
rect 10030 2722 10565 2790
rect 10030 2676 10394 2722
rect 10440 2676 10508 2722
rect 10554 2676 10565 2722
rect 10030 2608 10565 2676
rect 10030 2562 10394 2608
rect 10440 2562 10508 2608
rect 10554 2562 10565 2608
rect 10030 2494 10565 2562
rect 10030 2448 10394 2494
rect 10440 2448 10508 2494
rect 10554 2448 10565 2494
rect 10030 2380 10565 2448
rect 10030 2334 10394 2380
rect 10440 2334 10508 2380
rect 10554 2334 10565 2380
rect 10030 2266 10565 2334
rect 10030 2220 10394 2266
rect 10440 2220 10508 2266
rect 10554 2220 10565 2266
rect 10030 2152 10565 2220
rect 10030 2106 10394 2152
rect 10440 2106 10508 2152
rect 10554 2106 10565 2152
rect 10030 2038 10565 2106
rect 10030 1992 10394 2038
rect 10440 1992 10508 2038
rect 10554 1992 10565 2038
rect 10030 1924 10565 1992
rect 10030 1878 10394 1924
rect 10440 1878 10508 1924
rect 10554 1878 10565 1924
rect 10030 1810 10565 1878
rect 10030 1764 10394 1810
rect 10440 1764 10508 1810
rect 10554 1764 10565 1810
rect 10030 1696 10565 1764
rect 10030 1650 10394 1696
rect 10440 1650 10508 1696
rect 10554 1650 10565 1696
rect 10030 1582 10565 1650
rect 10030 1536 10394 1582
rect 10440 1536 10508 1582
rect 10554 1536 10565 1582
rect 10030 1468 10565 1536
rect 10030 1422 10394 1468
rect 10440 1422 10508 1468
rect 10554 1422 10565 1468
rect 10030 1354 10565 1422
rect 10030 1308 10394 1354
rect 10440 1308 10508 1354
rect 10554 1308 10565 1354
rect 10030 1240 10565 1308
rect 10030 1194 10394 1240
rect 10440 1194 10508 1240
rect 10554 1194 10565 1240
rect 10030 1126 10565 1194
rect 10030 1080 10394 1126
rect 10440 1080 10508 1126
rect 10554 1080 10565 1126
rect 10030 1012 10565 1080
rect 10030 966 10394 1012
rect 10440 966 10508 1012
rect 10554 966 10565 1012
rect 10030 898 10565 966
rect 10030 852 10394 898
rect 10440 852 10508 898
rect 10554 852 10565 898
rect 10030 784 10565 852
rect 10030 738 10394 784
rect 10440 738 10508 784
rect 10554 738 10565 784
rect 10030 670 10565 738
rect 10030 658 10394 670
rect 9973 624 10394 658
rect 10440 624 10508 670
rect 10554 624 10565 670
rect 9973 621 10565 624
rect 5561 588 7477 599
rect 5561 542 5572 588
rect 7466 542 7477 588
rect 5561 531 7477 542
rect 7997 588 9913 599
rect 7997 542 8008 588
rect 9902 542 9913 588
rect 7997 531 9913 542
rect 5561 399 9913 531
rect 10383 556 10565 621
rect 10383 510 10394 556
rect 10440 510 10508 556
rect 10554 510 10565 556
rect 10383 442 10565 510
rect 4915 282 4926 328
rect 4972 282 5040 328
rect 5086 282 5097 328
rect 4915 226 5097 282
rect 10383 396 10394 442
rect 10440 396 10508 442
rect 10554 396 10565 442
rect 10383 328 10565 396
rect 10383 282 10394 328
rect 10440 282 10508 328
rect 10554 282 10565 328
rect 10383 226 10565 282
rect 4915 214 10565 226
rect 4915 168 4926 214
rect 4972 168 5040 214
rect 5086 168 5222 214
rect 5268 168 5336 214
rect 5382 168 5450 214
rect 5496 168 5564 214
rect 5610 168 5678 214
rect 5724 168 5792 214
rect 5838 168 5906 214
rect 5952 168 6020 214
rect 6066 168 6134 214
rect 6180 168 6248 214
rect 6294 168 6362 214
rect 6408 168 6476 214
rect 6522 168 6590 214
rect 6636 168 6704 214
rect 6750 168 6818 214
rect 6864 168 6932 214
rect 6978 168 7046 214
rect 7092 168 7160 214
rect 7206 168 7274 214
rect 7320 168 7388 214
rect 7434 168 7502 214
rect 7548 168 7616 214
rect 7662 168 7730 214
rect 7776 168 7844 214
rect 7890 168 7958 214
rect 8004 168 8072 214
rect 8118 168 8186 214
rect 8232 168 8300 214
rect 8346 168 8414 214
rect 8460 168 8528 214
rect 8574 168 8642 214
rect 8688 168 8756 214
rect 8802 168 8870 214
rect 8916 168 8984 214
rect 9030 168 9098 214
rect 9144 168 9212 214
rect 9258 168 9326 214
rect 9372 168 9440 214
rect 9486 168 9554 214
rect 9600 168 9668 214
rect 9714 168 9782 214
rect 9828 168 9896 214
rect 9942 168 10010 214
rect 10056 168 10124 214
rect 10170 168 10238 214
rect 10284 168 10394 214
rect 10440 168 10508 214
rect 10554 168 10565 214
rect 4915 100 10565 168
rect 4915 54 4926 100
rect 4972 54 5040 100
rect 5086 54 5222 100
rect 5268 54 5336 100
rect 5382 54 5450 100
rect 5496 54 5564 100
rect 5610 54 5678 100
rect 5724 54 5792 100
rect 5838 54 5906 100
rect 5952 54 6020 100
rect 6066 54 6134 100
rect 6180 54 6248 100
rect 6294 54 6362 100
rect 6408 54 6476 100
rect 6522 54 6590 100
rect 6636 54 6704 100
rect 6750 54 6818 100
rect 6864 54 6932 100
rect 6978 54 7046 100
rect 7092 54 7160 100
rect 7206 54 7274 100
rect 7320 54 7388 100
rect 7434 54 7502 100
rect 7548 54 7616 100
rect 7662 54 7730 100
rect 7776 54 7844 100
rect 7890 54 7958 100
rect 8004 54 8072 100
rect 8118 54 8186 100
rect 8232 54 8300 100
rect 8346 54 8414 100
rect 8460 54 8528 100
rect 8574 54 8642 100
rect 8688 54 8756 100
rect 8802 54 8870 100
rect 8916 54 8984 100
rect 9030 54 9098 100
rect 9144 54 9212 100
rect 9258 54 9326 100
rect 9372 54 9440 100
rect 9486 54 9554 100
rect 9600 54 9668 100
rect 9714 54 9782 100
rect 9828 54 9896 100
rect 9942 54 10010 100
rect 10056 54 10124 100
rect 10170 54 10238 100
rect 10284 54 10394 100
rect 10440 54 10508 100
rect 10554 54 10565 100
rect 4915 42 10565 54
use M1_PSUB_CDNS_40661954729136  M1_PSUB_CDNS_40661954729136_0
timestamp 1698431365
transform 1 0 10474 0 1 6176
box 0 0 1 1
use M1_PSUB_CDNS_40661954729137  M1_PSUB_CDNS_40661954729137_0
timestamp 1698431365
transform 0 -1 7748 1 0 12218
box 0 0 1 1
use M1_PSUB_CDNS_40661954729137  M1_PSUB_CDNS_40661954729137_1
timestamp 1698431365
transform 0 -1 7745 1 0 6127
box 0 0 1 1
use M1_PSUB_CDNS_40661954729137  M1_PSUB_CDNS_40661954729137_2
timestamp 1698431365
transform 0 -1 7753 1 0 134
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_0
timestamp 1698431365
transform 1 0 7955 0 -1 5621
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_1
timestamp 1698431365
transform 1 0 5519 0 -1 5621
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_2
timestamp 1698431365
transform 1 0 7955 0 1 6633
box 0 0 1 1
use nmoscap_6p0_CDNS_406619547290  nmoscap_6p0_CDNS_406619547290_3
timestamp 1698431365
transform 1 0 5519 0 1 6633
box 0 0 1 1
<< properties >>
string GDS_END 4793568
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4778802
<< end >>
