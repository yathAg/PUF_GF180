magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 2102 870
rect -86 352 215 377
rect 923 352 2102 377
<< pwell >>
rect -86 -86 2102 352
<< mvnmos >>
rect 124 68 244 232
rect 392 93 512 257
rect 616 93 736 257
rect 884 68 1004 232
rect 1109 68 1229 232
rect 1313 68 1433 232
rect 1537 68 1657 232
rect 1721 68 1841 232
<< mvpmos >>
rect 144 497 244 716
rect 412 497 512 716
rect 616 497 716 716
rect 884 497 984 716
rect 1129 519 1229 716
rect 1333 519 1433 716
rect 1537 519 1637 716
rect 1741 519 1841 716
<< mvndiff >>
rect 304 244 392 257
rect 304 232 317 244
rect 36 152 124 232
rect 36 106 49 152
rect 95 106 124 152
rect 36 68 124 106
rect 244 198 317 232
rect 363 198 392 244
rect 244 93 392 198
rect 512 152 616 257
rect 512 106 541 152
rect 587 106 616 152
rect 512 93 616 106
rect 736 244 824 257
rect 736 198 765 244
rect 811 232 824 244
rect 811 198 884 232
rect 736 93 884 198
rect 244 68 332 93
rect 804 68 884 93
rect 1004 152 1109 232
rect 1004 106 1034 152
rect 1080 106 1109 152
rect 1004 68 1109 106
rect 1229 68 1313 232
rect 1433 127 1537 232
rect 1433 81 1462 127
rect 1508 81 1537 127
rect 1433 68 1537 81
rect 1657 68 1721 232
rect 1841 152 1929 232
rect 1841 106 1870 152
rect 1916 106 1929 152
rect 1841 68 1929 106
<< mvpdiff >>
rect 56 678 144 716
rect 56 538 69 678
rect 115 538 144 678
rect 56 497 144 538
rect 244 497 412 716
rect 512 644 616 716
rect 512 598 541 644
rect 587 598 616 644
rect 512 497 616 598
rect 716 497 884 716
rect 984 687 1129 716
rect 984 641 1034 687
rect 1080 641 1129 687
rect 984 519 1129 641
rect 1229 644 1333 716
rect 1229 598 1258 644
rect 1304 598 1333 644
rect 1229 519 1333 598
rect 1433 687 1537 716
rect 1433 641 1462 687
rect 1508 641 1537 687
rect 1433 519 1537 641
rect 1637 644 1741 716
rect 1637 598 1666 644
rect 1712 598 1741 644
rect 1637 519 1741 598
rect 1841 678 1929 716
rect 1841 538 1870 678
rect 1916 538 1929 678
rect 1841 519 1929 538
rect 984 497 1064 519
<< mvndiffc >>
rect 49 106 95 152
rect 317 198 363 244
rect 541 106 587 152
rect 765 198 811 244
rect 1034 106 1080 152
rect 1462 81 1508 127
rect 1870 106 1916 152
<< mvpdiffc >>
rect 69 538 115 678
rect 541 598 587 644
rect 1034 641 1080 687
rect 1258 598 1304 644
rect 1462 641 1508 687
rect 1666 598 1712 644
rect 1870 538 1916 678
<< polysilicon >>
rect 144 716 244 760
rect 412 716 512 760
rect 616 716 716 760
rect 884 716 984 760
rect 1129 716 1229 760
rect 1333 716 1433 760
rect 1537 716 1637 760
rect 1741 716 1841 760
rect 144 401 244 497
rect 412 415 512 497
rect 412 401 439 415
rect 124 367 244 401
rect 124 321 174 367
rect 220 321 244 367
rect 124 232 244 321
rect 392 369 439 401
rect 485 401 512 415
rect 616 415 716 497
rect 616 401 643 415
rect 485 369 643 401
rect 689 401 716 415
rect 884 415 984 497
rect 689 369 736 401
rect 392 348 736 369
rect 392 257 512 348
rect 616 257 736 348
rect 884 369 915 415
rect 961 401 984 415
rect 1129 401 1229 519
rect 1333 415 1433 519
rect 1333 401 1360 415
rect 961 369 1004 401
rect 884 232 1004 369
rect 1109 394 1229 401
rect 1109 348 1153 394
rect 1199 348 1229 394
rect 1109 232 1229 348
rect 1313 369 1360 401
rect 1406 401 1433 415
rect 1537 415 1637 519
rect 1537 401 1564 415
rect 1406 369 1564 401
rect 1610 401 1637 415
rect 1741 401 1841 519
rect 1610 369 1657 401
rect 1313 348 1657 369
rect 1313 232 1433 348
rect 1537 232 1657 348
rect 1721 394 1841 401
rect 1721 348 1776 394
rect 1822 348 1841 394
rect 1721 232 1841 348
rect 124 24 244 68
rect 392 24 512 93
rect 616 24 736 93
rect 884 24 1004 68
rect 1109 24 1229 68
rect 1313 24 1433 68
rect 1537 24 1657 68
rect 1721 24 1841 68
<< polycontact >>
rect 174 321 220 367
rect 439 369 485 415
rect 643 369 689 415
rect 915 369 961 415
rect 1153 348 1199 394
rect 1360 369 1406 415
rect 1564 369 1610 415
rect 1776 348 1822 394
<< metal1 >>
rect 0 724 2016 844
rect 69 678 115 724
rect 1023 687 1091 724
rect 426 644 972 656
rect 426 598 541 644
rect 587 598 972 644
rect 1023 641 1034 687
rect 1080 641 1091 687
rect 1451 687 1519 724
rect 1258 644 1304 655
rect 426 584 972 598
rect 69 497 115 538
rect 926 536 972 584
rect 1451 641 1462 687
rect 1508 641 1519 687
rect 1870 678 1916 724
rect 1666 644 1712 655
rect 1258 536 1304 598
rect 1666 536 1712 598
rect 165 470 876 536
rect 926 476 1712 536
rect 1870 519 1916 538
rect 926 474 1096 476
rect 165 367 229 470
rect 824 424 876 470
rect 165 321 174 367
rect 220 321 229 367
rect 312 415 774 424
rect 312 369 439 415
rect 485 369 643 415
rect 689 369 774 415
rect 312 358 774 369
rect 824 415 980 424
rect 824 369 915 415
rect 961 369 980 415
rect 824 358 980 369
rect 165 232 229 321
rect 1030 312 1096 474
rect 306 244 1096 312
rect 1144 394 1208 430
rect 1144 348 1153 394
rect 1199 348 1208 394
rect 1256 415 1664 428
rect 1256 369 1360 415
rect 1406 369 1564 415
rect 1610 369 1664 415
rect 1256 360 1664 369
rect 1773 394 1884 438
rect 1144 311 1208 348
rect 1773 348 1776 394
rect 1822 348 1884 394
rect 1773 311 1884 348
rect 1144 265 1884 311
rect 306 198 317 244
rect 363 198 374 244
rect 754 198 765 244
rect 811 198 822 244
rect 1144 238 1297 265
rect 1676 238 1884 265
rect 1347 173 1616 219
rect 1347 152 1393 173
rect 36 106 49 152
rect 95 106 541 152
rect 587 106 1034 152
rect 1080 106 1393 152
rect 1570 152 1616 173
rect 1451 81 1462 127
rect 1508 81 1519 127
rect 1570 106 1870 152
rect 1916 106 1929 152
rect 1451 60 1519 81
rect 0 -60 2016 60
<< labels >>
flabel metal1 s 165 470 876 536 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel metal1 s 426 655 972 656 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 312 358 774 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1773 430 1884 438 0 FreeSans 400 0 0 0 B
port 3 nsew default input
flabel metal1 s 1256 360 1664 428 0 FreeSans 400 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 724 2016 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1451 60 1519 127 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 824 424 876 470 1 A2
port 2 nsew default input
rlabel metal1 s 165 424 229 470 1 A2
port 2 nsew default input
rlabel metal1 s 824 358 980 424 1 A2
port 2 nsew default input
rlabel metal1 s 165 358 229 424 1 A2
port 2 nsew default input
rlabel metal1 s 165 232 229 358 1 A2
port 2 nsew default input
rlabel metal1 s 1773 311 1884 430 1 B
port 3 nsew default input
rlabel metal1 s 1144 311 1208 430 1 B
port 3 nsew default input
rlabel metal1 s 1144 265 1884 311 1 B
port 3 nsew default input
rlabel metal1 s 1676 238 1884 265 1 B
port 3 nsew default input
rlabel metal1 s 1144 238 1297 265 1 B
port 3 nsew default input
rlabel metal1 s 1666 584 1712 655 1 ZN
port 5 nsew default output
rlabel metal1 s 1258 584 1304 655 1 ZN
port 5 nsew default output
rlabel metal1 s 426 584 972 655 1 ZN
port 5 nsew default output
rlabel metal1 s 1666 536 1712 584 1 ZN
port 5 nsew default output
rlabel metal1 s 1258 536 1304 584 1 ZN
port 5 nsew default output
rlabel metal1 s 926 536 972 584 1 ZN
port 5 nsew default output
rlabel metal1 s 926 476 1712 536 1 ZN
port 5 nsew default output
rlabel metal1 s 926 474 1096 476 1 ZN
port 5 nsew default output
rlabel metal1 s 1030 312 1096 474 1 ZN
port 5 nsew default output
rlabel metal1 s 306 244 1096 312 1 ZN
port 5 nsew default output
rlabel metal1 s 754 198 822 244 1 ZN
port 5 nsew default output
rlabel metal1 s 306 198 374 244 1 ZN
port 5 nsew default output
rlabel metal1 s 1870 641 1916 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1451 641 1519 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1023 641 1091 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 641 115 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1870 519 1916 641 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 519 115 641 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 497 115 519 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -60 2016 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 784
string GDS_END 97542
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 92760
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
