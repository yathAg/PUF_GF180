magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
use M1_NACTIVE4310591302024_512x8m81  M1_NACTIVE4310591302024_512x8m81_0
timestamp 1698431365
transform 1 0 1337 0 1 4210
box 0 0 1 1
use M1_POLY24310591302059_512x8m81  M1_POLY24310591302059_512x8m81_0
timestamp 1698431365
transform 1 0 865 0 1 7450
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1698431365
transform -1 0 824 0 1 4092
box 0 0 1 1
use M2_M1$$43376684_512x8m81  M2_M1$$43376684_512x8m81_0
timestamp 1698431365
transform -1 0 599 0 1 2099
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_0
timestamp 1698431365
transform 1 0 1113 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_1
timestamp 1698431365
transform 1 0 881 0 1 10532
box 0 0 1 1
use M2_M1$$43379756_512x8m81  M2_M1$$43379756_512x8m81_2
timestamp 1698431365
transform 1 0 441 0 1 10532
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_0
timestamp 1698431365
transform 1 0 441 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_1
timestamp 1698431365
transform 1 0 889 0 1 9494
box 0 0 1 1
use M2_M1$$43380780_512x8m81  M2_M1$$43380780_512x8m81_2
timestamp 1698431365
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_0
timestamp 1698431365
transform 1 0 1054 0 1 6153
box 0 0 1 1
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_1
timestamp 1698431365
transform 1 0 602 0 1 6153
box 0 0 1 1
use M2_M1$$47500332_512x8m81  M2_M1$$47500332_512x8m81_2
timestamp 1698431365
transform 1 0 1337 0 1 6153
box 0 0 1 1
use M2_M1$$47640620_512x8m81  M2_M1$$47640620_512x8m81_0
timestamp 1698431365
transform 1 0 1337 0 1 1526
box 0 0 1 1
use M2_M1$$47640620_512x8m81  M2_M1$$47640620_512x8m81_1
timestamp 1698431365
transform 1 0 1054 0 1 1526
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_0
timestamp 1698431365
transform 1 0 1337 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_1
timestamp 1698431365
transform 1 0 1054 0 1 2505
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_2
timestamp 1698431365
transform 1 0 441 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_3
timestamp 1698431365
transform 1 0 889 0 1 9494
box 0 0 1 1
use M3_M2$$47108140_512x8m81  M3_M2$$47108140_512x8m81_4
timestamp 1698431365
transform 1 0 1337 0 1 9494
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_0
timestamp 1698431365
transform 1 0 1337 0 1 438
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_1
timestamp 1698431365
transform 1 0 1054 0 1 438
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_2
timestamp 1698431365
transform 1 0 881 0 1 10532
box 0 0 1 1
use M3_M2$$47333420_512x8m81  M3_M2$$47333420_512x8m81_3
timestamp 1698431365
transform 1 0 441 0 1 10532
box 0 0 1 1
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_0
timestamp 1698431365
transform 1 0 1054 0 1 6153
box 0 0 1 1
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_1
timestamp 1698431365
transform 1 0 602 0 1 6153
box 0 0 1 1
use M3_M2$$47644716_512x8m81  M3_M2$$47644716_512x8m81_2
timestamp 1698431365
transform 1 0 1337 0 1 6153
box 0 0 1 1
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_0
timestamp 1698431365
transform -1 0 1254 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_1
timestamp 1698431365
transform -1 0 806 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_2
timestamp 1698431365
transform -1 0 582 0 -1 11038
box -31 0 -30 1
use nmos_1p2$$47641644_512x8m81  nmos_1p2$$47641644_512x8m81_3
timestamp 1698431365
transform -1 0 1030 0 -1 11038
box -31 0 -30 1
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_0
timestamp 1698431365
transform -1 0 1030 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_1
timestamp 1698431365
transform -1 0 806 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_2
timestamp 1698431365
transform -1 0 582 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47513644_512x8m81  pmos_1p2$$47513644_512x8m81_3
timestamp 1698431365
transform -1 0 1254 0 -1 9850
box -31 0 -30 1
use pmos_1p2$$47642668_512x8m81  pmos_1p2$$47642668_512x8m81_0
timestamp 1698431365
transform -1 0 964 0 1 3908
box -31 0 -30 1
use pmos_1p2$$47643692_512x8m81  pmos_1p2$$47643692_512x8m81_0
timestamp 1698431365
transform -1 0 740 0 1 3908
box -31 0 -30 1
<< properties >>
string GDS_END 560808
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 552470
<< end >>
