magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 3558 870
<< pwell >>
rect -86 -86 3558 352
<< mvnmos >>
rect 179 68 299 140
rect 403 68 523 140
rect 571 68 691 140
rect 1027 68 1147 140
rect 1195 68 1315 140
rect 1419 68 1539 140
rect 1587 68 1707 140
rect 2063 68 2183 141
rect 2231 68 2351 141
rect 2492 68 2612 232
rect 2755 68 2875 232
rect 2979 68 3099 232
rect 3203 68 3323 232
<< mvpmos >>
rect 179 644 279 716
rect 403 644 503 716
rect 571 644 671 716
rect 1007 644 1107 716
rect 1175 644 1275 716
rect 1459 644 1559 716
rect 1627 644 1727 716
rect 2063 622 2163 694
rect 2231 622 2331 694
rect 2561 472 2661 716
rect 2775 472 2875 716
rect 2979 472 3079 716
rect 3193 472 3293 716
<< mvndiff >>
rect 47 180 119 193
rect 47 134 60 180
rect 106 140 119 180
rect 751 200 823 213
rect 751 154 764 200
rect 810 154 823 200
rect 751 140 823 154
rect 106 134 179 140
rect 47 68 179 134
rect 299 127 403 140
rect 299 81 328 127
rect 374 81 403 127
rect 299 68 403 81
rect 523 68 571 140
rect 691 68 823 140
rect 895 200 967 213
rect 895 154 908 200
rect 954 154 967 200
rect 895 140 967 154
rect 1767 200 1839 213
rect 1767 154 1780 200
rect 1826 154 1839 200
rect 1767 140 1839 154
rect 895 68 1027 140
rect 1147 68 1195 140
rect 1315 127 1419 140
rect 1315 81 1344 127
rect 1390 81 1419 127
rect 1315 68 1419 81
rect 1539 68 1587 140
rect 1707 68 1839 140
rect 1931 200 2003 213
rect 1931 154 1944 200
rect 1990 154 2003 200
rect 1931 141 2003 154
rect 2412 141 2492 232
rect 1931 68 2063 141
rect 2183 68 2231 141
rect 2351 128 2492 141
rect 2351 82 2385 128
rect 2431 82 2492 128
rect 2351 68 2492 82
rect 2612 192 2755 232
rect 2612 146 2680 192
rect 2726 146 2755 192
rect 2612 68 2755 146
rect 2875 128 2979 232
rect 2875 82 2904 128
rect 2950 82 2979 128
rect 2875 68 2979 82
rect 3099 192 3203 232
rect 3099 146 3128 192
rect 3174 146 3203 192
rect 3099 68 3203 146
rect 3323 128 3411 232
rect 3323 82 3352 128
rect 3398 82 3411 128
rect 3323 68 3411 82
<< mvpdiff >>
rect 47 644 179 716
rect 279 703 403 716
rect 279 657 308 703
rect 354 657 403 703
rect 279 644 403 657
rect 503 644 571 716
rect 671 644 803 716
rect 47 621 119 644
rect 47 575 60 621
rect 106 575 119 621
rect 47 562 119 575
rect 731 621 803 644
rect 731 575 744 621
rect 790 575 803 621
rect 731 562 803 575
rect 875 644 1007 716
rect 1107 644 1175 716
rect 1275 703 1459 716
rect 1275 657 1304 703
rect 1350 657 1459 703
rect 1275 644 1459 657
rect 1559 644 1627 716
rect 1727 644 1859 716
rect 2481 694 2561 716
rect 875 621 947 644
rect 875 575 888 621
rect 934 575 947 621
rect 875 562 947 575
rect 1787 621 1859 644
rect 1787 575 1800 621
rect 1846 575 1859 621
rect 1787 562 1859 575
rect 1931 622 2063 694
rect 2163 622 2231 694
rect 2331 681 2561 694
rect 2331 635 2360 681
rect 2406 635 2561 681
rect 2331 622 2561 635
rect 1931 621 2003 622
rect 1931 575 1944 621
rect 1990 575 2003 621
rect 1931 562 2003 575
rect 2481 472 2561 622
rect 2661 639 2775 716
rect 2661 593 2690 639
rect 2736 593 2775 639
rect 2661 531 2775 593
rect 2661 485 2690 531
rect 2736 485 2775 531
rect 2661 472 2775 485
rect 2875 681 2979 716
rect 2875 635 2904 681
rect 2950 635 2979 681
rect 2875 472 2979 635
rect 3079 639 3193 716
rect 3079 593 3108 639
rect 3154 593 3193 639
rect 3079 531 3193 593
rect 3079 485 3108 531
rect 3154 485 3193 531
rect 3079 472 3193 485
rect 3293 681 3381 716
rect 3293 541 3322 681
rect 3368 541 3381 681
rect 3293 472 3381 541
<< mvndiffc >>
rect 60 134 106 180
rect 764 154 810 200
rect 328 81 374 127
rect 908 154 954 200
rect 1780 154 1826 200
rect 1344 81 1390 127
rect 1944 154 1990 200
rect 2385 82 2431 128
rect 2680 146 2726 192
rect 2904 82 2950 128
rect 3128 146 3174 192
rect 3352 82 3398 128
<< mvpdiffc >>
rect 308 657 354 703
rect 60 575 106 621
rect 744 575 790 621
rect 1304 657 1350 703
rect 888 575 934 621
rect 1800 575 1846 621
rect 2360 635 2406 681
rect 1944 575 1990 621
rect 2690 593 2736 639
rect 2690 485 2736 531
rect 2904 635 2950 681
rect 3108 593 3154 639
rect 3108 485 3154 531
rect 3322 541 3368 681
<< polysilicon >>
rect 179 716 279 760
rect 403 716 503 760
rect 571 716 671 760
rect 1007 716 1107 760
rect 1175 716 1275 760
rect 1459 716 1559 760
rect 1627 716 1727 760
rect 179 303 279 644
rect 179 257 192 303
rect 238 257 279 303
rect 179 184 279 257
rect 403 483 503 644
rect 571 483 671 644
rect 2063 694 2163 738
rect 2231 694 2331 738
rect 2561 716 2661 760
rect 2775 716 2875 760
rect 2979 716 3079 760
rect 3193 716 3293 760
rect 403 470 671 483
rect 403 424 416 470
rect 462 424 596 470
rect 642 424 671 470
rect 403 411 671 424
rect 403 184 503 411
rect 571 184 671 411
rect 1007 371 1107 644
rect 1175 371 1275 644
rect 1007 350 1275 371
rect 1007 304 1020 350
rect 1160 304 1275 350
rect 1007 290 1275 304
rect 179 140 299 184
rect 403 140 523 184
rect 571 140 691 184
rect 1027 140 1147 290
rect 1195 184 1275 290
rect 1459 371 1559 644
rect 1627 371 1727 644
rect 1459 350 1727 371
rect 1459 304 1472 350
rect 1612 304 1727 350
rect 1459 290 1727 304
rect 2063 377 2163 622
rect 2231 377 2331 622
rect 2063 364 2331 377
rect 2561 365 2661 472
rect 2775 365 2875 472
rect 2979 365 3079 472
rect 3193 365 3293 472
rect 2063 318 2076 364
rect 2216 318 2331 364
rect 2063 305 2331 318
rect 1459 184 1539 290
rect 1195 140 1315 184
rect 1419 140 1539 184
rect 1587 140 1707 290
rect 2063 185 2163 305
rect 2231 185 2331 305
rect 2492 352 3293 365
rect 2492 306 2505 352
rect 2927 311 3293 352
rect 2927 306 3323 311
rect 2492 292 3323 306
rect 2492 232 2612 292
rect 2755 232 2875 292
rect 2979 232 3099 292
rect 3203 232 3323 292
rect 2063 141 2183 185
rect 2231 141 2351 185
rect 179 24 299 68
rect 403 24 523 68
rect 571 24 691 68
rect 1027 24 1147 68
rect 1195 24 1315 68
rect 1419 24 1539 68
rect 1587 24 1707 68
rect 2063 24 2183 68
rect 2231 24 2351 68
rect 2492 24 2612 68
rect 2755 24 2875 68
rect 2979 24 3099 68
rect 3203 24 3323 68
<< polycontact >>
rect 192 257 238 303
rect 416 424 462 470
rect 596 424 642 470
rect 1020 304 1160 350
rect 1472 304 1612 350
rect 2076 318 2216 364
rect 2505 306 2927 352
<< metal1 >>
rect 0 724 3472 844
rect 297 703 365 724
rect 297 657 308 703
rect 354 657 365 703
rect 1293 703 1361 724
rect 1293 657 1304 703
rect 1350 657 1361 703
rect 2349 681 2417 724
rect 2349 635 2360 681
rect 2406 635 2417 681
rect 2893 681 2961 724
rect 744 621 790 632
rect 1780 621 1857 632
rect 49 575 60 621
rect 106 575 117 621
rect 49 481 117 575
rect 877 575 888 621
rect 934 575 1252 621
rect 49 470 653 481
rect 49 424 416 470
rect 462 424 596 470
rect 642 424 653 470
rect 49 413 653 424
rect 49 180 95 413
rect 744 361 790 575
rect 744 350 1160 361
rect 186 303 681 320
rect 186 257 192 303
rect 238 257 681 303
rect 186 240 681 257
rect 744 304 1020 350
rect 744 293 1160 304
rect 1206 350 1252 575
rect 1780 575 1800 621
rect 1846 575 1857 621
rect 1780 564 1857 575
rect 1944 621 1990 632
rect 1780 375 1826 564
rect 1944 493 1990 575
rect 2679 593 2690 639
rect 2736 593 2747 639
rect 2893 635 2904 681
rect 2950 635 2961 681
rect 3311 681 3379 724
rect 3108 639 3230 651
rect 2679 532 2747 593
rect 3154 593 3230 639
rect 3108 532 3230 593
rect 3311 541 3322 681
rect 3368 541 3379 681
rect 2679 531 3230 532
rect 1944 447 2338 493
rect 2679 485 2690 531
rect 2736 485 3108 531
rect 3154 485 3230 531
rect 1780 364 2216 375
rect 1206 304 1472 350
rect 1612 304 1623 350
rect 1780 318 2076 364
rect 1780 307 2216 318
rect 2274 352 2338 447
rect 744 200 821 293
rect 1206 200 1252 304
rect 49 134 60 180
rect 106 134 117 180
rect 744 154 764 200
rect 810 154 821 200
rect 897 154 908 200
rect 954 154 1252 200
rect 1780 200 1826 307
rect 2274 306 2505 352
rect 2927 306 2938 352
rect 2274 211 2338 306
rect 3108 231 3230 485
rect 1780 143 1826 154
rect 1944 200 2338 211
rect 1990 154 2338 200
rect 1944 143 2338 154
rect 2679 192 3230 231
rect 2679 146 2680 192
rect 2726 185 3128 192
rect 3108 146 3128 185
rect 3174 146 3230 192
rect 2385 128 2431 139
rect 2679 135 2726 146
rect 317 81 328 127
rect 374 81 385 127
rect 317 60 385 81
rect 1333 81 1344 127
rect 1390 81 1401 127
rect 1333 60 1401 81
rect 2385 60 2431 82
rect 2904 128 2950 139
rect 2904 60 2950 82
rect 3352 128 3398 139
rect 3352 60 3398 82
rect 0 -60 3472 60
<< labels >>
flabel metal1 s 3108 639 3230 651 0 FreeSans 400 0 0 0 Z
port 2 nsew default output
flabel metal1 s 3352 127 3398 139 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 186 240 681 320 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 3472 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 4 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 5 nsew ground bidirectional
rlabel metal1 s 3108 532 3230 639 1 Z
port 2 nsew default output
rlabel metal1 s 2679 532 2747 639 1 Z
port 2 nsew default output
rlabel metal1 s 2679 485 3230 532 1 Z
port 2 nsew default output
rlabel metal1 s 3108 231 3230 485 1 Z
port 2 nsew default output
rlabel metal1 s 2679 185 3230 231 1 Z
port 2 nsew default output
rlabel metal1 s 3108 146 3230 185 1 Z
port 2 nsew default output
rlabel metal1 s 2679 146 2726 185 1 Z
port 2 nsew default output
rlabel metal1 s 2679 135 2726 146 1 Z
port 2 nsew default output
rlabel metal1 s 3311 657 3379 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2893 657 2961 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2349 657 2417 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1293 657 1361 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3311 635 3379 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2893 635 2961 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2349 635 2417 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3311 541 3379 635 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2904 127 2950 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2385 127 2431 139 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3352 60 3398 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2904 60 2950 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2385 60 2431 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1333 60 1401 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3472 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 784
string GDS_END 1122016
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1115372
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
