magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< metal1 >>
rect -44 7318 200 7400
rect -44 7266 0 7318
rect 156 7266 200 7318
rect -44 7194 200 7266
rect -44 7142 0 7194
rect 156 7142 200 7194
rect -44 7070 200 7142
rect -44 7018 0 7070
rect 156 7018 200 7070
rect -44 6946 200 7018
rect -44 6894 0 6946
rect 156 6894 200 6946
rect -44 6822 200 6894
rect -44 6770 0 6822
rect 156 6770 200 6822
rect -44 6698 200 6770
rect -44 6646 0 6698
rect 156 6646 200 6698
rect -44 6574 200 6646
rect -44 6522 0 6574
rect 156 6522 200 6574
rect -44 6450 200 6522
rect -44 6398 0 6450
rect 156 6398 200 6450
rect -44 6326 200 6398
rect -44 6274 0 6326
rect 156 6274 200 6326
rect -44 6202 200 6274
rect -44 6150 0 6202
rect 156 6150 200 6202
rect -44 6078 200 6150
rect -44 6026 0 6078
rect 156 6026 200 6078
rect -44 5954 200 6026
rect -44 5902 0 5954
rect 156 5902 200 5954
rect -44 5830 200 5902
rect -44 5778 0 5830
rect 156 5778 200 5830
rect -44 5706 200 5778
rect -44 5654 0 5706
rect 156 5654 200 5706
rect -44 5582 200 5654
rect -44 5530 0 5582
rect 156 5530 200 5582
rect -44 5458 200 5530
rect -44 5406 0 5458
rect 156 5406 200 5458
rect -44 5334 200 5406
rect -44 5282 0 5334
rect 156 5282 200 5334
rect -44 5210 200 5282
rect -44 5158 0 5210
rect 156 5158 200 5210
rect -44 5086 200 5158
rect -44 5034 0 5086
rect 156 5034 200 5086
rect -44 4962 200 5034
rect -44 4910 0 4962
rect 156 4910 200 4962
rect -44 4838 200 4910
rect -44 4786 0 4838
rect 156 4786 200 4838
rect -44 4714 200 4786
rect -44 4662 0 4714
rect 156 4662 200 4714
rect -44 4590 200 4662
rect -44 4538 0 4590
rect 156 4538 200 4590
rect -44 4466 200 4538
rect -44 4414 0 4466
rect 156 4414 200 4466
rect -44 4342 200 4414
rect -44 4290 0 4342
rect 156 4290 200 4342
rect -44 4218 200 4290
rect -44 4166 0 4218
rect 156 4166 200 4218
rect -44 4094 200 4166
rect -44 4042 0 4094
rect 156 4042 200 4094
rect -44 3970 200 4042
rect -44 3918 0 3970
rect 156 3918 200 3970
rect -44 3846 200 3918
rect -44 3794 0 3846
rect 156 3794 200 3846
rect -44 3722 200 3794
rect -44 3670 0 3722
rect 156 3670 200 3722
rect -44 3598 200 3670
rect -44 3546 0 3598
rect 156 3546 200 3598
rect -44 3474 200 3546
rect -44 3422 0 3474
rect 156 3422 200 3474
rect -44 3350 200 3422
rect -44 3298 0 3350
rect 156 3298 200 3350
rect -44 3226 200 3298
rect -44 3174 0 3226
rect 156 3174 200 3226
rect -44 3102 200 3174
rect -44 3050 0 3102
rect 156 3050 200 3102
rect -44 2978 200 3050
rect -44 2926 0 2978
rect 156 2926 200 2978
rect -44 2854 200 2926
rect -44 2802 0 2854
rect 156 2802 200 2854
rect -44 2730 200 2802
rect -44 2678 0 2730
rect 156 2678 200 2730
rect -44 2606 200 2678
rect -44 2554 0 2606
rect 156 2554 200 2606
rect -44 2482 200 2554
rect -44 2430 0 2482
rect 156 2430 200 2482
rect -44 2358 200 2430
rect -44 2306 0 2358
rect 156 2306 200 2358
rect -44 2234 200 2306
rect -44 2182 0 2234
rect 156 2182 200 2234
rect -44 2110 200 2182
rect -44 2058 0 2110
rect 156 2058 200 2110
rect -44 1986 200 2058
rect -44 1934 0 1986
rect 156 1934 200 1986
rect -44 1862 200 1934
rect -44 1810 0 1862
rect 156 1810 200 1862
rect -44 1738 200 1810
rect -44 1686 0 1738
rect 156 1686 200 1738
rect -44 1614 200 1686
rect -44 1562 0 1614
rect 156 1562 200 1614
rect -44 1490 200 1562
rect -44 1438 0 1490
rect 156 1438 200 1490
rect -44 1366 200 1438
rect -44 1314 0 1366
rect 156 1314 200 1366
rect -44 1242 200 1314
rect -44 1190 0 1242
rect 156 1190 200 1242
rect -44 1118 200 1190
rect -44 1066 0 1118
rect 156 1066 200 1118
rect -44 994 200 1066
rect -44 942 0 994
rect 156 942 200 994
rect -44 870 200 942
rect -44 818 0 870
rect 156 818 200 870
rect -44 746 200 818
rect -44 694 0 746
rect 156 694 200 746
rect -44 622 200 694
rect -44 570 0 622
rect 156 570 200 622
rect -44 498 200 570
rect -44 446 0 498
rect 156 446 200 498
rect -44 374 200 446
rect -44 322 0 374
rect 156 322 200 374
rect -44 250 200 322
rect -44 198 0 250
rect 156 198 200 250
rect -44 126 200 198
rect -44 74 0 126
rect 156 74 200 126
rect -44 0 200 74
rect 360 7299 2004 7400
rect 360 7247 412 7299
rect 464 7247 536 7299
rect 588 7247 660 7299
rect 712 7247 784 7299
rect 836 7247 908 7299
rect 960 7247 1032 7299
rect 1084 7247 1156 7299
rect 1208 7247 1280 7299
rect 1332 7247 1404 7299
rect 1456 7247 1528 7299
rect 1580 7247 1652 7299
rect 1704 7247 1776 7299
rect 1828 7247 1900 7299
rect 1952 7247 2004 7299
rect 360 7175 2004 7247
rect 360 7123 412 7175
rect 464 7123 536 7175
rect 588 7123 660 7175
rect 712 7123 784 7175
rect 836 7123 908 7175
rect 960 7123 1032 7175
rect 1084 7123 1156 7175
rect 1208 7123 1280 7175
rect 1332 7123 1404 7175
rect 1456 7123 1528 7175
rect 1580 7123 1652 7175
rect 1704 7123 1776 7175
rect 1828 7123 1900 7175
rect 1952 7123 2004 7175
rect 360 7051 2004 7123
rect 360 6999 412 7051
rect 464 6999 536 7051
rect 588 6999 660 7051
rect 712 6999 784 7051
rect 836 6999 908 7051
rect 960 6999 1032 7051
rect 1084 6999 1156 7051
rect 1208 6999 1280 7051
rect 1332 6999 1404 7051
rect 1456 6999 1528 7051
rect 1580 6999 1652 7051
rect 1704 6999 1776 7051
rect 1828 6999 1900 7051
rect 1952 6999 2004 7051
rect 360 6927 2004 6999
rect 360 6875 412 6927
rect 464 6875 536 6927
rect 588 6875 660 6927
rect 712 6875 784 6927
rect 836 6875 908 6927
rect 960 6875 1032 6927
rect 1084 6875 1156 6927
rect 1208 6875 1280 6927
rect 1332 6875 1404 6927
rect 1456 6875 1528 6927
rect 1580 6875 1652 6927
rect 1704 6875 1776 6927
rect 1828 6875 1900 6927
rect 1952 6875 2004 6927
rect 360 6803 2004 6875
rect 360 6751 412 6803
rect 464 6751 536 6803
rect 588 6751 660 6803
rect 712 6751 784 6803
rect 836 6751 908 6803
rect 960 6751 1032 6803
rect 1084 6751 1156 6803
rect 1208 6751 1280 6803
rect 1332 6751 1404 6803
rect 1456 6751 1528 6803
rect 1580 6751 1652 6803
rect 1704 6751 1776 6803
rect 1828 6751 1900 6803
rect 1952 6751 2004 6803
rect 360 6679 2004 6751
rect 360 6627 412 6679
rect 464 6627 536 6679
rect 588 6627 660 6679
rect 712 6627 784 6679
rect 836 6627 908 6679
rect 960 6627 1032 6679
rect 1084 6627 1156 6679
rect 1208 6627 1280 6679
rect 1332 6627 1404 6679
rect 1456 6627 1528 6679
rect 1580 6627 1652 6679
rect 1704 6627 1776 6679
rect 1828 6627 1900 6679
rect 1952 6627 2004 6679
rect 360 6555 2004 6627
rect 360 6503 412 6555
rect 464 6503 536 6555
rect 588 6503 660 6555
rect 712 6503 784 6555
rect 836 6503 908 6555
rect 960 6503 1032 6555
rect 1084 6503 1156 6555
rect 1208 6503 1280 6555
rect 1332 6503 1404 6555
rect 1456 6503 1528 6555
rect 1580 6503 1652 6555
rect 1704 6503 1776 6555
rect 1828 6503 1900 6555
rect 1952 6503 2004 6555
rect 360 6431 2004 6503
rect 360 6379 412 6431
rect 464 6379 536 6431
rect 588 6379 660 6431
rect 712 6379 784 6431
rect 836 6379 908 6431
rect 960 6379 1032 6431
rect 1084 6379 1156 6431
rect 1208 6379 1280 6431
rect 1332 6379 1404 6431
rect 1456 6379 1528 6431
rect 1580 6379 1652 6431
rect 1704 6379 1776 6431
rect 1828 6379 1900 6431
rect 1952 6379 2004 6431
rect 360 6307 2004 6379
rect 360 6255 412 6307
rect 464 6255 536 6307
rect 588 6255 660 6307
rect 712 6255 784 6307
rect 836 6255 908 6307
rect 960 6255 1032 6307
rect 1084 6255 1156 6307
rect 1208 6255 1280 6307
rect 1332 6255 1404 6307
rect 1456 6255 1528 6307
rect 1580 6255 1652 6307
rect 1704 6255 1776 6307
rect 1828 6255 1900 6307
rect 1952 6255 2004 6307
rect 360 6183 2004 6255
rect 360 6131 412 6183
rect 464 6131 536 6183
rect 588 6131 660 6183
rect 712 6131 784 6183
rect 836 6131 908 6183
rect 960 6131 1032 6183
rect 1084 6131 1156 6183
rect 1208 6131 1280 6183
rect 1332 6131 1404 6183
rect 1456 6131 1528 6183
rect 1580 6131 1652 6183
rect 1704 6131 1776 6183
rect 1828 6131 1900 6183
rect 1952 6131 2004 6183
rect 360 6059 2004 6131
rect 360 6007 412 6059
rect 464 6007 536 6059
rect 588 6007 660 6059
rect 712 6007 784 6059
rect 836 6007 908 6059
rect 960 6007 1032 6059
rect 1084 6007 1156 6059
rect 1208 6007 1280 6059
rect 1332 6007 1404 6059
rect 1456 6007 1528 6059
rect 1580 6007 1652 6059
rect 1704 6007 1776 6059
rect 1828 6007 1900 6059
rect 1952 6007 2004 6059
rect 360 5935 2004 6007
rect 360 5883 412 5935
rect 464 5883 536 5935
rect 588 5883 660 5935
rect 712 5883 784 5935
rect 836 5883 908 5935
rect 960 5883 1032 5935
rect 1084 5883 1156 5935
rect 1208 5883 1280 5935
rect 1332 5883 1404 5935
rect 1456 5883 1528 5935
rect 1580 5883 1652 5935
rect 1704 5883 1776 5935
rect 1828 5883 1900 5935
rect 1952 5883 2004 5935
rect 360 5811 2004 5883
rect 360 5759 412 5811
rect 464 5759 536 5811
rect 588 5759 660 5811
rect 712 5759 784 5811
rect 836 5759 908 5811
rect 960 5759 1032 5811
rect 1084 5759 1156 5811
rect 1208 5759 1280 5811
rect 1332 5759 1404 5811
rect 1456 5759 1528 5811
rect 1580 5759 1652 5811
rect 1704 5759 1776 5811
rect 1828 5759 1900 5811
rect 1952 5759 2004 5811
rect 360 5687 2004 5759
rect 360 5635 412 5687
rect 464 5635 536 5687
rect 588 5635 660 5687
rect 712 5635 784 5687
rect 836 5635 908 5687
rect 960 5635 1032 5687
rect 1084 5635 1156 5687
rect 1208 5635 1280 5687
rect 1332 5635 1404 5687
rect 1456 5635 1528 5687
rect 1580 5635 1652 5687
rect 1704 5635 1776 5687
rect 1828 5635 1900 5687
rect 1952 5635 2004 5687
rect 360 5563 2004 5635
rect 360 5511 412 5563
rect 464 5511 536 5563
rect 588 5511 660 5563
rect 712 5511 784 5563
rect 836 5511 908 5563
rect 960 5511 1032 5563
rect 1084 5511 1156 5563
rect 1208 5511 1280 5563
rect 1332 5511 1404 5563
rect 1456 5511 1528 5563
rect 1580 5511 1652 5563
rect 1704 5511 1776 5563
rect 1828 5511 1900 5563
rect 1952 5511 2004 5563
rect 360 5439 2004 5511
rect 360 5387 412 5439
rect 464 5387 536 5439
rect 588 5387 660 5439
rect 712 5387 784 5439
rect 836 5387 908 5439
rect 960 5387 1032 5439
rect 1084 5387 1156 5439
rect 1208 5387 1280 5439
rect 1332 5387 1404 5439
rect 1456 5387 1528 5439
rect 1580 5387 1652 5439
rect 1704 5387 1776 5439
rect 1828 5387 1900 5439
rect 1952 5387 2004 5439
rect 360 5315 2004 5387
rect 360 5263 412 5315
rect 464 5263 536 5315
rect 588 5263 660 5315
rect 712 5263 784 5315
rect 836 5263 908 5315
rect 960 5263 1032 5315
rect 1084 5263 1156 5315
rect 1208 5263 1280 5315
rect 1332 5263 1404 5315
rect 1456 5263 1528 5315
rect 1580 5263 1652 5315
rect 1704 5263 1776 5315
rect 1828 5263 1900 5315
rect 1952 5263 2004 5315
rect 360 5191 2004 5263
rect 360 5139 412 5191
rect 464 5139 536 5191
rect 588 5139 660 5191
rect 712 5139 784 5191
rect 836 5139 908 5191
rect 960 5139 1032 5191
rect 1084 5139 1156 5191
rect 1208 5139 1280 5191
rect 1332 5139 1404 5191
rect 1456 5139 1528 5191
rect 1580 5139 1652 5191
rect 1704 5139 1776 5191
rect 1828 5139 1900 5191
rect 1952 5139 2004 5191
rect 360 5067 2004 5139
rect 360 5015 412 5067
rect 464 5015 536 5067
rect 588 5015 660 5067
rect 712 5015 784 5067
rect 836 5015 908 5067
rect 960 5015 1032 5067
rect 1084 5015 1156 5067
rect 1208 5015 1280 5067
rect 1332 5015 1404 5067
rect 1456 5015 1528 5067
rect 1580 5015 1652 5067
rect 1704 5015 1776 5067
rect 1828 5015 1900 5067
rect 1952 5015 2004 5067
rect 360 4943 2004 5015
rect 360 4891 412 4943
rect 464 4891 536 4943
rect 588 4891 660 4943
rect 712 4891 784 4943
rect 836 4891 908 4943
rect 960 4891 1032 4943
rect 1084 4891 1156 4943
rect 1208 4891 1280 4943
rect 1332 4891 1404 4943
rect 1456 4891 1528 4943
rect 1580 4891 1652 4943
rect 1704 4891 1776 4943
rect 1828 4891 1900 4943
rect 1952 4891 2004 4943
rect 360 4819 2004 4891
rect 360 4767 412 4819
rect 464 4767 536 4819
rect 588 4767 660 4819
rect 712 4767 784 4819
rect 836 4767 908 4819
rect 960 4767 1032 4819
rect 1084 4767 1156 4819
rect 1208 4767 1280 4819
rect 1332 4767 1404 4819
rect 1456 4767 1528 4819
rect 1580 4767 1652 4819
rect 1704 4767 1776 4819
rect 1828 4767 1900 4819
rect 1952 4767 2004 4819
rect 360 4695 2004 4767
rect 360 4643 412 4695
rect 464 4643 536 4695
rect 588 4643 660 4695
rect 712 4643 784 4695
rect 836 4643 908 4695
rect 960 4643 1032 4695
rect 1084 4643 1156 4695
rect 1208 4643 1280 4695
rect 1332 4643 1404 4695
rect 1456 4643 1528 4695
rect 1580 4643 1652 4695
rect 1704 4643 1776 4695
rect 1828 4643 1900 4695
rect 1952 4643 2004 4695
rect 360 4571 2004 4643
rect 360 4519 412 4571
rect 464 4519 536 4571
rect 588 4519 660 4571
rect 712 4519 784 4571
rect 836 4519 908 4571
rect 960 4519 1032 4571
rect 1084 4519 1156 4571
rect 1208 4519 1280 4571
rect 1332 4519 1404 4571
rect 1456 4519 1528 4571
rect 1580 4519 1652 4571
rect 1704 4519 1776 4571
rect 1828 4519 1900 4571
rect 1952 4519 2004 4571
rect 360 4447 2004 4519
rect 360 4395 412 4447
rect 464 4395 536 4447
rect 588 4395 660 4447
rect 712 4395 784 4447
rect 836 4395 908 4447
rect 960 4395 1032 4447
rect 1084 4395 1156 4447
rect 1208 4395 1280 4447
rect 1332 4395 1404 4447
rect 1456 4395 1528 4447
rect 1580 4395 1652 4447
rect 1704 4395 1776 4447
rect 1828 4395 1900 4447
rect 1952 4395 2004 4447
rect 360 4323 2004 4395
rect 360 4271 412 4323
rect 464 4271 536 4323
rect 588 4271 660 4323
rect 712 4271 784 4323
rect 836 4271 908 4323
rect 960 4271 1032 4323
rect 1084 4271 1156 4323
rect 1208 4271 1280 4323
rect 1332 4271 1404 4323
rect 1456 4271 1528 4323
rect 1580 4271 1652 4323
rect 1704 4271 1776 4323
rect 1828 4271 1900 4323
rect 1952 4271 2004 4323
rect 360 4199 2004 4271
rect 360 4147 412 4199
rect 464 4147 536 4199
rect 588 4147 660 4199
rect 712 4147 784 4199
rect 836 4147 908 4199
rect 960 4147 1032 4199
rect 1084 4147 1156 4199
rect 1208 4147 1280 4199
rect 1332 4147 1404 4199
rect 1456 4147 1528 4199
rect 1580 4147 1652 4199
rect 1704 4147 1776 4199
rect 1828 4147 1900 4199
rect 1952 4147 2004 4199
rect 360 4075 2004 4147
rect 360 4023 412 4075
rect 464 4023 536 4075
rect 588 4023 660 4075
rect 712 4023 784 4075
rect 836 4023 908 4075
rect 960 4023 1032 4075
rect 1084 4023 1156 4075
rect 1208 4023 1280 4075
rect 1332 4023 1404 4075
rect 1456 4023 1528 4075
rect 1580 4023 1652 4075
rect 1704 4023 1776 4075
rect 1828 4023 1900 4075
rect 1952 4023 2004 4075
rect 360 3951 2004 4023
rect 360 3899 412 3951
rect 464 3899 536 3951
rect 588 3899 660 3951
rect 712 3899 784 3951
rect 836 3899 908 3951
rect 960 3899 1032 3951
rect 1084 3899 1156 3951
rect 1208 3899 1280 3951
rect 1332 3899 1404 3951
rect 1456 3899 1528 3951
rect 1580 3899 1652 3951
rect 1704 3899 1776 3951
rect 1828 3899 1900 3951
rect 1952 3899 2004 3951
rect 360 3827 2004 3899
rect 360 3775 412 3827
rect 464 3775 536 3827
rect 588 3775 660 3827
rect 712 3775 784 3827
rect 836 3775 908 3827
rect 960 3775 1032 3827
rect 1084 3775 1156 3827
rect 1208 3775 1280 3827
rect 1332 3775 1404 3827
rect 1456 3775 1528 3827
rect 1580 3775 1652 3827
rect 1704 3775 1776 3827
rect 1828 3775 1900 3827
rect 1952 3775 2004 3827
rect 360 3703 2004 3775
rect 360 3651 412 3703
rect 464 3651 536 3703
rect 588 3651 660 3703
rect 712 3651 784 3703
rect 836 3651 908 3703
rect 960 3651 1032 3703
rect 1084 3651 1156 3703
rect 1208 3651 1280 3703
rect 1332 3651 1404 3703
rect 1456 3651 1528 3703
rect 1580 3651 1652 3703
rect 1704 3651 1776 3703
rect 1828 3651 1900 3703
rect 1952 3651 2004 3703
rect 360 3579 2004 3651
rect 360 3527 412 3579
rect 464 3527 536 3579
rect 588 3527 660 3579
rect 712 3527 784 3579
rect 836 3527 908 3579
rect 960 3527 1032 3579
rect 1084 3527 1156 3579
rect 1208 3527 1280 3579
rect 1332 3527 1404 3579
rect 1456 3527 1528 3579
rect 1580 3527 1652 3579
rect 1704 3527 1776 3579
rect 1828 3527 1900 3579
rect 1952 3527 2004 3579
rect 360 3455 2004 3527
rect 360 3403 412 3455
rect 464 3403 536 3455
rect 588 3403 660 3455
rect 712 3403 784 3455
rect 836 3403 908 3455
rect 960 3403 1032 3455
rect 1084 3403 1156 3455
rect 1208 3403 1280 3455
rect 1332 3403 1404 3455
rect 1456 3403 1528 3455
rect 1580 3403 1652 3455
rect 1704 3403 1776 3455
rect 1828 3403 1900 3455
rect 1952 3403 2004 3455
rect 360 3331 2004 3403
rect 360 3279 412 3331
rect 464 3279 536 3331
rect 588 3279 660 3331
rect 712 3279 784 3331
rect 836 3279 908 3331
rect 960 3279 1032 3331
rect 1084 3279 1156 3331
rect 1208 3279 1280 3331
rect 1332 3279 1404 3331
rect 1456 3279 1528 3331
rect 1580 3279 1652 3331
rect 1704 3279 1776 3331
rect 1828 3279 1900 3331
rect 1952 3279 2004 3331
rect 360 3207 2004 3279
rect 360 3155 412 3207
rect 464 3155 536 3207
rect 588 3155 660 3207
rect 712 3155 784 3207
rect 836 3155 908 3207
rect 960 3155 1032 3207
rect 1084 3155 1156 3207
rect 1208 3155 1280 3207
rect 1332 3155 1404 3207
rect 1456 3155 1528 3207
rect 1580 3155 1652 3207
rect 1704 3155 1776 3207
rect 1828 3155 1900 3207
rect 1952 3155 2004 3207
rect 360 3083 2004 3155
rect 360 3031 412 3083
rect 464 3031 536 3083
rect 588 3031 660 3083
rect 712 3031 784 3083
rect 836 3031 908 3083
rect 960 3031 1032 3083
rect 1084 3031 1156 3083
rect 1208 3031 1280 3083
rect 1332 3031 1404 3083
rect 1456 3031 1528 3083
rect 1580 3031 1652 3083
rect 1704 3031 1776 3083
rect 1828 3031 1900 3083
rect 1952 3031 2004 3083
rect 360 2959 2004 3031
rect 360 2907 412 2959
rect 464 2907 536 2959
rect 588 2907 660 2959
rect 712 2907 784 2959
rect 836 2907 908 2959
rect 960 2907 1032 2959
rect 1084 2907 1156 2959
rect 1208 2907 1280 2959
rect 1332 2907 1404 2959
rect 1456 2907 1528 2959
rect 1580 2907 1652 2959
rect 1704 2907 1776 2959
rect 1828 2907 1900 2959
rect 1952 2907 2004 2959
rect 360 2835 2004 2907
rect 360 2783 412 2835
rect 464 2783 536 2835
rect 588 2783 660 2835
rect 712 2783 784 2835
rect 836 2783 908 2835
rect 960 2783 1032 2835
rect 1084 2783 1156 2835
rect 1208 2783 1280 2835
rect 1332 2783 1404 2835
rect 1456 2783 1528 2835
rect 1580 2783 1652 2835
rect 1704 2783 1776 2835
rect 1828 2783 1900 2835
rect 1952 2783 2004 2835
rect 360 2711 2004 2783
rect 360 2659 412 2711
rect 464 2659 536 2711
rect 588 2659 660 2711
rect 712 2659 784 2711
rect 836 2659 908 2711
rect 960 2659 1032 2711
rect 1084 2659 1156 2711
rect 1208 2659 1280 2711
rect 1332 2659 1404 2711
rect 1456 2659 1528 2711
rect 1580 2659 1652 2711
rect 1704 2659 1776 2711
rect 1828 2659 1900 2711
rect 1952 2659 2004 2711
rect 360 2587 2004 2659
rect 360 2535 412 2587
rect 464 2535 536 2587
rect 588 2535 660 2587
rect 712 2535 784 2587
rect 836 2535 908 2587
rect 960 2535 1032 2587
rect 1084 2535 1156 2587
rect 1208 2535 1280 2587
rect 1332 2535 1404 2587
rect 1456 2535 1528 2587
rect 1580 2535 1652 2587
rect 1704 2535 1776 2587
rect 1828 2535 1900 2587
rect 1952 2535 2004 2587
rect 360 2463 2004 2535
rect 360 2411 412 2463
rect 464 2411 536 2463
rect 588 2411 660 2463
rect 712 2411 784 2463
rect 836 2411 908 2463
rect 960 2411 1032 2463
rect 1084 2411 1156 2463
rect 1208 2411 1280 2463
rect 1332 2411 1404 2463
rect 1456 2411 1528 2463
rect 1580 2411 1652 2463
rect 1704 2411 1776 2463
rect 1828 2411 1900 2463
rect 1952 2411 2004 2463
rect 360 2339 2004 2411
rect 360 2287 412 2339
rect 464 2287 536 2339
rect 588 2287 660 2339
rect 712 2287 784 2339
rect 836 2287 908 2339
rect 960 2287 1032 2339
rect 1084 2287 1156 2339
rect 1208 2287 1280 2339
rect 1332 2287 1404 2339
rect 1456 2287 1528 2339
rect 1580 2287 1652 2339
rect 1704 2287 1776 2339
rect 1828 2287 1900 2339
rect 1952 2287 2004 2339
rect 360 2215 2004 2287
rect 360 2163 412 2215
rect 464 2163 536 2215
rect 588 2163 660 2215
rect 712 2163 784 2215
rect 836 2163 908 2215
rect 960 2163 1032 2215
rect 1084 2163 1156 2215
rect 1208 2163 1280 2215
rect 1332 2163 1404 2215
rect 1456 2163 1528 2215
rect 1580 2163 1652 2215
rect 1704 2163 1776 2215
rect 1828 2163 1900 2215
rect 1952 2163 2004 2215
rect 360 2091 2004 2163
rect 360 2039 412 2091
rect 464 2039 536 2091
rect 588 2039 660 2091
rect 712 2039 784 2091
rect 836 2039 908 2091
rect 960 2039 1032 2091
rect 1084 2039 1156 2091
rect 1208 2039 1280 2091
rect 1332 2039 1404 2091
rect 1456 2039 1528 2091
rect 1580 2039 1652 2091
rect 1704 2039 1776 2091
rect 1828 2039 1900 2091
rect 1952 2039 2004 2091
rect 360 1967 2004 2039
rect 360 1915 412 1967
rect 464 1915 536 1967
rect 588 1915 660 1967
rect 712 1915 784 1967
rect 836 1915 908 1967
rect 960 1915 1032 1967
rect 1084 1915 1156 1967
rect 1208 1915 1280 1967
rect 1332 1915 1404 1967
rect 1456 1915 1528 1967
rect 1580 1915 1652 1967
rect 1704 1915 1776 1967
rect 1828 1915 1900 1967
rect 1952 1915 2004 1967
rect 360 1843 2004 1915
rect 360 1791 412 1843
rect 464 1791 536 1843
rect 588 1791 660 1843
rect 712 1791 784 1843
rect 836 1791 908 1843
rect 960 1791 1032 1843
rect 1084 1791 1156 1843
rect 1208 1791 1280 1843
rect 1332 1791 1404 1843
rect 1456 1791 1528 1843
rect 1580 1791 1652 1843
rect 1704 1791 1776 1843
rect 1828 1791 1900 1843
rect 1952 1791 2004 1843
rect 360 1719 2004 1791
rect 360 1667 412 1719
rect 464 1667 536 1719
rect 588 1667 660 1719
rect 712 1667 784 1719
rect 836 1667 908 1719
rect 960 1667 1032 1719
rect 1084 1667 1156 1719
rect 1208 1667 1280 1719
rect 1332 1667 1404 1719
rect 1456 1667 1528 1719
rect 1580 1667 1652 1719
rect 1704 1667 1776 1719
rect 1828 1667 1900 1719
rect 1952 1667 2004 1719
rect 360 1595 2004 1667
rect 360 1543 412 1595
rect 464 1543 536 1595
rect 588 1543 660 1595
rect 712 1543 784 1595
rect 836 1543 908 1595
rect 960 1543 1032 1595
rect 1084 1543 1156 1595
rect 1208 1543 1280 1595
rect 1332 1543 1404 1595
rect 1456 1543 1528 1595
rect 1580 1543 1652 1595
rect 1704 1543 1776 1595
rect 1828 1543 1900 1595
rect 1952 1543 2004 1595
rect 360 1471 2004 1543
rect 360 1419 412 1471
rect 464 1419 536 1471
rect 588 1419 660 1471
rect 712 1419 784 1471
rect 836 1419 908 1471
rect 960 1419 1032 1471
rect 1084 1419 1156 1471
rect 1208 1419 1280 1471
rect 1332 1419 1404 1471
rect 1456 1419 1528 1471
rect 1580 1419 1652 1471
rect 1704 1419 1776 1471
rect 1828 1419 1900 1471
rect 1952 1419 2004 1471
rect 360 1347 2004 1419
rect 360 1295 412 1347
rect 464 1295 536 1347
rect 588 1295 660 1347
rect 712 1295 784 1347
rect 836 1295 908 1347
rect 960 1295 1032 1347
rect 1084 1295 1156 1347
rect 1208 1295 1280 1347
rect 1332 1295 1404 1347
rect 1456 1295 1528 1347
rect 1580 1295 1652 1347
rect 1704 1295 1776 1347
rect 1828 1295 1900 1347
rect 1952 1295 2004 1347
rect 360 1223 2004 1295
rect 360 1171 412 1223
rect 464 1171 536 1223
rect 588 1171 660 1223
rect 712 1171 784 1223
rect 836 1171 908 1223
rect 960 1171 1032 1223
rect 1084 1171 1156 1223
rect 1208 1171 1280 1223
rect 1332 1171 1404 1223
rect 1456 1171 1528 1223
rect 1580 1171 1652 1223
rect 1704 1171 1776 1223
rect 1828 1171 1900 1223
rect 1952 1171 2004 1223
rect 360 1099 2004 1171
rect 360 1047 412 1099
rect 464 1047 536 1099
rect 588 1047 660 1099
rect 712 1047 784 1099
rect 836 1047 908 1099
rect 960 1047 1032 1099
rect 1084 1047 1156 1099
rect 1208 1047 1280 1099
rect 1332 1047 1404 1099
rect 1456 1047 1528 1099
rect 1580 1047 1652 1099
rect 1704 1047 1776 1099
rect 1828 1047 1900 1099
rect 1952 1047 2004 1099
rect 360 975 2004 1047
rect 360 923 412 975
rect 464 923 536 975
rect 588 923 660 975
rect 712 923 784 975
rect 836 923 908 975
rect 960 923 1032 975
rect 1084 923 1156 975
rect 1208 923 1280 975
rect 1332 923 1404 975
rect 1456 923 1528 975
rect 1580 923 1652 975
rect 1704 923 1776 975
rect 1828 923 1900 975
rect 1952 923 2004 975
rect 360 851 2004 923
rect 360 799 412 851
rect 464 799 536 851
rect 588 799 660 851
rect 712 799 784 851
rect 836 799 908 851
rect 960 799 1032 851
rect 1084 799 1156 851
rect 1208 799 1280 851
rect 1332 799 1404 851
rect 1456 799 1528 851
rect 1580 799 1652 851
rect 1704 799 1776 851
rect 1828 799 1900 851
rect 1952 799 2004 851
rect 360 727 2004 799
rect 360 675 412 727
rect 464 675 536 727
rect 588 675 660 727
rect 712 675 784 727
rect 836 675 908 727
rect 960 675 1032 727
rect 1084 675 1156 727
rect 1208 675 1280 727
rect 1332 675 1404 727
rect 1456 675 1528 727
rect 1580 675 1652 727
rect 1704 675 1776 727
rect 1828 675 1900 727
rect 1952 675 2004 727
rect 360 603 2004 675
rect 360 551 412 603
rect 464 551 536 603
rect 588 551 660 603
rect 712 551 784 603
rect 836 551 908 603
rect 960 551 1032 603
rect 1084 551 1156 603
rect 1208 551 1280 603
rect 1332 551 1404 603
rect 1456 551 1528 603
rect 1580 551 1652 603
rect 1704 551 1776 603
rect 1828 551 1900 603
rect 1952 551 2004 603
rect 360 479 2004 551
rect 360 427 412 479
rect 464 427 536 479
rect 588 427 660 479
rect 712 427 784 479
rect 836 427 908 479
rect 960 427 1032 479
rect 1084 427 1156 479
rect 1208 427 1280 479
rect 1332 427 1404 479
rect 1456 427 1528 479
rect 1580 427 1652 479
rect 1704 427 1776 479
rect 1828 427 1900 479
rect 1952 427 2004 479
rect 360 355 2004 427
rect 360 303 412 355
rect 464 303 536 355
rect 588 303 660 355
rect 712 303 784 355
rect 836 303 908 355
rect 960 303 1032 355
rect 1084 303 1156 355
rect 1208 303 1280 355
rect 1332 303 1404 355
rect 1456 303 1528 355
rect 1580 303 1652 355
rect 1704 303 1776 355
rect 1828 303 1900 355
rect 1952 303 2004 355
rect 360 231 2004 303
rect 360 179 412 231
rect 464 179 536 231
rect 588 179 660 231
rect 712 179 784 231
rect 836 179 908 231
rect 960 179 1032 231
rect 1084 179 1156 231
rect 1208 179 1280 231
rect 1332 179 1404 231
rect 1456 179 1528 231
rect 1580 179 1652 231
rect 1704 179 1776 231
rect 1828 179 1900 231
rect 1952 179 2004 231
rect 360 107 2004 179
rect 360 55 412 107
rect 464 55 536 107
rect 588 55 660 107
rect 712 55 784 107
rect 836 55 908 107
rect 960 55 1032 107
rect 1084 55 1156 107
rect 1208 55 1280 107
rect 1332 55 1404 107
rect 1456 55 1528 107
rect 1580 55 1652 107
rect 1704 55 1776 107
rect 1828 55 1900 107
rect 1952 55 2004 107
rect 360 0 2004 55
<< via1 >>
rect 0 7266 156 7318
rect 0 7142 156 7194
rect 0 7018 156 7070
rect 0 6894 156 6946
rect 0 6770 156 6822
rect 0 6646 156 6698
rect 0 6522 156 6574
rect 0 6398 156 6450
rect 0 6274 156 6326
rect 0 6150 156 6202
rect 0 6026 156 6078
rect 0 5902 156 5954
rect 0 5778 156 5830
rect 0 5654 156 5706
rect 0 5530 156 5582
rect 0 5406 156 5458
rect 0 5282 156 5334
rect 0 5158 156 5210
rect 0 5034 156 5086
rect 0 4910 156 4962
rect 0 4786 156 4838
rect 0 4662 156 4714
rect 0 4538 156 4590
rect 0 4414 156 4466
rect 0 4290 156 4342
rect 0 4166 156 4218
rect 0 4042 156 4094
rect 0 3918 156 3970
rect 0 3794 156 3846
rect 0 3670 156 3722
rect 0 3546 156 3598
rect 0 3422 156 3474
rect 0 3298 156 3350
rect 0 3174 156 3226
rect 0 3050 156 3102
rect 0 2926 156 2978
rect 0 2802 156 2854
rect 0 2678 156 2730
rect 0 2554 156 2606
rect 0 2430 156 2482
rect 0 2306 156 2358
rect 0 2182 156 2234
rect 0 2058 156 2110
rect 0 1934 156 1986
rect 0 1810 156 1862
rect 0 1686 156 1738
rect 0 1562 156 1614
rect 0 1438 156 1490
rect 0 1314 156 1366
rect 0 1190 156 1242
rect 0 1066 156 1118
rect 0 942 156 994
rect 0 818 156 870
rect 0 694 156 746
rect 0 570 156 622
rect 0 446 156 498
rect 0 322 156 374
rect 0 198 156 250
rect 0 74 156 126
rect 412 7247 464 7299
rect 536 7247 588 7299
rect 660 7247 712 7299
rect 784 7247 836 7299
rect 908 7247 960 7299
rect 1032 7247 1084 7299
rect 1156 7247 1208 7299
rect 1280 7247 1332 7299
rect 1404 7247 1456 7299
rect 1528 7247 1580 7299
rect 1652 7247 1704 7299
rect 1776 7247 1828 7299
rect 1900 7247 1952 7299
rect 412 7123 464 7175
rect 536 7123 588 7175
rect 660 7123 712 7175
rect 784 7123 836 7175
rect 908 7123 960 7175
rect 1032 7123 1084 7175
rect 1156 7123 1208 7175
rect 1280 7123 1332 7175
rect 1404 7123 1456 7175
rect 1528 7123 1580 7175
rect 1652 7123 1704 7175
rect 1776 7123 1828 7175
rect 1900 7123 1952 7175
rect 412 6999 464 7051
rect 536 6999 588 7051
rect 660 6999 712 7051
rect 784 6999 836 7051
rect 908 6999 960 7051
rect 1032 6999 1084 7051
rect 1156 6999 1208 7051
rect 1280 6999 1332 7051
rect 1404 6999 1456 7051
rect 1528 6999 1580 7051
rect 1652 6999 1704 7051
rect 1776 6999 1828 7051
rect 1900 6999 1952 7051
rect 412 6875 464 6927
rect 536 6875 588 6927
rect 660 6875 712 6927
rect 784 6875 836 6927
rect 908 6875 960 6927
rect 1032 6875 1084 6927
rect 1156 6875 1208 6927
rect 1280 6875 1332 6927
rect 1404 6875 1456 6927
rect 1528 6875 1580 6927
rect 1652 6875 1704 6927
rect 1776 6875 1828 6927
rect 1900 6875 1952 6927
rect 412 6751 464 6803
rect 536 6751 588 6803
rect 660 6751 712 6803
rect 784 6751 836 6803
rect 908 6751 960 6803
rect 1032 6751 1084 6803
rect 1156 6751 1208 6803
rect 1280 6751 1332 6803
rect 1404 6751 1456 6803
rect 1528 6751 1580 6803
rect 1652 6751 1704 6803
rect 1776 6751 1828 6803
rect 1900 6751 1952 6803
rect 412 6627 464 6679
rect 536 6627 588 6679
rect 660 6627 712 6679
rect 784 6627 836 6679
rect 908 6627 960 6679
rect 1032 6627 1084 6679
rect 1156 6627 1208 6679
rect 1280 6627 1332 6679
rect 1404 6627 1456 6679
rect 1528 6627 1580 6679
rect 1652 6627 1704 6679
rect 1776 6627 1828 6679
rect 1900 6627 1952 6679
rect 412 6503 464 6555
rect 536 6503 588 6555
rect 660 6503 712 6555
rect 784 6503 836 6555
rect 908 6503 960 6555
rect 1032 6503 1084 6555
rect 1156 6503 1208 6555
rect 1280 6503 1332 6555
rect 1404 6503 1456 6555
rect 1528 6503 1580 6555
rect 1652 6503 1704 6555
rect 1776 6503 1828 6555
rect 1900 6503 1952 6555
rect 412 6379 464 6431
rect 536 6379 588 6431
rect 660 6379 712 6431
rect 784 6379 836 6431
rect 908 6379 960 6431
rect 1032 6379 1084 6431
rect 1156 6379 1208 6431
rect 1280 6379 1332 6431
rect 1404 6379 1456 6431
rect 1528 6379 1580 6431
rect 1652 6379 1704 6431
rect 1776 6379 1828 6431
rect 1900 6379 1952 6431
rect 412 6255 464 6307
rect 536 6255 588 6307
rect 660 6255 712 6307
rect 784 6255 836 6307
rect 908 6255 960 6307
rect 1032 6255 1084 6307
rect 1156 6255 1208 6307
rect 1280 6255 1332 6307
rect 1404 6255 1456 6307
rect 1528 6255 1580 6307
rect 1652 6255 1704 6307
rect 1776 6255 1828 6307
rect 1900 6255 1952 6307
rect 412 6131 464 6183
rect 536 6131 588 6183
rect 660 6131 712 6183
rect 784 6131 836 6183
rect 908 6131 960 6183
rect 1032 6131 1084 6183
rect 1156 6131 1208 6183
rect 1280 6131 1332 6183
rect 1404 6131 1456 6183
rect 1528 6131 1580 6183
rect 1652 6131 1704 6183
rect 1776 6131 1828 6183
rect 1900 6131 1952 6183
rect 412 6007 464 6059
rect 536 6007 588 6059
rect 660 6007 712 6059
rect 784 6007 836 6059
rect 908 6007 960 6059
rect 1032 6007 1084 6059
rect 1156 6007 1208 6059
rect 1280 6007 1332 6059
rect 1404 6007 1456 6059
rect 1528 6007 1580 6059
rect 1652 6007 1704 6059
rect 1776 6007 1828 6059
rect 1900 6007 1952 6059
rect 412 5883 464 5935
rect 536 5883 588 5935
rect 660 5883 712 5935
rect 784 5883 836 5935
rect 908 5883 960 5935
rect 1032 5883 1084 5935
rect 1156 5883 1208 5935
rect 1280 5883 1332 5935
rect 1404 5883 1456 5935
rect 1528 5883 1580 5935
rect 1652 5883 1704 5935
rect 1776 5883 1828 5935
rect 1900 5883 1952 5935
rect 412 5759 464 5811
rect 536 5759 588 5811
rect 660 5759 712 5811
rect 784 5759 836 5811
rect 908 5759 960 5811
rect 1032 5759 1084 5811
rect 1156 5759 1208 5811
rect 1280 5759 1332 5811
rect 1404 5759 1456 5811
rect 1528 5759 1580 5811
rect 1652 5759 1704 5811
rect 1776 5759 1828 5811
rect 1900 5759 1952 5811
rect 412 5635 464 5687
rect 536 5635 588 5687
rect 660 5635 712 5687
rect 784 5635 836 5687
rect 908 5635 960 5687
rect 1032 5635 1084 5687
rect 1156 5635 1208 5687
rect 1280 5635 1332 5687
rect 1404 5635 1456 5687
rect 1528 5635 1580 5687
rect 1652 5635 1704 5687
rect 1776 5635 1828 5687
rect 1900 5635 1952 5687
rect 412 5511 464 5563
rect 536 5511 588 5563
rect 660 5511 712 5563
rect 784 5511 836 5563
rect 908 5511 960 5563
rect 1032 5511 1084 5563
rect 1156 5511 1208 5563
rect 1280 5511 1332 5563
rect 1404 5511 1456 5563
rect 1528 5511 1580 5563
rect 1652 5511 1704 5563
rect 1776 5511 1828 5563
rect 1900 5511 1952 5563
rect 412 5387 464 5439
rect 536 5387 588 5439
rect 660 5387 712 5439
rect 784 5387 836 5439
rect 908 5387 960 5439
rect 1032 5387 1084 5439
rect 1156 5387 1208 5439
rect 1280 5387 1332 5439
rect 1404 5387 1456 5439
rect 1528 5387 1580 5439
rect 1652 5387 1704 5439
rect 1776 5387 1828 5439
rect 1900 5387 1952 5439
rect 412 5263 464 5315
rect 536 5263 588 5315
rect 660 5263 712 5315
rect 784 5263 836 5315
rect 908 5263 960 5315
rect 1032 5263 1084 5315
rect 1156 5263 1208 5315
rect 1280 5263 1332 5315
rect 1404 5263 1456 5315
rect 1528 5263 1580 5315
rect 1652 5263 1704 5315
rect 1776 5263 1828 5315
rect 1900 5263 1952 5315
rect 412 5139 464 5191
rect 536 5139 588 5191
rect 660 5139 712 5191
rect 784 5139 836 5191
rect 908 5139 960 5191
rect 1032 5139 1084 5191
rect 1156 5139 1208 5191
rect 1280 5139 1332 5191
rect 1404 5139 1456 5191
rect 1528 5139 1580 5191
rect 1652 5139 1704 5191
rect 1776 5139 1828 5191
rect 1900 5139 1952 5191
rect 412 5015 464 5067
rect 536 5015 588 5067
rect 660 5015 712 5067
rect 784 5015 836 5067
rect 908 5015 960 5067
rect 1032 5015 1084 5067
rect 1156 5015 1208 5067
rect 1280 5015 1332 5067
rect 1404 5015 1456 5067
rect 1528 5015 1580 5067
rect 1652 5015 1704 5067
rect 1776 5015 1828 5067
rect 1900 5015 1952 5067
rect 412 4891 464 4943
rect 536 4891 588 4943
rect 660 4891 712 4943
rect 784 4891 836 4943
rect 908 4891 960 4943
rect 1032 4891 1084 4943
rect 1156 4891 1208 4943
rect 1280 4891 1332 4943
rect 1404 4891 1456 4943
rect 1528 4891 1580 4943
rect 1652 4891 1704 4943
rect 1776 4891 1828 4943
rect 1900 4891 1952 4943
rect 412 4767 464 4819
rect 536 4767 588 4819
rect 660 4767 712 4819
rect 784 4767 836 4819
rect 908 4767 960 4819
rect 1032 4767 1084 4819
rect 1156 4767 1208 4819
rect 1280 4767 1332 4819
rect 1404 4767 1456 4819
rect 1528 4767 1580 4819
rect 1652 4767 1704 4819
rect 1776 4767 1828 4819
rect 1900 4767 1952 4819
rect 412 4643 464 4695
rect 536 4643 588 4695
rect 660 4643 712 4695
rect 784 4643 836 4695
rect 908 4643 960 4695
rect 1032 4643 1084 4695
rect 1156 4643 1208 4695
rect 1280 4643 1332 4695
rect 1404 4643 1456 4695
rect 1528 4643 1580 4695
rect 1652 4643 1704 4695
rect 1776 4643 1828 4695
rect 1900 4643 1952 4695
rect 412 4519 464 4571
rect 536 4519 588 4571
rect 660 4519 712 4571
rect 784 4519 836 4571
rect 908 4519 960 4571
rect 1032 4519 1084 4571
rect 1156 4519 1208 4571
rect 1280 4519 1332 4571
rect 1404 4519 1456 4571
rect 1528 4519 1580 4571
rect 1652 4519 1704 4571
rect 1776 4519 1828 4571
rect 1900 4519 1952 4571
rect 412 4395 464 4447
rect 536 4395 588 4447
rect 660 4395 712 4447
rect 784 4395 836 4447
rect 908 4395 960 4447
rect 1032 4395 1084 4447
rect 1156 4395 1208 4447
rect 1280 4395 1332 4447
rect 1404 4395 1456 4447
rect 1528 4395 1580 4447
rect 1652 4395 1704 4447
rect 1776 4395 1828 4447
rect 1900 4395 1952 4447
rect 412 4271 464 4323
rect 536 4271 588 4323
rect 660 4271 712 4323
rect 784 4271 836 4323
rect 908 4271 960 4323
rect 1032 4271 1084 4323
rect 1156 4271 1208 4323
rect 1280 4271 1332 4323
rect 1404 4271 1456 4323
rect 1528 4271 1580 4323
rect 1652 4271 1704 4323
rect 1776 4271 1828 4323
rect 1900 4271 1952 4323
rect 412 4147 464 4199
rect 536 4147 588 4199
rect 660 4147 712 4199
rect 784 4147 836 4199
rect 908 4147 960 4199
rect 1032 4147 1084 4199
rect 1156 4147 1208 4199
rect 1280 4147 1332 4199
rect 1404 4147 1456 4199
rect 1528 4147 1580 4199
rect 1652 4147 1704 4199
rect 1776 4147 1828 4199
rect 1900 4147 1952 4199
rect 412 4023 464 4075
rect 536 4023 588 4075
rect 660 4023 712 4075
rect 784 4023 836 4075
rect 908 4023 960 4075
rect 1032 4023 1084 4075
rect 1156 4023 1208 4075
rect 1280 4023 1332 4075
rect 1404 4023 1456 4075
rect 1528 4023 1580 4075
rect 1652 4023 1704 4075
rect 1776 4023 1828 4075
rect 1900 4023 1952 4075
rect 412 3899 464 3951
rect 536 3899 588 3951
rect 660 3899 712 3951
rect 784 3899 836 3951
rect 908 3899 960 3951
rect 1032 3899 1084 3951
rect 1156 3899 1208 3951
rect 1280 3899 1332 3951
rect 1404 3899 1456 3951
rect 1528 3899 1580 3951
rect 1652 3899 1704 3951
rect 1776 3899 1828 3951
rect 1900 3899 1952 3951
rect 412 3775 464 3827
rect 536 3775 588 3827
rect 660 3775 712 3827
rect 784 3775 836 3827
rect 908 3775 960 3827
rect 1032 3775 1084 3827
rect 1156 3775 1208 3827
rect 1280 3775 1332 3827
rect 1404 3775 1456 3827
rect 1528 3775 1580 3827
rect 1652 3775 1704 3827
rect 1776 3775 1828 3827
rect 1900 3775 1952 3827
rect 412 3651 464 3703
rect 536 3651 588 3703
rect 660 3651 712 3703
rect 784 3651 836 3703
rect 908 3651 960 3703
rect 1032 3651 1084 3703
rect 1156 3651 1208 3703
rect 1280 3651 1332 3703
rect 1404 3651 1456 3703
rect 1528 3651 1580 3703
rect 1652 3651 1704 3703
rect 1776 3651 1828 3703
rect 1900 3651 1952 3703
rect 412 3527 464 3579
rect 536 3527 588 3579
rect 660 3527 712 3579
rect 784 3527 836 3579
rect 908 3527 960 3579
rect 1032 3527 1084 3579
rect 1156 3527 1208 3579
rect 1280 3527 1332 3579
rect 1404 3527 1456 3579
rect 1528 3527 1580 3579
rect 1652 3527 1704 3579
rect 1776 3527 1828 3579
rect 1900 3527 1952 3579
rect 412 3403 464 3455
rect 536 3403 588 3455
rect 660 3403 712 3455
rect 784 3403 836 3455
rect 908 3403 960 3455
rect 1032 3403 1084 3455
rect 1156 3403 1208 3455
rect 1280 3403 1332 3455
rect 1404 3403 1456 3455
rect 1528 3403 1580 3455
rect 1652 3403 1704 3455
rect 1776 3403 1828 3455
rect 1900 3403 1952 3455
rect 412 3279 464 3331
rect 536 3279 588 3331
rect 660 3279 712 3331
rect 784 3279 836 3331
rect 908 3279 960 3331
rect 1032 3279 1084 3331
rect 1156 3279 1208 3331
rect 1280 3279 1332 3331
rect 1404 3279 1456 3331
rect 1528 3279 1580 3331
rect 1652 3279 1704 3331
rect 1776 3279 1828 3331
rect 1900 3279 1952 3331
rect 412 3155 464 3207
rect 536 3155 588 3207
rect 660 3155 712 3207
rect 784 3155 836 3207
rect 908 3155 960 3207
rect 1032 3155 1084 3207
rect 1156 3155 1208 3207
rect 1280 3155 1332 3207
rect 1404 3155 1456 3207
rect 1528 3155 1580 3207
rect 1652 3155 1704 3207
rect 1776 3155 1828 3207
rect 1900 3155 1952 3207
rect 412 3031 464 3083
rect 536 3031 588 3083
rect 660 3031 712 3083
rect 784 3031 836 3083
rect 908 3031 960 3083
rect 1032 3031 1084 3083
rect 1156 3031 1208 3083
rect 1280 3031 1332 3083
rect 1404 3031 1456 3083
rect 1528 3031 1580 3083
rect 1652 3031 1704 3083
rect 1776 3031 1828 3083
rect 1900 3031 1952 3083
rect 412 2907 464 2959
rect 536 2907 588 2959
rect 660 2907 712 2959
rect 784 2907 836 2959
rect 908 2907 960 2959
rect 1032 2907 1084 2959
rect 1156 2907 1208 2959
rect 1280 2907 1332 2959
rect 1404 2907 1456 2959
rect 1528 2907 1580 2959
rect 1652 2907 1704 2959
rect 1776 2907 1828 2959
rect 1900 2907 1952 2959
rect 412 2783 464 2835
rect 536 2783 588 2835
rect 660 2783 712 2835
rect 784 2783 836 2835
rect 908 2783 960 2835
rect 1032 2783 1084 2835
rect 1156 2783 1208 2835
rect 1280 2783 1332 2835
rect 1404 2783 1456 2835
rect 1528 2783 1580 2835
rect 1652 2783 1704 2835
rect 1776 2783 1828 2835
rect 1900 2783 1952 2835
rect 412 2659 464 2711
rect 536 2659 588 2711
rect 660 2659 712 2711
rect 784 2659 836 2711
rect 908 2659 960 2711
rect 1032 2659 1084 2711
rect 1156 2659 1208 2711
rect 1280 2659 1332 2711
rect 1404 2659 1456 2711
rect 1528 2659 1580 2711
rect 1652 2659 1704 2711
rect 1776 2659 1828 2711
rect 1900 2659 1952 2711
rect 412 2535 464 2587
rect 536 2535 588 2587
rect 660 2535 712 2587
rect 784 2535 836 2587
rect 908 2535 960 2587
rect 1032 2535 1084 2587
rect 1156 2535 1208 2587
rect 1280 2535 1332 2587
rect 1404 2535 1456 2587
rect 1528 2535 1580 2587
rect 1652 2535 1704 2587
rect 1776 2535 1828 2587
rect 1900 2535 1952 2587
rect 412 2411 464 2463
rect 536 2411 588 2463
rect 660 2411 712 2463
rect 784 2411 836 2463
rect 908 2411 960 2463
rect 1032 2411 1084 2463
rect 1156 2411 1208 2463
rect 1280 2411 1332 2463
rect 1404 2411 1456 2463
rect 1528 2411 1580 2463
rect 1652 2411 1704 2463
rect 1776 2411 1828 2463
rect 1900 2411 1952 2463
rect 412 2287 464 2339
rect 536 2287 588 2339
rect 660 2287 712 2339
rect 784 2287 836 2339
rect 908 2287 960 2339
rect 1032 2287 1084 2339
rect 1156 2287 1208 2339
rect 1280 2287 1332 2339
rect 1404 2287 1456 2339
rect 1528 2287 1580 2339
rect 1652 2287 1704 2339
rect 1776 2287 1828 2339
rect 1900 2287 1952 2339
rect 412 2163 464 2215
rect 536 2163 588 2215
rect 660 2163 712 2215
rect 784 2163 836 2215
rect 908 2163 960 2215
rect 1032 2163 1084 2215
rect 1156 2163 1208 2215
rect 1280 2163 1332 2215
rect 1404 2163 1456 2215
rect 1528 2163 1580 2215
rect 1652 2163 1704 2215
rect 1776 2163 1828 2215
rect 1900 2163 1952 2215
rect 412 2039 464 2091
rect 536 2039 588 2091
rect 660 2039 712 2091
rect 784 2039 836 2091
rect 908 2039 960 2091
rect 1032 2039 1084 2091
rect 1156 2039 1208 2091
rect 1280 2039 1332 2091
rect 1404 2039 1456 2091
rect 1528 2039 1580 2091
rect 1652 2039 1704 2091
rect 1776 2039 1828 2091
rect 1900 2039 1952 2091
rect 412 1915 464 1967
rect 536 1915 588 1967
rect 660 1915 712 1967
rect 784 1915 836 1967
rect 908 1915 960 1967
rect 1032 1915 1084 1967
rect 1156 1915 1208 1967
rect 1280 1915 1332 1967
rect 1404 1915 1456 1967
rect 1528 1915 1580 1967
rect 1652 1915 1704 1967
rect 1776 1915 1828 1967
rect 1900 1915 1952 1967
rect 412 1791 464 1843
rect 536 1791 588 1843
rect 660 1791 712 1843
rect 784 1791 836 1843
rect 908 1791 960 1843
rect 1032 1791 1084 1843
rect 1156 1791 1208 1843
rect 1280 1791 1332 1843
rect 1404 1791 1456 1843
rect 1528 1791 1580 1843
rect 1652 1791 1704 1843
rect 1776 1791 1828 1843
rect 1900 1791 1952 1843
rect 412 1667 464 1719
rect 536 1667 588 1719
rect 660 1667 712 1719
rect 784 1667 836 1719
rect 908 1667 960 1719
rect 1032 1667 1084 1719
rect 1156 1667 1208 1719
rect 1280 1667 1332 1719
rect 1404 1667 1456 1719
rect 1528 1667 1580 1719
rect 1652 1667 1704 1719
rect 1776 1667 1828 1719
rect 1900 1667 1952 1719
rect 412 1543 464 1595
rect 536 1543 588 1595
rect 660 1543 712 1595
rect 784 1543 836 1595
rect 908 1543 960 1595
rect 1032 1543 1084 1595
rect 1156 1543 1208 1595
rect 1280 1543 1332 1595
rect 1404 1543 1456 1595
rect 1528 1543 1580 1595
rect 1652 1543 1704 1595
rect 1776 1543 1828 1595
rect 1900 1543 1952 1595
rect 412 1419 464 1471
rect 536 1419 588 1471
rect 660 1419 712 1471
rect 784 1419 836 1471
rect 908 1419 960 1471
rect 1032 1419 1084 1471
rect 1156 1419 1208 1471
rect 1280 1419 1332 1471
rect 1404 1419 1456 1471
rect 1528 1419 1580 1471
rect 1652 1419 1704 1471
rect 1776 1419 1828 1471
rect 1900 1419 1952 1471
rect 412 1295 464 1347
rect 536 1295 588 1347
rect 660 1295 712 1347
rect 784 1295 836 1347
rect 908 1295 960 1347
rect 1032 1295 1084 1347
rect 1156 1295 1208 1347
rect 1280 1295 1332 1347
rect 1404 1295 1456 1347
rect 1528 1295 1580 1347
rect 1652 1295 1704 1347
rect 1776 1295 1828 1347
rect 1900 1295 1952 1347
rect 412 1171 464 1223
rect 536 1171 588 1223
rect 660 1171 712 1223
rect 784 1171 836 1223
rect 908 1171 960 1223
rect 1032 1171 1084 1223
rect 1156 1171 1208 1223
rect 1280 1171 1332 1223
rect 1404 1171 1456 1223
rect 1528 1171 1580 1223
rect 1652 1171 1704 1223
rect 1776 1171 1828 1223
rect 1900 1171 1952 1223
rect 412 1047 464 1099
rect 536 1047 588 1099
rect 660 1047 712 1099
rect 784 1047 836 1099
rect 908 1047 960 1099
rect 1032 1047 1084 1099
rect 1156 1047 1208 1099
rect 1280 1047 1332 1099
rect 1404 1047 1456 1099
rect 1528 1047 1580 1099
rect 1652 1047 1704 1099
rect 1776 1047 1828 1099
rect 1900 1047 1952 1099
rect 412 923 464 975
rect 536 923 588 975
rect 660 923 712 975
rect 784 923 836 975
rect 908 923 960 975
rect 1032 923 1084 975
rect 1156 923 1208 975
rect 1280 923 1332 975
rect 1404 923 1456 975
rect 1528 923 1580 975
rect 1652 923 1704 975
rect 1776 923 1828 975
rect 1900 923 1952 975
rect 412 799 464 851
rect 536 799 588 851
rect 660 799 712 851
rect 784 799 836 851
rect 908 799 960 851
rect 1032 799 1084 851
rect 1156 799 1208 851
rect 1280 799 1332 851
rect 1404 799 1456 851
rect 1528 799 1580 851
rect 1652 799 1704 851
rect 1776 799 1828 851
rect 1900 799 1952 851
rect 412 675 464 727
rect 536 675 588 727
rect 660 675 712 727
rect 784 675 836 727
rect 908 675 960 727
rect 1032 675 1084 727
rect 1156 675 1208 727
rect 1280 675 1332 727
rect 1404 675 1456 727
rect 1528 675 1580 727
rect 1652 675 1704 727
rect 1776 675 1828 727
rect 1900 675 1952 727
rect 412 551 464 603
rect 536 551 588 603
rect 660 551 712 603
rect 784 551 836 603
rect 908 551 960 603
rect 1032 551 1084 603
rect 1156 551 1208 603
rect 1280 551 1332 603
rect 1404 551 1456 603
rect 1528 551 1580 603
rect 1652 551 1704 603
rect 1776 551 1828 603
rect 1900 551 1952 603
rect 412 427 464 479
rect 536 427 588 479
rect 660 427 712 479
rect 784 427 836 479
rect 908 427 960 479
rect 1032 427 1084 479
rect 1156 427 1208 479
rect 1280 427 1332 479
rect 1404 427 1456 479
rect 1528 427 1580 479
rect 1652 427 1704 479
rect 1776 427 1828 479
rect 1900 427 1952 479
rect 412 303 464 355
rect 536 303 588 355
rect 660 303 712 355
rect 784 303 836 355
rect 908 303 960 355
rect 1032 303 1084 355
rect 1156 303 1208 355
rect 1280 303 1332 355
rect 1404 303 1456 355
rect 1528 303 1580 355
rect 1652 303 1704 355
rect 1776 303 1828 355
rect 1900 303 1952 355
rect 412 179 464 231
rect 536 179 588 231
rect 660 179 712 231
rect 784 179 836 231
rect 908 179 960 231
rect 1032 179 1084 231
rect 1156 179 1208 231
rect 1280 179 1332 231
rect 1404 179 1456 231
rect 1528 179 1580 231
rect 1652 179 1704 231
rect 1776 179 1828 231
rect 1900 179 1952 231
rect 412 55 464 107
rect 536 55 588 107
rect 660 55 712 107
rect 784 55 836 107
rect 908 55 960 107
rect 1032 55 1084 107
rect 1156 55 1208 107
rect 1280 55 1332 107
rect 1404 55 1456 107
rect 1528 55 1580 107
rect 1652 55 1704 107
rect 1776 55 1828 107
rect 1900 55 1952 107
<< metal2 >>
rect -44 7318 200 7400
rect -44 7307 0 7318
rect 156 7307 200 7318
rect -44 7251 -2 7307
rect 158 7251 200 7307
rect -44 7194 200 7251
rect -44 7183 0 7194
rect 156 7183 200 7194
rect -44 7127 -2 7183
rect 158 7127 200 7183
rect -44 7070 200 7127
rect -44 7059 0 7070
rect 156 7059 200 7070
rect -44 7003 -2 7059
rect 158 7003 200 7059
rect -44 6946 200 7003
rect -44 6935 0 6946
rect 156 6935 200 6946
rect -44 6879 -2 6935
rect 158 6879 200 6935
rect -44 6822 200 6879
rect -44 6811 0 6822
rect 156 6811 200 6822
rect -44 6755 -2 6811
rect 158 6755 200 6811
rect -44 6698 200 6755
rect -44 6687 0 6698
rect 156 6687 200 6698
rect -44 6631 -2 6687
rect 158 6631 200 6687
rect -44 6574 200 6631
rect -44 6563 0 6574
rect 156 6563 200 6574
rect -44 6507 -2 6563
rect 158 6507 200 6563
rect -44 6450 200 6507
rect -44 6439 0 6450
rect 156 6439 200 6450
rect -44 6383 -2 6439
rect 158 6383 200 6439
rect -44 6326 200 6383
rect -44 6315 0 6326
rect 156 6315 200 6326
rect -44 6259 -2 6315
rect 158 6259 200 6315
rect -44 6202 200 6259
rect -44 6191 0 6202
rect 156 6191 200 6202
rect -44 6135 -2 6191
rect 158 6135 200 6191
rect -44 6078 200 6135
rect -44 6067 0 6078
rect 156 6067 200 6078
rect -44 6011 -2 6067
rect 158 6011 200 6067
rect -44 5954 200 6011
rect -44 5943 0 5954
rect 156 5943 200 5954
rect -44 5887 -2 5943
rect 158 5887 200 5943
rect -44 5830 200 5887
rect -44 5819 0 5830
rect 156 5819 200 5830
rect -44 5763 -2 5819
rect 158 5763 200 5819
rect -44 5706 200 5763
rect -44 5654 0 5706
rect 156 5654 200 5706
rect -44 5582 200 5654
rect -44 5530 0 5582
rect 156 5530 200 5582
rect -44 5458 200 5530
rect -44 5456 0 5458
rect 156 5456 200 5458
rect -44 5400 -2 5456
rect 158 5400 200 5456
rect -44 5334 200 5400
rect -44 5332 0 5334
rect 156 5332 200 5334
rect -44 5276 -2 5332
rect 158 5276 200 5332
rect -44 5210 200 5276
rect -44 5208 0 5210
rect 156 5208 200 5210
rect -44 5152 -2 5208
rect 158 5152 200 5208
rect -44 5086 200 5152
rect -44 5084 0 5086
rect 156 5084 200 5086
rect -44 5028 -2 5084
rect 158 5028 200 5084
rect -44 4962 200 5028
rect -44 4960 0 4962
rect 156 4960 200 4962
rect -44 4904 -2 4960
rect 158 4904 200 4960
rect -44 4838 200 4904
rect -44 4836 0 4838
rect 156 4836 200 4838
rect -44 4780 -2 4836
rect 158 4780 200 4836
rect -44 4714 200 4780
rect -44 4712 0 4714
rect 156 4712 200 4714
rect -44 4656 -2 4712
rect 158 4656 200 4712
rect -44 4590 200 4656
rect -44 4588 0 4590
rect 156 4588 200 4590
rect -44 4532 -2 4588
rect 158 4532 200 4588
rect -44 4466 200 4532
rect -44 4464 0 4466
rect 156 4464 200 4466
rect -44 4408 -2 4464
rect 158 4408 200 4464
rect -44 4342 200 4408
rect -44 4340 0 4342
rect 156 4340 200 4342
rect -44 4284 -2 4340
rect 158 4284 200 4340
rect -44 4218 200 4284
rect -44 4216 0 4218
rect 156 4216 200 4218
rect -44 4160 -2 4216
rect 158 4160 200 4216
rect -44 4094 200 4160
rect -44 4092 0 4094
rect 156 4092 200 4094
rect -44 4036 -2 4092
rect 158 4036 200 4092
rect -44 3970 200 4036
rect -44 3968 0 3970
rect 156 3968 200 3970
rect -44 3912 -2 3968
rect 158 3912 200 3968
rect -44 3846 200 3912
rect -44 3844 0 3846
rect 156 3844 200 3846
rect -44 3788 -2 3844
rect 158 3788 200 3844
rect -44 3722 200 3788
rect -44 3720 0 3722
rect 156 3720 200 3722
rect -44 3664 -2 3720
rect 158 3664 200 3720
rect -44 3598 200 3664
rect -44 3596 0 3598
rect 156 3596 200 3598
rect -44 3540 -2 3596
rect 158 3540 200 3596
rect -44 3474 200 3540
rect -44 3472 0 3474
rect 156 3472 200 3474
rect -44 3416 -2 3472
rect 158 3416 200 3472
rect -44 3350 200 3416
rect -44 3348 0 3350
rect 156 3348 200 3350
rect -44 3292 -2 3348
rect 158 3292 200 3348
rect -44 3226 200 3292
rect -44 3224 0 3226
rect 156 3224 200 3226
rect -44 3168 -2 3224
rect 158 3168 200 3224
rect -44 3102 200 3168
rect -44 3100 0 3102
rect 156 3100 200 3102
rect -44 3044 -2 3100
rect 158 3044 200 3100
rect -44 2978 200 3044
rect -44 2976 0 2978
rect 156 2976 200 2978
rect -44 2920 -2 2976
rect 158 2920 200 2976
rect -44 2854 200 2920
rect -44 2852 0 2854
rect 156 2852 200 2854
rect -44 2796 -2 2852
rect 158 2796 200 2852
rect -44 2730 200 2796
rect -44 2728 0 2730
rect 156 2728 200 2730
rect -44 2672 -2 2728
rect 158 2672 200 2728
rect -44 2606 200 2672
rect -44 2604 0 2606
rect 156 2604 200 2606
rect -44 2548 -2 2604
rect 158 2548 200 2604
rect -44 2482 200 2548
rect -44 2430 0 2482
rect 156 2430 200 2482
rect -44 2358 200 2430
rect -44 2306 0 2358
rect 156 2306 200 2358
rect -44 2235 200 2306
rect -44 2179 -2 2235
rect 158 2179 200 2235
rect -44 2111 200 2179
rect -44 2055 -2 2111
rect 158 2055 200 2111
rect -44 1987 200 2055
rect -44 1931 -2 1987
rect 158 1931 200 1987
rect -44 1863 200 1931
rect -44 1807 -2 1863
rect 158 1807 200 1863
rect -44 1739 200 1807
rect -44 1683 -2 1739
rect 158 1683 200 1739
rect -44 1615 200 1683
rect -44 1559 -2 1615
rect 158 1559 200 1615
rect -44 1491 200 1559
rect -44 1435 -2 1491
rect 158 1435 200 1491
rect -44 1367 200 1435
rect -44 1311 -2 1367
rect 158 1311 200 1367
rect -44 1243 200 1311
rect -44 1187 -2 1243
rect 158 1187 200 1243
rect -44 1119 200 1187
rect -44 1063 -2 1119
rect 158 1063 200 1119
rect -44 995 200 1063
rect -44 939 -2 995
rect 158 939 200 995
rect -44 871 200 939
rect -44 815 -2 871
rect 158 815 200 871
rect -44 747 200 815
rect -44 691 -2 747
rect 158 691 200 747
rect -44 623 200 691
rect -44 567 -2 623
rect 158 567 200 623
rect -44 499 200 567
rect -44 443 -2 499
rect 158 443 200 499
rect -44 375 200 443
rect -44 319 -2 375
rect 158 319 200 375
rect -44 251 200 319
rect -44 195 -2 251
rect 158 195 200 251
rect -44 127 200 195
rect -44 71 -2 127
rect 158 71 200 127
rect -44 0 200 71
rect 360 7299 2004 7400
rect 360 7247 412 7299
rect 464 7247 536 7299
rect 588 7247 660 7299
rect 712 7247 784 7299
rect 836 7247 908 7299
rect 960 7247 1032 7299
rect 1084 7247 1156 7299
rect 1208 7247 1280 7299
rect 1332 7247 1404 7299
rect 1456 7247 1528 7299
rect 1580 7247 1652 7299
rect 1704 7247 1776 7299
rect 1828 7247 1900 7299
rect 1952 7247 2004 7299
rect 360 7175 2004 7247
rect 360 7123 412 7175
rect 464 7123 536 7175
rect 588 7123 660 7175
rect 712 7123 784 7175
rect 836 7123 908 7175
rect 960 7123 1032 7175
rect 1084 7123 1156 7175
rect 1208 7123 1280 7175
rect 1332 7123 1404 7175
rect 1456 7123 1528 7175
rect 1580 7123 1652 7175
rect 1704 7123 1776 7175
rect 1828 7123 1900 7175
rect 1952 7123 2004 7175
rect 360 7051 2004 7123
rect 360 6999 412 7051
rect 464 6999 536 7051
rect 588 6999 660 7051
rect 712 6999 784 7051
rect 836 6999 908 7051
rect 960 6999 1032 7051
rect 1084 6999 1156 7051
rect 1208 6999 1280 7051
rect 1332 6999 1404 7051
rect 1456 6999 1528 7051
rect 1580 6999 1652 7051
rect 1704 6999 1776 7051
rect 1828 6999 1900 7051
rect 1952 6999 2004 7051
rect 360 6927 2004 6999
rect 360 6875 412 6927
rect 464 6875 536 6927
rect 588 6875 660 6927
rect 712 6875 784 6927
rect 836 6875 908 6927
rect 960 6875 1032 6927
rect 1084 6875 1156 6927
rect 1208 6875 1280 6927
rect 1332 6875 1404 6927
rect 1456 6875 1528 6927
rect 1580 6875 1652 6927
rect 1704 6875 1776 6927
rect 1828 6875 1900 6927
rect 1952 6875 2004 6927
rect 360 6803 2004 6875
rect 360 6751 412 6803
rect 464 6751 536 6803
rect 588 6751 660 6803
rect 712 6751 784 6803
rect 836 6751 908 6803
rect 960 6751 1032 6803
rect 1084 6751 1156 6803
rect 1208 6751 1280 6803
rect 1332 6751 1404 6803
rect 1456 6751 1528 6803
rect 1580 6751 1652 6803
rect 1704 6751 1776 6803
rect 1828 6751 1900 6803
rect 1952 6751 2004 6803
rect 360 6679 2004 6751
rect 360 6627 412 6679
rect 464 6627 536 6679
rect 588 6627 660 6679
rect 712 6627 784 6679
rect 836 6627 908 6679
rect 960 6627 1032 6679
rect 1084 6627 1156 6679
rect 1208 6627 1280 6679
rect 1332 6627 1404 6679
rect 1456 6627 1528 6679
rect 1580 6627 1652 6679
rect 1704 6627 1776 6679
rect 1828 6627 1900 6679
rect 1952 6627 2004 6679
rect 360 6555 2004 6627
rect 360 6503 412 6555
rect 464 6503 536 6555
rect 588 6503 660 6555
rect 712 6503 784 6555
rect 836 6503 908 6555
rect 960 6503 1032 6555
rect 1084 6503 1156 6555
rect 1208 6503 1280 6555
rect 1332 6503 1404 6555
rect 1456 6503 1528 6555
rect 1580 6503 1652 6555
rect 1704 6503 1776 6555
rect 1828 6503 1900 6555
rect 1952 6503 2004 6555
rect 360 6431 2004 6503
rect 360 6379 412 6431
rect 464 6379 536 6431
rect 588 6379 660 6431
rect 712 6379 784 6431
rect 836 6379 908 6431
rect 960 6379 1032 6431
rect 1084 6379 1156 6431
rect 1208 6379 1280 6431
rect 1332 6379 1404 6431
rect 1456 6379 1528 6431
rect 1580 6379 1652 6431
rect 1704 6379 1776 6431
rect 1828 6379 1900 6431
rect 1952 6379 2004 6431
rect 360 6307 2004 6379
rect 360 6255 412 6307
rect 464 6255 536 6307
rect 588 6255 660 6307
rect 712 6255 784 6307
rect 836 6255 908 6307
rect 960 6255 1032 6307
rect 1084 6255 1156 6307
rect 1208 6255 1280 6307
rect 1332 6255 1404 6307
rect 1456 6255 1528 6307
rect 1580 6255 1652 6307
rect 1704 6255 1776 6307
rect 1828 6255 1900 6307
rect 1952 6255 2004 6307
rect 360 6183 2004 6255
rect 360 6131 412 6183
rect 464 6131 536 6183
rect 588 6131 660 6183
rect 712 6131 784 6183
rect 836 6131 908 6183
rect 960 6131 1032 6183
rect 1084 6131 1156 6183
rect 1208 6131 1280 6183
rect 1332 6131 1404 6183
rect 1456 6131 1528 6183
rect 1580 6131 1652 6183
rect 1704 6131 1776 6183
rect 1828 6131 1900 6183
rect 1952 6131 2004 6183
rect 360 6059 2004 6131
rect 360 6007 412 6059
rect 464 6007 536 6059
rect 588 6007 660 6059
rect 712 6007 784 6059
rect 836 6007 908 6059
rect 960 6007 1032 6059
rect 1084 6007 1156 6059
rect 1208 6007 1280 6059
rect 1332 6007 1404 6059
rect 1456 6007 1528 6059
rect 1580 6007 1652 6059
rect 1704 6007 1776 6059
rect 1828 6007 1900 6059
rect 1952 6007 2004 6059
rect 360 5935 2004 6007
rect 360 5883 412 5935
rect 464 5883 536 5935
rect 588 5883 660 5935
rect 712 5883 784 5935
rect 836 5883 908 5935
rect 960 5883 1032 5935
rect 1084 5883 1156 5935
rect 1208 5883 1280 5935
rect 1332 5883 1404 5935
rect 1456 5883 1528 5935
rect 1580 5883 1652 5935
rect 1704 5883 1776 5935
rect 1828 5883 1900 5935
rect 1952 5883 2004 5935
rect 360 5811 2004 5883
rect 360 5759 412 5811
rect 464 5759 536 5811
rect 588 5759 660 5811
rect 712 5759 784 5811
rect 836 5759 908 5811
rect 960 5759 1032 5811
rect 1084 5759 1156 5811
rect 1208 5759 1280 5811
rect 1332 5759 1404 5811
rect 1456 5759 1528 5811
rect 1580 5759 1652 5811
rect 1704 5759 1776 5811
rect 1828 5759 1900 5811
rect 1952 5759 2004 5811
rect 360 5687 2004 5759
rect 360 5635 412 5687
rect 464 5635 536 5687
rect 588 5635 660 5687
rect 712 5635 784 5687
rect 836 5635 908 5687
rect 960 5635 1032 5687
rect 1084 5635 1156 5687
rect 1208 5635 1280 5687
rect 1332 5635 1404 5687
rect 1456 5635 1528 5687
rect 1580 5635 1652 5687
rect 1704 5635 1776 5687
rect 1828 5635 1900 5687
rect 1952 5635 2004 5687
rect 360 5563 2004 5635
rect 360 5511 412 5563
rect 464 5511 536 5563
rect 588 5511 660 5563
rect 712 5511 784 5563
rect 836 5511 908 5563
rect 960 5511 1032 5563
rect 1084 5511 1156 5563
rect 1208 5511 1280 5563
rect 1332 5511 1404 5563
rect 1456 5511 1528 5563
rect 1580 5511 1652 5563
rect 1704 5511 1776 5563
rect 1828 5511 1900 5563
rect 1952 5511 2004 5563
rect 360 5439 2004 5511
rect 360 5387 412 5439
rect 464 5387 536 5439
rect 588 5387 660 5439
rect 712 5387 784 5439
rect 836 5387 908 5439
rect 960 5387 1032 5439
rect 1084 5387 1156 5439
rect 1208 5387 1280 5439
rect 1332 5387 1404 5439
rect 1456 5387 1528 5439
rect 1580 5387 1652 5439
rect 1704 5387 1776 5439
rect 1828 5387 1900 5439
rect 1952 5387 2004 5439
rect 360 5315 2004 5387
rect 360 5263 412 5315
rect 464 5263 536 5315
rect 588 5263 660 5315
rect 712 5263 784 5315
rect 836 5263 908 5315
rect 960 5263 1032 5315
rect 1084 5263 1156 5315
rect 1208 5263 1280 5315
rect 1332 5263 1404 5315
rect 1456 5263 1528 5315
rect 1580 5263 1652 5315
rect 1704 5263 1776 5315
rect 1828 5263 1900 5315
rect 1952 5263 2004 5315
rect 360 5191 2004 5263
rect 360 5139 412 5191
rect 464 5139 536 5191
rect 588 5139 660 5191
rect 712 5139 784 5191
rect 836 5139 908 5191
rect 960 5139 1032 5191
rect 1084 5139 1156 5191
rect 1208 5139 1280 5191
rect 1332 5139 1404 5191
rect 1456 5139 1528 5191
rect 1580 5139 1652 5191
rect 1704 5139 1776 5191
rect 1828 5139 1900 5191
rect 1952 5139 2004 5191
rect 360 5067 2004 5139
rect 360 5015 412 5067
rect 464 5015 536 5067
rect 588 5015 660 5067
rect 712 5015 784 5067
rect 836 5015 908 5067
rect 960 5015 1032 5067
rect 1084 5015 1156 5067
rect 1208 5015 1280 5067
rect 1332 5015 1404 5067
rect 1456 5015 1528 5067
rect 1580 5015 1652 5067
rect 1704 5015 1776 5067
rect 1828 5015 1900 5067
rect 1952 5015 2004 5067
rect 360 4943 2004 5015
rect 360 4891 412 4943
rect 464 4891 536 4943
rect 588 4891 660 4943
rect 712 4891 784 4943
rect 836 4891 908 4943
rect 960 4891 1032 4943
rect 1084 4891 1156 4943
rect 1208 4891 1280 4943
rect 1332 4891 1404 4943
rect 1456 4891 1528 4943
rect 1580 4891 1652 4943
rect 1704 4891 1776 4943
rect 1828 4891 1900 4943
rect 1952 4891 2004 4943
rect 360 4819 2004 4891
rect 360 4767 412 4819
rect 464 4767 536 4819
rect 588 4767 660 4819
rect 712 4767 784 4819
rect 836 4767 908 4819
rect 960 4767 1032 4819
rect 1084 4767 1156 4819
rect 1208 4767 1280 4819
rect 1332 4767 1404 4819
rect 1456 4767 1528 4819
rect 1580 4767 1652 4819
rect 1704 4767 1776 4819
rect 1828 4767 1900 4819
rect 1952 4767 2004 4819
rect 360 4695 2004 4767
rect 360 4643 412 4695
rect 464 4643 536 4695
rect 588 4643 660 4695
rect 712 4643 784 4695
rect 836 4643 908 4695
rect 960 4643 1032 4695
rect 1084 4643 1156 4695
rect 1208 4643 1280 4695
rect 1332 4643 1404 4695
rect 1456 4643 1528 4695
rect 1580 4643 1652 4695
rect 1704 4643 1776 4695
rect 1828 4643 1900 4695
rect 1952 4643 2004 4695
rect 360 4571 2004 4643
rect 360 4519 412 4571
rect 464 4519 536 4571
rect 588 4519 660 4571
rect 712 4519 784 4571
rect 836 4519 908 4571
rect 960 4519 1032 4571
rect 1084 4519 1156 4571
rect 1208 4519 1280 4571
rect 1332 4519 1404 4571
rect 1456 4519 1528 4571
rect 1580 4519 1652 4571
rect 1704 4519 1776 4571
rect 1828 4519 1900 4571
rect 1952 4519 2004 4571
rect 360 4447 2004 4519
rect 360 4395 412 4447
rect 464 4395 536 4447
rect 588 4395 660 4447
rect 712 4395 784 4447
rect 836 4395 908 4447
rect 960 4395 1032 4447
rect 1084 4395 1156 4447
rect 1208 4395 1280 4447
rect 1332 4395 1404 4447
rect 1456 4395 1528 4447
rect 1580 4395 1652 4447
rect 1704 4395 1776 4447
rect 1828 4395 1900 4447
rect 1952 4395 2004 4447
rect 360 4323 2004 4395
rect 360 4271 412 4323
rect 464 4271 536 4323
rect 588 4271 660 4323
rect 712 4271 784 4323
rect 836 4271 908 4323
rect 960 4271 1032 4323
rect 1084 4271 1156 4323
rect 1208 4271 1280 4323
rect 1332 4271 1404 4323
rect 1456 4271 1528 4323
rect 1580 4271 1652 4323
rect 1704 4271 1776 4323
rect 1828 4271 1900 4323
rect 1952 4271 2004 4323
rect 360 4199 2004 4271
rect 360 4147 412 4199
rect 464 4147 536 4199
rect 588 4147 660 4199
rect 712 4147 784 4199
rect 836 4147 908 4199
rect 960 4147 1032 4199
rect 1084 4147 1156 4199
rect 1208 4147 1280 4199
rect 1332 4147 1404 4199
rect 1456 4147 1528 4199
rect 1580 4147 1652 4199
rect 1704 4147 1776 4199
rect 1828 4147 1900 4199
rect 1952 4147 2004 4199
rect 360 4075 2004 4147
rect 360 4023 412 4075
rect 464 4023 536 4075
rect 588 4023 660 4075
rect 712 4023 784 4075
rect 836 4023 908 4075
rect 960 4023 1032 4075
rect 1084 4023 1156 4075
rect 1208 4023 1280 4075
rect 1332 4023 1404 4075
rect 1456 4023 1528 4075
rect 1580 4023 1652 4075
rect 1704 4023 1776 4075
rect 1828 4023 1900 4075
rect 1952 4023 2004 4075
rect 360 3951 2004 4023
rect 360 3899 412 3951
rect 464 3899 536 3951
rect 588 3899 660 3951
rect 712 3899 784 3951
rect 836 3899 908 3951
rect 960 3899 1032 3951
rect 1084 3899 1156 3951
rect 1208 3899 1280 3951
rect 1332 3899 1404 3951
rect 1456 3899 1528 3951
rect 1580 3899 1652 3951
rect 1704 3899 1776 3951
rect 1828 3899 1900 3951
rect 1952 3899 2004 3951
rect 360 3827 2004 3899
rect 360 3775 412 3827
rect 464 3775 536 3827
rect 588 3775 660 3827
rect 712 3775 784 3827
rect 836 3775 908 3827
rect 960 3775 1032 3827
rect 1084 3775 1156 3827
rect 1208 3775 1280 3827
rect 1332 3775 1404 3827
rect 1456 3775 1528 3827
rect 1580 3775 1652 3827
rect 1704 3775 1776 3827
rect 1828 3775 1900 3827
rect 1952 3775 2004 3827
rect 360 3703 2004 3775
rect 360 3651 412 3703
rect 464 3651 536 3703
rect 588 3651 660 3703
rect 712 3651 784 3703
rect 836 3651 908 3703
rect 960 3651 1032 3703
rect 1084 3651 1156 3703
rect 1208 3651 1280 3703
rect 1332 3651 1404 3703
rect 1456 3651 1528 3703
rect 1580 3651 1652 3703
rect 1704 3651 1776 3703
rect 1828 3651 1900 3703
rect 1952 3651 2004 3703
rect 360 3579 2004 3651
rect 360 3527 412 3579
rect 464 3527 536 3579
rect 588 3527 660 3579
rect 712 3527 784 3579
rect 836 3527 908 3579
rect 960 3527 1032 3579
rect 1084 3527 1156 3579
rect 1208 3527 1280 3579
rect 1332 3527 1404 3579
rect 1456 3527 1528 3579
rect 1580 3527 1652 3579
rect 1704 3527 1776 3579
rect 1828 3527 1900 3579
rect 1952 3527 2004 3579
rect 360 3455 2004 3527
rect 360 3403 412 3455
rect 464 3403 536 3455
rect 588 3403 660 3455
rect 712 3403 784 3455
rect 836 3403 908 3455
rect 960 3403 1032 3455
rect 1084 3403 1156 3455
rect 1208 3403 1280 3455
rect 1332 3403 1404 3455
rect 1456 3403 1528 3455
rect 1580 3403 1652 3455
rect 1704 3403 1776 3455
rect 1828 3403 1900 3455
rect 1952 3403 2004 3455
rect 360 3331 2004 3403
rect 360 3279 412 3331
rect 464 3279 536 3331
rect 588 3279 660 3331
rect 712 3279 784 3331
rect 836 3279 908 3331
rect 960 3279 1032 3331
rect 1084 3279 1156 3331
rect 1208 3279 1280 3331
rect 1332 3279 1404 3331
rect 1456 3279 1528 3331
rect 1580 3279 1652 3331
rect 1704 3279 1776 3331
rect 1828 3279 1900 3331
rect 1952 3279 2004 3331
rect 360 3207 2004 3279
rect 360 3155 412 3207
rect 464 3155 536 3207
rect 588 3155 660 3207
rect 712 3155 784 3207
rect 836 3155 908 3207
rect 960 3155 1032 3207
rect 1084 3155 1156 3207
rect 1208 3155 1280 3207
rect 1332 3155 1404 3207
rect 1456 3155 1528 3207
rect 1580 3155 1652 3207
rect 1704 3155 1776 3207
rect 1828 3155 1900 3207
rect 1952 3155 2004 3207
rect 360 3083 2004 3155
rect 360 3031 412 3083
rect 464 3031 536 3083
rect 588 3031 660 3083
rect 712 3031 784 3083
rect 836 3031 908 3083
rect 960 3031 1032 3083
rect 1084 3031 1156 3083
rect 1208 3031 1280 3083
rect 1332 3031 1404 3083
rect 1456 3031 1528 3083
rect 1580 3031 1652 3083
rect 1704 3031 1776 3083
rect 1828 3031 1900 3083
rect 1952 3031 2004 3083
rect 360 2959 2004 3031
rect 360 2907 412 2959
rect 464 2907 536 2959
rect 588 2907 660 2959
rect 712 2907 784 2959
rect 836 2907 908 2959
rect 960 2907 1032 2959
rect 1084 2907 1156 2959
rect 1208 2907 1280 2959
rect 1332 2907 1404 2959
rect 1456 2907 1528 2959
rect 1580 2907 1652 2959
rect 1704 2907 1776 2959
rect 1828 2907 1900 2959
rect 1952 2907 2004 2959
rect 360 2835 2004 2907
rect 360 2783 412 2835
rect 464 2783 536 2835
rect 588 2783 660 2835
rect 712 2783 784 2835
rect 836 2783 908 2835
rect 960 2783 1032 2835
rect 1084 2783 1156 2835
rect 1208 2783 1280 2835
rect 1332 2783 1404 2835
rect 1456 2783 1528 2835
rect 1580 2783 1652 2835
rect 1704 2783 1776 2835
rect 1828 2783 1900 2835
rect 1952 2783 2004 2835
rect 360 2711 2004 2783
rect 360 2659 412 2711
rect 464 2659 536 2711
rect 588 2659 660 2711
rect 712 2659 784 2711
rect 836 2659 908 2711
rect 960 2659 1032 2711
rect 1084 2659 1156 2711
rect 1208 2659 1280 2711
rect 1332 2659 1404 2711
rect 1456 2659 1528 2711
rect 1580 2659 1652 2711
rect 1704 2659 1776 2711
rect 1828 2659 1900 2711
rect 1952 2659 2004 2711
rect 360 2587 2004 2659
rect 360 2535 412 2587
rect 464 2535 536 2587
rect 588 2535 660 2587
rect 712 2535 784 2587
rect 836 2535 908 2587
rect 960 2535 1032 2587
rect 1084 2535 1156 2587
rect 1208 2535 1280 2587
rect 1332 2535 1404 2587
rect 1456 2535 1528 2587
rect 1580 2535 1652 2587
rect 1704 2535 1776 2587
rect 1828 2535 1900 2587
rect 1952 2535 2004 2587
rect 360 2463 2004 2535
rect 360 2411 412 2463
rect 464 2411 536 2463
rect 588 2411 660 2463
rect 712 2411 784 2463
rect 836 2411 908 2463
rect 960 2411 1032 2463
rect 1084 2411 1156 2463
rect 1208 2411 1280 2463
rect 1332 2411 1404 2463
rect 1456 2411 1528 2463
rect 1580 2411 1652 2463
rect 1704 2411 1776 2463
rect 1828 2411 1900 2463
rect 1952 2411 2004 2463
rect 360 2339 2004 2411
rect 360 2287 412 2339
rect 464 2287 536 2339
rect 588 2287 660 2339
rect 712 2287 784 2339
rect 836 2287 908 2339
rect 960 2287 1032 2339
rect 1084 2287 1156 2339
rect 1208 2287 1280 2339
rect 1332 2287 1404 2339
rect 1456 2287 1528 2339
rect 1580 2287 1652 2339
rect 1704 2287 1776 2339
rect 1828 2287 1900 2339
rect 1952 2287 2004 2339
rect 360 2215 2004 2287
rect 360 2163 412 2215
rect 464 2163 536 2215
rect 588 2163 660 2215
rect 712 2163 784 2215
rect 836 2163 908 2215
rect 960 2163 1032 2215
rect 1084 2163 1156 2215
rect 1208 2163 1280 2215
rect 1332 2163 1404 2215
rect 1456 2163 1528 2215
rect 1580 2163 1652 2215
rect 1704 2163 1776 2215
rect 1828 2163 1900 2215
rect 1952 2163 2004 2215
rect 360 2091 2004 2163
rect 360 2039 412 2091
rect 464 2039 536 2091
rect 588 2039 660 2091
rect 712 2039 784 2091
rect 836 2039 908 2091
rect 960 2039 1032 2091
rect 1084 2039 1156 2091
rect 1208 2039 1280 2091
rect 1332 2039 1404 2091
rect 1456 2039 1528 2091
rect 1580 2039 1652 2091
rect 1704 2039 1776 2091
rect 1828 2039 1900 2091
rect 1952 2039 2004 2091
rect 360 1967 2004 2039
rect 360 1915 412 1967
rect 464 1915 536 1967
rect 588 1915 660 1967
rect 712 1915 784 1967
rect 836 1915 908 1967
rect 960 1915 1032 1967
rect 1084 1915 1156 1967
rect 1208 1915 1280 1967
rect 1332 1915 1404 1967
rect 1456 1915 1528 1967
rect 1580 1915 1652 1967
rect 1704 1915 1776 1967
rect 1828 1915 1900 1967
rect 1952 1915 2004 1967
rect 360 1843 2004 1915
rect 360 1791 412 1843
rect 464 1791 536 1843
rect 588 1791 660 1843
rect 712 1791 784 1843
rect 836 1791 908 1843
rect 960 1791 1032 1843
rect 1084 1791 1156 1843
rect 1208 1791 1280 1843
rect 1332 1791 1404 1843
rect 1456 1791 1528 1843
rect 1580 1791 1652 1843
rect 1704 1791 1776 1843
rect 1828 1791 1900 1843
rect 1952 1791 2004 1843
rect 360 1719 2004 1791
rect 360 1667 412 1719
rect 464 1667 536 1719
rect 588 1667 660 1719
rect 712 1667 784 1719
rect 836 1667 908 1719
rect 960 1667 1032 1719
rect 1084 1667 1156 1719
rect 1208 1667 1280 1719
rect 1332 1667 1404 1719
rect 1456 1667 1528 1719
rect 1580 1667 1652 1719
rect 1704 1667 1776 1719
rect 1828 1667 1900 1719
rect 1952 1667 2004 1719
rect 360 1595 2004 1667
rect 360 1543 412 1595
rect 464 1543 536 1595
rect 588 1543 660 1595
rect 712 1543 784 1595
rect 836 1543 908 1595
rect 960 1543 1032 1595
rect 1084 1543 1156 1595
rect 1208 1543 1280 1595
rect 1332 1543 1404 1595
rect 1456 1543 1528 1595
rect 1580 1543 1652 1595
rect 1704 1543 1776 1595
rect 1828 1543 1900 1595
rect 1952 1543 2004 1595
rect 360 1471 2004 1543
rect 360 1419 412 1471
rect 464 1419 536 1471
rect 588 1419 660 1471
rect 712 1419 784 1471
rect 836 1419 908 1471
rect 960 1419 1032 1471
rect 1084 1419 1156 1471
rect 1208 1419 1280 1471
rect 1332 1419 1404 1471
rect 1456 1419 1528 1471
rect 1580 1419 1652 1471
rect 1704 1419 1776 1471
rect 1828 1419 1900 1471
rect 1952 1419 2004 1471
rect 360 1347 2004 1419
rect 360 1295 412 1347
rect 464 1295 536 1347
rect 588 1295 660 1347
rect 712 1295 784 1347
rect 836 1295 908 1347
rect 960 1295 1032 1347
rect 1084 1295 1156 1347
rect 1208 1295 1280 1347
rect 1332 1295 1404 1347
rect 1456 1295 1528 1347
rect 1580 1295 1652 1347
rect 1704 1295 1776 1347
rect 1828 1295 1900 1347
rect 1952 1295 2004 1347
rect 360 1223 2004 1295
rect 360 1171 412 1223
rect 464 1171 536 1223
rect 588 1171 660 1223
rect 712 1171 784 1223
rect 836 1171 908 1223
rect 960 1171 1032 1223
rect 1084 1171 1156 1223
rect 1208 1171 1280 1223
rect 1332 1171 1404 1223
rect 1456 1171 1528 1223
rect 1580 1171 1652 1223
rect 1704 1171 1776 1223
rect 1828 1171 1900 1223
rect 1952 1171 2004 1223
rect 360 1099 2004 1171
rect 360 1047 412 1099
rect 464 1047 536 1099
rect 588 1047 660 1099
rect 712 1047 784 1099
rect 836 1047 908 1099
rect 960 1047 1032 1099
rect 1084 1047 1156 1099
rect 1208 1047 1280 1099
rect 1332 1047 1404 1099
rect 1456 1047 1528 1099
rect 1580 1047 1652 1099
rect 1704 1047 1776 1099
rect 1828 1047 1900 1099
rect 1952 1047 2004 1099
rect 360 975 2004 1047
rect 360 923 412 975
rect 464 923 536 975
rect 588 923 660 975
rect 712 923 784 975
rect 836 923 908 975
rect 960 923 1032 975
rect 1084 923 1156 975
rect 1208 923 1280 975
rect 1332 923 1404 975
rect 1456 923 1528 975
rect 1580 923 1652 975
rect 1704 923 1776 975
rect 1828 923 1900 975
rect 1952 923 2004 975
rect 360 851 2004 923
rect 360 799 412 851
rect 464 799 536 851
rect 588 799 660 851
rect 712 799 784 851
rect 836 799 908 851
rect 960 799 1032 851
rect 1084 799 1156 851
rect 1208 799 1280 851
rect 1332 799 1404 851
rect 1456 799 1528 851
rect 1580 799 1652 851
rect 1704 799 1776 851
rect 1828 799 1900 851
rect 1952 799 2004 851
rect 360 727 2004 799
rect 360 675 412 727
rect 464 675 536 727
rect 588 675 660 727
rect 712 675 784 727
rect 836 675 908 727
rect 960 675 1032 727
rect 1084 675 1156 727
rect 1208 675 1280 727
rect 1332 675 1404 727
rect 1456 675 1528 727
rect 1580 675 1652 727
rect 1704 675 1776 727
rect 1828 675 1900 727
rect 1952 675 2004 727
rect 360 603 2004 675
rect 360 551 412 603
rect 464 551 536 603
rect 588 551 660 603
rect 712 551 784 603
rect 836 551 908 603
rect 960 551 1032 603
rect 1084 551 1156 603
rect 1208 551 1280 603
rect 1332 551 1404 603
rect 1456 551 1528 603
rect 1580 551 1652 603
rect 1704 551 1776 603
rect 1828 551 1900 603
rect 1952 551 2004 603
rect 360 479 2004 551
rect 360 427 412 479
rect 464 427 536 479
rect 588 427 660 479
rect 712 427 784 479
rect 836 427 908 479
rect 960 427 1032 479
rect 1084 427 1156 479
rect 1208 427 1280 479
rect 1332 427 1404 479
rect 1456 427 1528 479
rect 1580 427 1652 479
rect 1704 427 1776 479
rect 1828 427 1900 479
rect 1952 427 2004 479
rect 360 355 2004 427
rect 360 303 412 355
rect 464 303 536 355
rect 588 303 660 355
rect 712 303 784 355
rect 836 303 908 355
rect 960 303 1032 355
rect 1084 303 1156 355
rect 1208 303 1280 355
rect 1332 303 1404 355
rect 1456 303 1528 355
rect 1580 303 1652 355
rect 1704 303 1776 355
rect 1828 303 1900 355
rect 1952 303 2004 355
rect 360 231 2004 303
rect 360 179 412 231
rect 464 179 536 231
rect 588 179 660 231
rect 712 179 784 231
rect 836 179 908 231
rect 960 179 1032 231
rect 1084 179 1156 231
rect 1208 179 1280 231
rect 1332 179 1404 231
rect 1456 179 1528 231
rect 1580 179 1652 231
rect 1704 179 1776 231
rect 1828 179 1900 231
rect 1952 179 2004 231
rect 360 107 2004 179
rect 360 55 412 107
rect 464 55 536 107
rect 588 55 660 107
rect 712 55 784 107
rect 836 55 908 107
rect 960 55 1032 107
rect 1084 55 1156 107
rect 1208 55 1280 107
rect 1332 55 1404 107
rect 1456 55 1528 107
rect 1580 55 1652 107
rect 1704 55 1776 107
rect 1828 55 1900 107
rect 1952 55 2004 107
rect 360 0 2004 55
<< via2 >>
rect -2 7266 0 7307
rect 0 7266 156 7307
rect 156 7266 158 7307
rect -2 7251 158 7266
rect -2 7142 0 7183
rect 0 7142 156 7183
rect 156 7142 158 7183
rect -2 7127 158 7142
rect -2 7018 0 7059
rect 0 7018 156 7059
rect 156 7018 158 7059
rect -2 7003 158 7018
rect -2 6894 0 6935
rect 0 6894 156 6935
rect 156 6894 158 6935
rect -2 6879 158 6894
rect -2 6770 0 6811
rect 0 6770 156 6811
rect 156 6770 158 6811
rect -2 6755 158 6770
rect -2 6646 0 6687
rect 0 6646 156 6687
rect 156 6646 158 6687
rect -2 6631 158 6646
rect -2 6522 0 6563
rect 0 6522 156 6563
rect 156 6522 158 6563
rect -2 6507 158 6522
rect -2 6398 0 6439
rect 0 6398 156 6439
rect 156 6398 158 6439
rect -2 6383 158 6398
rect -2 6274 0 6315
rect 0 6274 156 6315
rect 156 6274 158 6315
rect -2 6259 158 6274
rect -2 6150 0 6191
rect 0 6150 156 6191
rect 156 6150 158 6191
rect -2 6135 158 6150
rect -2 6026 0 6067
rect 0 6026 156 6067
rect 156 6026 158 6067
rect -2 6011 158 6026
rect -2 5902 0 5943
rect 0 5902 156 5943
rect 156 5902 158 5943
rect -2 5887 158 5902
rect -2 5778 0 5819
rect 0 5778 156 5819
rect 156 5778 158 5819
rect -2 5763 158 5778
rect -2 5406 0 5456
rect 0 5406 156 5456
rect 156 5406 158 5456
rect -2 5400 158 5406
rect -2 5282 0 5332
rect 0 5282 156 5332
rect 156 5282 158 5332
rect -2 5276 158 5282
rect -2 5158 0 5208
rect 0 5158 156 5208
rect 156 5158 158 5208
rect -2 5152 158 5158
rect -2 5034 0 5084
rect 0 5034 156 5084
rect 156 5034 158 5084
rect -2 5028 158 5034
rect -2 4910 0 4960
rect 0 4910 156 4960
rect 156 4910 158 4960
rect -2 4904 158 4910
rect -2 4786 0 4836
rect 0 4786 156 4836
rect 156 4786 158 4836
rect -2 4780 158 4786
rect -2 4662 0 4712
rect 0 4662 156 4712
rect 156 4662 158 4712
rect -2 4656 158 4662
rect -2 4538 0 4588
rect 0 4538 156 4588
rect 156 4538 158 4588
rect -2 4532 158 4538
rect -2 4414 0 4464
rect 0 4414 156 4464
rect 156 4414 158 4464
rect -2 4408 158 4414
rect -2 4290 0 4340
rect 0 4290 156 4340
rect 156 4290 158 4340
rect -2 4284 158 4290
rect -2 4166 0 4216
rect 0 4166 156 4216
rect 156 4166 158 4216
rect -2 4160 158 4166
rect -2 4042 0 4092
rect 0 4042 156 4092
rect 156 4042 158 4092
rect -2 4036 158 4042
rect -2 3918 0 3968
rect 0 3918 156 3968
rect 156 3918 158 3968
rect -2 3912 158 3918
rect -2 3794 0 3844
rect 0 3794 156 3844
rect 156 3794 158 3844
rect -2 3788 158 3794
rect -2 3670 0 3720
rect 0 3670 156 3720
rect 156 3670 158 3720
rect -2 3664 158 3670
rect -2 3546 0 3596
rect 0 3546 156 3596
rect 156 3546 158 3596
rect -2 3540 158 3546
rect -2 3422 0 3472
rect 0 3422 156 3472
rect 156 3422 158 3472
rect -2 3416 158 3422
rect -2 3298 0 3348
rect 0 3298 156 3348
rect 156 3298 158 3348
rect -2 3292 158 3298
rect -2 3174 0 3224
rect 0 3174 156 3224
rect 156 3174 158 3224
rect -2 3168 158 3174
rect -2 3050 0 3100
rect 0 3050 156 3100
rect 156 3050 158 3100
rect -2 3044 158 3050
rect -2 2926 0 2976
rect 0 2926 156 2976
rect 156 2926 158 2976
rect -2 2920 158 2926
rect -2 2802 0 2852
rect 0 2802 156 2852
rect 156 2802 158 2852
rect -2 2796 158 2802
rect -2 2678 0 2728
rect 0 2678 156 2728
rect 156 2678 158 2728
rect -2 2672 158 2678
rect -2 2554 0 2604
rect 0 2554 156 2604
rect 156 2554 158 2604
rect -2 2548 158 2554
rect -2 2234 158 2235
rect -2 2182 0 2234
rect 0 2182 156 2234
rect 156 2182 158 2234
rect -2 2179 158 2182
rect -2 2110 158 2111
rect -2 2058 0 2110
rect 0 2058 156 2110
rect 156 2058 158 2110
rect -2 2055 158 2058
rect -2 1986 158 1987
rect -2 1934 0 1986
rect 0 1934 156 1986
rect 156 1934 158 1986
rect -2 1931 158 1934
rect -2 1862 158 1863
rect -2 1810 0 1862
rect 0 1810 156 1862
rect 156 1810 158 1862
rect -2 1807 158 1810
rect -2 1738 158 1739
rect -2 1686 0 1738
rect 0 1686 156 1738
rect 156 1686 158 1738
rect -2 1683 158 1686
rect -2 1614 158 1615
rect -2 1562 0 1614
rect 0 1562 156 1614
rect 156 1562 158 1614
rect -2 1559 158 1562
rect -2 1490 158 1491
rect -2 1438 0 1490
rect 0 1438 156 1490
rect 156 1438 158 1490
rect -2 1435 158 1438
rect -2 1366 158 1367
rect -2 1314 0 1366
rect 0 1314 156 1366
rect 156 1314 158 1366
rect -2 1311 158 1314
rect -2 1242 158 1243
rect -2 1190 0 1242
rect 0 1190 156 1242
rect 156 1190 158 1242
rect -2 1187 158 1190
rect -2 1118 158 1119
rect -2 1066 0 1118
rect 0 1066 156 1118
rect 156 1066 158 1118
rect -2 1063 158 1066
rect -2 994 158 995
rect -2 942 0 994
rect 0 942 156 994
rect 156 942 158 994
rect -2 939 158 942
rect -2 870 158 871
rect -2 818 0 870
rect 0 818 156 870
rect 156 818 158 870
rect -2 815 158 818
rect -2 746 158 747
rect -2 694 0 746
rect 0 694 156 746
rect 156 694 158 746
rect -2 691 158 694
rect -2 622 158 623
rect -2 570 0 622
rect 0 570 156 622
rect 156 570 158 622
rect -2 567 158 570
rect -2 498 158 499
rect -2 446 0 498
rect 0 446 156 498
rect 156 446 158 498
rect -2 443 158 446
rect -2 374 158 375
rect -2 322 0 374
rect 0 322 156 374
rect 156 322 158 374
rect -2 319 158 322
rect -2 250 158 251
rect -2 198 0 250
rect 0 198 156 250
rect 156 198 158 250
rect -2 195 158 198
rect -2 126 158 127
rect -2 74 0 126
rect 0 74 156 126
rect 156 74 158 126
rect -2 71 158 74
<< metal3 >>
rect -12 7307 168 7317
rect -12 7251 -2 7307
rect 158 7251 168 7307
rect -12 7183 168 7251
rect -12 7127 -2 7183
rect 158 7127 168 7183
rect -12 7059 168 7127
rect -12 7003 -2 7059
rect 158 7003 168 7059
rect -12 6935 168 7003
rect -12 6879 -2 6935
rect 158 6879 168 6935
rect -12 6811 168 6879
rect -12 6755 -2 6811
rect 158 6755 168 6811
rect -12 6687 168 6755
rect -12 6631 -2 6687
rect 158 6631 168 6687
rect -12 6563 168 6631
rect -12 6507 -2 6563
rect 158 6507 168 6563
rect -12 6439 168 6507
rect -12 6383 -2 6439
rect 158 6383 168 6439
rect -12 6315 168 6383
rect -12 6259 -2 6315
rect 158 6259 168 6315
rect -12 6191 168 6259
rect -12 6135 -2 6191
rect 158 6135 168 6191
rect -12 6067 168 6135
rect -12 6011 -2 6067
rect 158 6011 168 6067
rect -12 5943 168 6011
rect -12 5887 -2 5943
rect 158 5887 168 5943
rect -12 5819 168 5887
rect -12 5763 -2 5819
rect 158 5763 168 5819
rect -12 5753 168 5763
rect -12 5456 168 5466
rect -12 5400 -2 5456
rect 158 5400 168 5456
rect -12 5332 168 5400
rect -12 5276 -2 5332
rect 158 5276 168 5332
rect -12 5208 168 5276
rect -12 5152 -2 5208
rect 158 5152 168 5208
rect -12 5084 168 5152
rect -12 5028 -2 5084
rect 158 5028 168 5084
rect -12 4960 168 5028
rect -12 4904 -2 4960
rect 158 4904 168 4960
rect -12 4836 168 4904
rect -12 4780 -2 4836
rect 158 4780 168 4836
rect -12 4712 168 4780
rect -12 4656 -2 4712
rect 158 4656 168 4712
rect -12 4588 168 4656
rect -12 4532 -2 4588
rect 158 4532 168 4588
rect -12 4464 168 4532
rect -12 4408 -2 4464
rect 158 4408 168 4464
rect -12 4340 168 4408
rect -12 4284 -2 4340
rect 158 4284 168 4340
rect -12 4216 168 4284
rect -12 4160 -2 4216
rect 158 4160 168 4216
rect -12 4092 168 4160
rect -12 4036 -2 4092
rect 158 4036 168 4092
rect -12 3968 168 4036
rect -12 3912 -2 3968
rect 158 3912 168 3968
rect -12 3844 168 3912
rect -12 3788 -2 3844
rect 158 3788 168 3844
rect -12 3720 168 3788
rect -12 3664 -2 3720
rect 158 3664 168 3720
rect -12 3596 168 3664
rect -12 3540 -2 3596
rect 158 3540 168 3596
rect -12 3472 168 3540
rect -12 3416 -2 3472
rect 158 3416 168 3472
rect -12 3348 168 3416
rect -12 3292 -2 3348
rect 158 3292 168 3348
rect -12 3224 168 3292
rect -12 3168 -2 3224
rect 158 3168 168 3224
rect -12 3100 168 3168
rect -12 3044 -2 3100
rect 158 3044 168 3100
rect -12 2976 168 3044
rect -12 2920 -2 2976
rect 158 2920 168 2976
rect -12 2852 168 2920
rect -12 2796 -2 2852
rect 158 2796 168 2852
rect -12 2728 168 2796
rect -12 2672 -2 2728
rect 158 2672 168 2728
rect -12 2604 168 2672
rect -12 2548 -2 2604
rect 158 2548 168 2604
rect -12 2538 168 2548
rect -12 2235 168 2245
rect -12 2179 -2 2235
rect 158 2179 168 2235
rect -12 2111 168 2179
rect -12 2055 -2 2111
rect 158 2055 168 2111
rect -12 1987 168 2055
rect -12 1931 -2 1987
rect 158 1931 168 1987
rect -12 1863 168 1931
rect -12 1807 -2 1863
rect 158 1807 168 1863
rect -12 1739 168 1807
rect -12 1683 -2 1739
rect 158 1683 168 1739
rect -12 1615 168 1683
rect -12 1559 -2 1615
rect 158 1559 168 1615
rect -12 1491 168 1559
rect -12 1435 -2 1491
rect 158 1435 168 1491
rect -12 1367 168 1435
rect -12 1311 -2 1367
rect 158 1311 168 1367
rect -12 1243 168 1311
rect -12 1187 -2 1243
rect 158 1187 168 1243
rect -12 1119 168 1187
rect -12 1063 -2 1119
rect 158 1063 168 1119
rect -12 995 168 1063
rect -12 939 -2 995
rect 158 939 168 995
rect -12 871 168 939
rect -12 815 -2 871
rect 158 815 168 871
rect -12 747 168 815
rect -12 691 -2 747
rect 158 691 168 747
rect -12 623 168 691
rect -12 567 -2 623
rect 158 567 168 623
rect -12 499 168 567
rect -12 443 -2 499
rect 158 443 168 499
rect -12 375 168 443
rect -12 319 -2 375
rect 158 319 168 375
rect -12 251 168 319
rect -12 195 -2 251
rect 158 195 168 251
rect -12 127 168 195
rect -12 71 -2 127
rect 158 71 168 127
rect -12 61 168 71
use M2_M1_CDNS_40661953145304  M2_M1_CDNS_40661953145304_0
timestamp 1698431365
transform 1 0 78 0 1 3696
box 0 0 1 1
use M2_M1_CDNS_40661953145307  M2_M1_CDNS_40661953145307_0
timestamp 1698431365
transform 1 0 1182 0 1 3677
box 0 0 1 1
use M3_M2_CDNS_40661953145303  M3_M2_CDNS_40661953145303_0
timestamp 1698431365
transform 1 0 78 0 1 6535
box 0 0 1 1
use M3_M2_CDNS_40661953145305  M3_M2_CDNS_40661953145305_0
timestamp 1698431365
transform 1 0 78 0 1 4002
box 0 0 1 1
use M3_M2_CDNS_40661953145306  M3_M2_CDNS_40661953145306_0
timestamp 1698431365
transform 1 0 78 0 1 1153
box 0 0 1 1
<< properties >>
string GDS_END 2050434
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2049924
<< end >>
