magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 4342 870
rect -86 352 1249 377
rect 2000 352 4342 377
<< pwell >>
rect 1249 352 2000 377
rect -86 -86 4342 352
<< mvnmos >>
rect 124 156 244 228
rect 348 156 468 228
rect 516 156 636 228
rect 740 156 860 228
rect 908 156 1028 228
rect 1168 135 1288 228
rect 1631 139 1751 232
rect 2043 158 2163 230
rect 2267 158 2387 230
rect 2435 158 2555 230
rect 2716 158 2836 230
rect 2940 158 3060 230
rect 3164 158 3284 230
rect 3332 158 3452 230
rect 3644 143 3764 230
rect 4012 69 4132 232
<< mvpmos >>
rect 124 502 224 628
rect 348 502 448 628
rect 496 502 596 628
rect 700 502 800 628
rect 888 502 988 628
rect 1188 502 1288 686
rect 1651 497 1751 660
rect 2032 502 2132 628
rect 2246 502 2346 628
rect 2424 502 2524 628
rect 2716 502 2818 628
rect 2950 502 3050 628
rect 3164 502 3264 628
rect 3312 502 3412 628
rect 3564 487 3664 628
rect 4032 472 4132 715
<< mvndiff >>
rect 1348 244 1424 257
rect 1348 228 1361 244
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 228
rect 636 215 740 228
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 228
rect 1028 215 1168 228
rect 1028 169 1070 215
rect 1116 169 1168 215
rect 1028 156 1168 169
rect 1088 135 1168 156
rect 1288 198 1361 228
rect 1407 198 1424 244
rect 1811 244 1883 257
rect 1811 232 1824 244
rect 1288 135 1424 198
rect 1543 198 1631 232
rect 1543 152 1556 198
rect 1602 152 1631 198
rect 1543 139 1631 152
rect 1751 198 1824 232
rect 1870 198 1883 244
rect 1751 139 1883 198
rect 1955 217 2043 230
rect 1955 171 1968 217
rect 2014 171 2043 217
rect 1955 158 2043 171
rect 2163 217 2267 230
rect 2163 171 2192 217
rect 2238 171 2267 217
rect 2163 158 2267 171
rect 2387 158 2435 230
rect 2555 217 2716 230
rect 2555 171 2607 217
rect 2653 171 2716 217
rect 2555 158 2716 171
rect 2836 217 2940 230
rect 2836 171 2865 217
rect 2911 171 2940 217
rect 2836 158 2940 171
rect 3060 217 3164 230
rect 3060 171 3089 217
rect 3135 171 3164 217
rect 3060 158 3164 171
rect 3284 158 3332 230
rect 3452 158 3644 230
rect 3512 143 3644 158
rect 3764 209 3852 230
rect 3764 163 3793 209
rect 3839 163 3852 209
rect 3764 143 3852 163
rect 3924 180 4012 232
rect 3512 119 3584 143
rect 3512 73 3525 119
rect 3571 73 3584 119
rect 3924 134 3937 180
rect 3983 134 4012 180
rect 3512 60 3584 73
rect 3924 69 4012 134
rect 4132 180 4220 232
rect 4132 134 4161 180
rect 4207 134 4220 180
rect 4132 69 4220 134
<< mvpdiff >>
rect 1048 686 1120 701
rect 1512 716 1586 729
rect 1048 682 1188 686
rect 1048 636 1061 682
rect 1107 636 1188 682
rect 1048 628 1188 636
rect 36 590 124 628
rect 36 544 49 590
rect 95 544 124 590
rect 36 502 124 544
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 502 348 569
rect 448 502 496 628
rect 596 587 700 628
rect 596 541 625 587
rect 671 541 700 587
rect 596 502 700 541
rect 800 502 888 628
rect 988 502 1188 628
rect 1288 561 1376 686
rect 1288 515 1317 561
rect 1363 515 1376 561
rect 1288 502 1376 515
rect 1512 670 1525 716
rect 1571 670 1586 716
rect 1512 660 1586 670
rect 1512 497 1651 660
rect 1751 561 1839 660
rect 2584 645 2656 658
rect 2584 628 2597 645
rect 1751 515 1780 561
rect 1826 515 1839 561
rect 1751 497 1839 515
rect 1944 595 2032 628
rect 1944 549 1957 595
rect 2003 549 2032 595
rect 1944 502 2032 549
rect 2132 563 2246 628
rect 2132 517 2171 563
rect 2217 517 2246 563
rect 2132 502 2246 517
rect 2346 502 2424 628
rect 2524 599 2597 628
rect 2643 628 2656 645
rect 3924 662 4032 715
rect 2643 599 2716 628
rect 2524 502 2716 599
rect 2818 563 2950 628
rect 2818 517 2865 563
rect 2911 517 2950 563
rect 2818 502 2950 517
rect 3050 563 3164 628
rect 3050 517 3089 563
rect 3135 517 3164 563
rect 3050 502 3164 517
rect 3264 502 3312 628
rect 3412 615 3564 628
rect 3412 569 3461 615
rect 3507 569 3564 615
rect 3412 502 3564 569
rect 3472 487 3564 502
rect 3664 579 3752 628
rect 3664 533 3693 579
rect 3739 533 3752 579
rect 3664 487 3752 533
rect 3924 616 3947 662
rect 3993 616 4032 662
rect 3924 557 4032 616
rect 3924 511 3947 557
rect 3993 511 4032 557
rect 3924 472 4032 511
rect 4132 662 4220 715
rect 4132 616 4161 662
rect 4207 616 4220 662
rect 4132 557 4220 616
rect 4132 511 4161 557
rect 4207 511 4220 557
rect 4132 472 4220 511
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1070 169 1116 215
rect 1361 198 1407 244
rect 1556 152 1602 198
rect 1824 198 1870 244
rect 1968 171 2014 217
rect 2192 171 2238 217
rect 2607 171 2653 217
rect 2865 171 2911 217
rect 3089 171 3135 217
rect 3793 163 3839 209
rect 3525 73 3571 119
rect 3937 134 3983 180
rect 4161 134 4207 180
<< mvpdiffc >>
rect 1061 636 1107 682
rect 49 544 95 590
rect 263 569 309 615
rect 625 541 671 587
rect 1317 515 1363 561
rect 1525 670 1571 716
rect 1780 515 1826 561
rect 1957 549 2003 595
rect 2171 517 2217 563
rect 2597 599 2643 645
rect 2865 517 2911 563
rect 3089 517 3135 563
rect 3461 569 3507 615
rect 3693 533 3739 579
rect 3947 616 3993 662
rect 3947 511 3993 557
rect 4161 616 4207 662
rect 4161 511 4207 557
<< polysilicon >>
rect 124 720 800 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 700 628 800 720
rect 888 628 988 692
rect 1188 686 1288 730
rect 1651 720 3050 760
rect 1651 660 1751 720
rect 124 351 224 502
rect 124 305 149 351
rect 195 305 224 351
rect 124 272 224 305
rect 348 351 448 502
rect 348 305 375 351
rect 421 305 448 351
rect 496 403 596 502
rect 700 458 800 502
rect 888 458 988 502
rect 496 357 509 403
rect 555 371 596 403
rect 908 434 988 458
rect 1188 442 1288 502
rect 2032 628 2132 672
rect 2246 628 2346 720
rect 2424 628 2524 672
rect 2716 628 2818 672
rect 2950 628 3050 720
rect 4032 715 4132 759
rect 3164 628 3264 672
rect 3312 628 3412 672
rect 3564 628 3664 672
rect 908 388 926 434
rect 972 388 988 434
rect 555 357 860 371
rect 496 325 860 357
rect 348 272 448 305
rect 124 228 244 272
rect 348 228 468 272
rect 516 228 636 272
rect 740 228 860 325
rect 908 272 988 388
rect 1168 424 1288 442
rect 1651 432 1751 497
rect 1651 427 1674 432
rect 1168 378 1209 424
rect 1255 378 1288 424
rect 908 228 1028 272
rect 1168 228 1288 378
rect 1631 386 1674 427
rect 1720 386 1751 432
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1631 232 1751 386
rect 2032 451 2132 502
rect 2246 458 2346 502
rect 2424 460 2524 502
rect 2032 405 2065 451
rect 2111 405 2132 451
rect 2032 389 2132 405
rect 2424 414 2455 460
rect 2501 442 2524 460
rect 2501 414 2555 442
rect 2032 343 2352 389
rect 2424 386 2555 414
rect 2267 292 2352 343
rect 2043 230 2163 274
rect 2267 230 2387 292
rect 2435 230 2555 386
rect 2716 340 2818 502
rect 2950 442 3050 502
rect 3164 469 3264 502
rect 2950 402 3109 442
rect 3164 423 3192 469
rect 3238 423 3264 469
rect 3312 458 3412 502
rect 3164 410 3264 423
rect 2716 294 2736 340
rect 2782 294 2818 340
rect 3068 362 3109 402
rect 3068 322 3224 362
rect 2716 276 2818 294
rect 2940 309 3016 322
rect 2716 230 2836 276
rect 2940 263 2957 309
rect 3003 274 3016 309
rect 3164 274 3224 322
rect 3332 337 3412 458
rect 3564 389 3664 487
rect 4032 402 4132 472
rect 4032 389 4051 402
rect 3564 343 3577 389
rect 3623 365 3664 389
rect 3623 343 3704 365
rect 3332 309 3452 337
rect 3564 325 3704 343
rect 3003 263 3060 274
rect 2940 230 3060 263
rect 3164 230 3284 274
rect 3332 263 3393 309
rect 3439 263 3452 309
rect 3332 230 3452 263
rect 3644 274 3704 325
rect 4012 356 4051 389
rect 4097 356 4132 402
rect 3644 230 3764 274
rect 4012 232 4132 356
rect 1168 91 1288 135
rect 124 24 636 64
rect 1631 70 1751 139
rect 2043 70 2163 158
rect 2267 114 2387 158
rect 2435 114 2555 158
rect 2716 114 2836 158
rect 2940 107 3060 158
rect 3164 114 3284 158
rect 3332 114 3452 158
rect 1631 24 2163 70
rect 3644 99 3764 143
rect 4012 25 4132 69
<< polycontact >>
rect 149 305 195 351
rect 375 305 421 351
rect 509 357 555 403
rect 926 388 972 434
rect 1209 378 1255 424
rect 1674 386 1720 432
rect 2065 405 2111 451
rect 2455 414 2501 460
rect 3192 423 3238 469
rect 2736 294 2782 340
rect 2957 263 3003 309
rect 3577 343 3623 389
rect 3393 263 3439 309
rect 4051 356 4097 402
<< metal1 >>
rect 0 724 4256 844
rect 252 615 320 724
rect 1050 682 1118 724
rect 1050 636 1061 682
rect 1107 636 1118 682
rect 1514 716 1582 724
rect 1514 670 1525 716
rect 1571 670 1582 716
rect 49 590 95 603
rect 252 569 263 615
rect 309 569 320 615
rect 1175 624 1464 664
rect 1674 624 2003 670
rect 1175 618 1720 624
rect 1175 587 1221 618
rect 49 523 95 544
rect 606 541 625 587
rect 671 541 1221 587
rect 1418 578 1720 618
rect 1957 595 2003 624
rect 1317 561 1363 572
rect 49 477 555 523
rect 1780 561 1826 572
rect 1363 515 1720 532
rect 1317 486 1720 515
rect 49 215 95 477
rect 49 158 95 169
rect 141 351 206 430
rect 141 305 149 351
rect 195 305 206 351
rect 141 119 206 305
rect 365 351 430 430
rect 365 305 375 351
rect 421 305 430 351
rect 509 403 555 477
rect 682 434 1017 443
rect 682 388 926 434
rect 972 388 1017 434
rect 682 359 1017 388
rect 1093 424 1326 440
rect 1093 378 1209 424
rect 1255 378 1326 424
rect 1093 359 1326 378
rect 509 325 555 357
rect 273 215 319 228
rect 273 60 319 169
rect 365 119 430 305
rect 885 261 1264 307
rect 885 215 931 261
rect 654 169 665 215
rect 711 169 931 215
rect 1059 169 1070 215
rect 1116 169 1127 215
rect 1059 60 1127 169
rect 1218 152 1264 261
rect 1372 255 1418 486
rect 1674 432 1720 486
rect 1674 375 1720 386
rect 1957 538 2003 549
rect 2065 630 2498 678
rect 1780 410 1826 515
rect 2065 451 2111 630
rect 1780 405 2065 410
rect 1780 364 2111 405
rect 2171 563 2217 574
rect 1350 244 1418 255
rect 1350 198 1361 244
rect 1407 198 1418 244
rect 1464 261 1721 307
rect 1464 152 1510 261
rect 1218 106 1510 152
rect 1556 198 1602 209
rect 1556 60 1602 152
rect 1675 152 1721 261
rect 1813 255 1859 364
rect 2171 340 2217 517
rect 2452 553 2498 630
rect 2586 645 2654 724
rect 2586 599 2597 645
rect 2643 599 2654 645
rect 2734 632 3249 678
rect 2734 553 2780 632
rect 2452 506 2780 553
rect 2865 563 2911 574
rect 2865 460 2911 517
rect 2440 414 2455 460
rect 2501 414 2911 460
rect 2171 294 2736 340
rect 2782 294 2793 340
rect 1813 244 1881 255
rect 1813 198 1824 244
rect 1870 198 1881 244
rect 1968 217 2014 228
rect 1968 152 2014 171
rect 2192 217 2238 294
rect 2865 217 2911 414
rect 2957 309 3003 632
rect 2957 252 3003 263
rect 3089 563 3135 574
rect 3089 355 3135 517
rect 3181 469 3249 632
rect 3450 615 3518 724
rect 3450 569 3461 615
rect 3507 569 3518 615
rect 3947 662 3993 724
rect 3693 579 3739 590
rect 3181 423 3192 469
rect 3238 423 3249 469
rect 3181 414 3249 423
rect 3301 463 3634 510
rect 3301 355 3347 463
rect 3089 308 3347 355
rect 3566 389 3634 463
rect 3566 343 3577 389
rect 3623 343 3634 389
rect 3693 402 3739 533
rect 3947 557 3993 616
rect 3947 492 3993 511
rect 4158 662 4230 673
rect 4158 616 4161 662
rect 4207 616 4230 662
rect 4158 557 4230 616
rect 4158 511 4161 557
rect 4207 511 4230 557
rect 3693 356 4051 402
rect 4097 356 4108 402
rect 3566 334 3634 343
rect 3393 309 3439 320
rect 2192 160 2238 171
rect 2596 171 2607 217
rect 2653 171 2664 217
rect 1675 106 2014 152
rect 2596 60 2664 171
rect 2865 160 2911 171
rect 3089 217 3135 308
rect 3393 246 3439 263
rect 3793 246 3839 356
rect 3393 209 3839 246
rect 3393 199 3793 209
rect 3089 160 3135 171
rect 3793 152 3839 163
rect 3937 180 3983 199
rect 3525 119 3571 136
rect 3525 60 3571 73
rect 3937 60 3983 134
rect 4158 180 4230 511
rect 4158 134 4161 180
rect 4207 134 4230 180
rect 4158 123 4230 134
rect 0 -60 4256 60
<< labels >>
flabel metal1 s 4158 123 4230 673 0 FreeSans 400 0 0 0 Q
port 5 nsew default output
flabel metal1 s 141 119 206 430 0 FreeSans 400 0 0 0 SE
port 2 nsew default input
flabel metal1 s 365 119 430 430 0 FreeSans 400 0 0 0 SI
port 3 nsew default input
flabel metal1 s 0 724 4256 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 273 217 319 228 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1093 359 1326 440 0 FreeSans 400 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 682 359 1017 443 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 3947 670 3993 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 670 3518 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 670 2654 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1514 670 1582 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 670 1118 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 636 3993 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 636 3518 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 636 2654 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 636 1118 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 636 320 670 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 599 3993 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 599 3518 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 599 2654 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 599 320 636 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 569 3993 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 569 3518 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 599 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 492 3993 569 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2596 215 2664 217 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 215 319 217 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2596 209 2664 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1059 209 1127 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 209 319 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2596 199 2664 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1556 199 1602 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1059 199 1127 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 199 319 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 136 3983 199 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2596 136 2664 199 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1556 136 1602 199 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1059 136 1127 199 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 136 319 199 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3937 60 3983 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3525 60 3571 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2596 60 2664 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1556 60 1602 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1059 60 1127 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 136 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string GDS_END 191330
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 182370
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
