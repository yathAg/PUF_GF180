magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 352 310 870
<< pwell >>
rect -86 -86 310 352
<< metal1 >>
rect 0 724 224 844
rect 28 162 95 542
rect 0 -60 224 60
<< labels >>
rlabel metal1 s 28 162 95 542 6 I
port 1 nsew default input
rlabel metal1 s 0 724 224 844 6 VDD
port 2 nsew power bidirectional abutment
rlabel nwell s -86 352 310 870 6 VNW
port 3 nsew power bidirectional
rlabel pwell s -86 -86 310 352 6 VPW
port 4 nsew ground bidirectional
rlabel metal1 s 0 -60 224 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 224 784
string LEFclass core ANTENNACELL
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1248338
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1246732
<< end >>
