magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< isosubstrate >>
rect 251 53100 14727 57210
rect 2457 47163 12521 53100
rect 601 42936 14377 47163
rect 957 26552 12844 42936
rect 957 1096 14021 26552
<< nwell >>
rect 2457 52160 12521 52716
rect 2457 48116 3013 52160
rect 11965 48116 12521 52160
rect 2457 47560 12521 48116
<< pwell >>
rect 747 53655 3923 56655
rect 4183 53655 7359 56655
rect 7619 53655 10795 56655
rect 11055 53655 14231 56655
<< mvndiff >>
rect 747 56618 835 56655
rect 747 53692 760 56618
rect 806 53692 835 56618
rect 747 53655 835 53692
rect 3835 56618 3923 56655
rect 3835 53692 3864 56618
rect 3910 53692 3923 56618
rect 3835 53655 3923 53692
rect 4183 56618 4271 56655
rect 4183 53692 4196 56618
rect 4242 53692 4271 56618
rect 4183 53655 4271 53692
rect 7271 56618 7359 56655
rect 7271 53692 7300 56618
rect 7346 53692 7359 56618
rect 7271 53655 7359 53692
rect 7619 56618 7707 56655
rect 7619 53692 7632 56618
rect 7678 53692 7707 56618
rect 7619 53655 7707 53692
rect 10707 56618 10795 56655
rect 10707 53692 10736 56618
rect 10782 53692 10795 56618
rect 10707 53655 10795 53692
rect 11055 56618 11143 56655
rect 11055 53692 11068 56618
rect 11114 53692 11143 56618
rect 11055 53655 11143 53692
rect 14143 56618 14231 56655
rect 14143 53692 14172 56618
rect 14218 53692 14231 56618
rect 14143 53655 14231 53692
<< mvndiffc >>
rect 760 53692 806 56618
rect 3864 53692 3910 56618
rect 4196 53692 4242 56618
rect 7300 53692 7346 56618
rect 7632 53692 7678 56618
rect 10736 53692 10782 56618
rect 11068 53692 11114 56618
rect 14172 53692 14218 56618
<< psubdiff >>
rect 334 57105 14644 57127
rect 334 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57037 14576 57059
rect 402 53273 424 57037
rect 14554 53273 14576 57037
rect 402 53251 14576 53273
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14644 57105
rect 334 53183 14644 53205
rect 246 52611 2236 52633
rect 246 47665 268 52611
rect 2214 47665 2236 52611
rect 246 47643 2236 47665
rect 3094 52029 11884 52051
rect 3094 51983 3142 52029
rect 11836 51983 11884 52029
rect 3094 51900 11884 51983
rect 3094 48376 3116 51900
rect 3162 51875 11816 51900
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51807 11662 51829
rect 3316 51271 3338 51807
rect 11640 51271 11662 51807
rect 3316 51249 11662 51271
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51095 11816 51203
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 50941 11816 51049
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50873 11662 50895
rect 3316 50337 3338 50873
rect 11640 50337 11662 50873
rect 3316 50315 11662 50337
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50161 11816 50269
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50007 11816 50115
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49939 11662 49961
rect 3316 49403 3338 49939
rect 11640 49403 11662 49939
rect 3316 49381 11662 49403
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49227 11816 49335
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49073 11816 49181
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49005 11662 49027
rect 3316 48469 3338 49005
rect 11640 48469 11662 49005
rect 3316 48447 11662 48469
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48376 11816 48401
rect 11862 48376 11884 51900
rect 3094 48293 11884 48376
rect 3094 48247 3142 48293
rect 11836 48247 11884 48293
rect 3094 48225 11884 48247
rect 12742 52611 14732 52633
rect 12742 47665 12764 52611
rect 14710 47665 14732 52611
rect 12742 47643 14732 47665
rect 246 42647 736 42669
rect 246 1201 268 42647
rect 714 1201 736 42647
rect 13001 42647 13991 42669
rect 13001 27201 13023 42647
rect 13969 27201 13991 42647
rect 13001 27179 13991 27201
rect 14242 42647 14732 42669
rect 246 1179 736 1201
rect 14242 1201 14264 42647
rect 14710 1201 14732 42647
rect 14242 1179 14732 1201
<< nsubdiff >>
rect 2540 52611 12438 52633
rect 2540 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52243 12070 52265
rect 2908 48033 2930 52243
rect 12048 48033 12070 52243
rect 2908 48011 12070 48033
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12438 52611
rect 2540 47643 12438 47665
<< psubdiffcont >>
rect 356 53205 402 57105
rect 510 57059 14468 57105
rect 510 53205 14468 53251
rect 14576 53205 14622 57105
rect 268 47665 2214 52611
rect 3142 51983 11836 52029
rect 3116 48376 3162 51900
rect 3270 51234 3316 51844
rect 3424 51829 11554 51875
rect 3424 51203 11554 51249
rect 11662 51234 11708 51844
rect 3330 51049 11648 51095
rect 3270 50300 3316 50910
rect 3424 50895 11554 50941
rect 3424 50269 11554 50315
rect 11662 50300 11708 50910
rect 3330 50115 11648 50161
rect 3270 49366 3316 49976
rect 3424 49961 11554 50007
rect 3424 49335 11554 49381
rect 11662 49366 11708 49976
rect 3330 49181 11648 49227
rect 3270 48432 3316 49042
rect 3424 49027 11554 49073
rect 3424 48401 11554 48447
rect 11662 48432 11708 49042
rect 11816 48376 11862 51900
rect 3142 48247 11836 48293
rect 12764 47665 14710 52611
rect 268 1201 714 42647
rect 13023 27201 13969 42647
rect 14264 1201 14710 42647
<< nsubdiffcont >>
rect 2562 47665 2908 52611
rect 3016 52265 11962 52611
rect 3016 47665 11962 48011
rect 12070 47665 12416 52611
<< mvnmoscap >>
rect 835 53655 3835 56655
rect 4271 53655 7271 56655
rect 7707 53655 10707 56655
rect 11143 53655 14143 56655
<< polysilicon >>
rect 835 56734 3835 56747
rect 835 56688 888 56734
rect 3782 56688 3835 56734
rect 835 56655 3835 56688
rect 4271 56734 7271 56747
rect 4271 56688 4324 56734
rect 7218 56688 7271 56734
rect 4271 56655 7271 56688
rect 7707 56734 10707 56747
rect 7707 56688 7760 56734
rect 10654 56688 10707 56734
rect 7707 56655 10707 56688
rect 11143 56734 14143 56747
rect 11143 56688 11196 56734
rect 14090 56688 14143 56734
rect 11143 56655 14143 56688
rect 835 53622 3835 53655
rect 835 53576 888 53622
rect 3782 53576 3835 53622
rect 835 53563 3835 53576
rect 4271 53622 7271 53655
rect 4271 53576 4324 53622
rect 7218 53576 7271 53622
rect 4271 53563 7271 53576
rect 7707 53622 10707 53655
rect 7707 53576 7760 53622
rect 10654 53576 10707 53622
rect 7707 53563 10707 53576
rect 11143 53622 14143 53655
rect 11143 53576 11196 53622
rect 14090 53576 14143 53622
rect 11143 53563 14143 53576
<< polycontact >>
rect 888 56688 3782 56734
rect 4324 56688 7218 56734
rect 7760 56688 10654 56734
rect 11196 56688 14090 56734
rect 888 53576 3782 53622
rect 4324 53576 7218 53622
rect 7760 53576 10654 53622
rect 11196 53576 14090 53622
<< mvndiode >>
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51498 11489 51580
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50564 11489 50646
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49630 11489 49712
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48696 11489 48778
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
<< mvndiodec >>
rect 3502 51580 11476 51626
rect 3502 51452 11476 51498
rect 3502 50646 11476 50692
rect 3502 50518 11476 50564
rect 3502 49712 11476 49758
rect 3502 49584 11476 49630
rect 3502 48778 11476 48824
rect 3502 48650 11476 48696
<< metal1 >>
rect 2489 57116 2673 57120
rect 4859 57116 5043 57120
rect 7235 57116 7743 57120
rect 9935 57116 10119 57120
rect 12305 57116 12489 57120
rect 345 57108 14633 57116
rect 345 57105 2501 57108
rect 2553 57105 2609 57108
rect 2661 57105 4871 57108
rect 4923 57105 4979 57108
rect 5031 57105 7247 57108
rect 7299 57105 7355 57108
rect 7407 57105 7463 57108
rect 7515 57105 7571 57108
rect 7623 57105 7679 57108
rect 7731 57105 9947 57108
rect 9999 57105 10055 57108
rect 10107 57105 12317 57108
rect 12369 57105 12425 57108
rect 12477 57105 14633 57108
rect 345 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57056 2501 57059
rect 2553 57056 2609 57059
rect 2661 57056 4871 57059
rect 4923 57056 4979 57059
rect 5031 57056 7247 57059
rect 7299 57056 7355 57059
rect 7407 57056 7463 57059
rect 7515 57056 7571 57059
rect 7623 57056 7679 57059
rect 7731 57056 9947 57059
rect 9999 57056 10055 57059
rect 10107 57056 12317 57059
rect 12369 57056 12425 57059
rect 12477 57056 14576 57059
rect 402 57048 14576 57056
rect 402 56655 413 57048
rect 2489 57044 2673 57048
rect 4859 57044 5043 57048
rect 7235 57044 7743 57048
rect 9935 57044 10119 57048
rect 12305 57044 12489 57048
rect 877 56734 3793 56745
rect 877 56688 888 56734
rect 3782 56688 3793 56734
rect 877 56677 3793 56688
rect 877 56669 1877 56677
rect 402 56618 817 56655
rect 402 53692 760 56618
rect 806 53692 817 56618
rect 402 53505 817 53692
rect 877 56617 917 56669
rect 969 56617 1041 56669
rect 1093 56617 1165 56669
rect 1217 56617 1289 56669
rect 1341 56617 1413 56669
rect 1465 56617 1537 56669
rect 1589 56617 1661 56669
rect 1713 56617 1785 56669
rect 1837 56617 1877 56669
rect 877 56545 1877 56617
rect 877 56493 917 56545
rect 969 56493 1041 56545
rect 1093 56493 1165 56545
rect 1217 56493 1289 56545
rect 1341 56493 1413 56545
rect 1465 56493 1537 56545
rect 1589 56493 1661 56545
rect 1713 56493 1785 56545
rect 1837 56493 1877 56545
rect 877 56421 1877 56493
rect 877 56369 917 56421
rect 969 56369 1041 56421
rect 1093 56369 1165 56421
rect 1217 56369 1289 56421
rect 1341 56369 1413 56421
rect 1465 56369 1537 56421
rect 1589 56369 1661 56421
rect 1713 56369 1785 56421
rect 1837 56369 1877 56421
rect 877 56297 1877 56369
rect 877 56245 917 56297
rect 969 56245 1041 56297
rect 1093 56245 1165 56297
rect 1217 56245 1289 56297
rect 1341 56245 1413 56297
rect 1465 56245 1537 56297
rect 1589 56245 1661 56297
rect 1713 56245 1785 56297
rect 1837 56245 1877 56297
rect 877 56173 1877 56245
rect 877 56121 917 56173
rect 969 56121 1041 56173
rect 1093 56121 1165 56173
rect 1217 56121 1289 56173
rect 1341 56121 1413 56173
rect 1465 56121 1537 56173
rect 1589 56121 1661 56173
rect 1713 56121 1785 56173
rect 1837 56121 1877 56173
rect 877 56049 1877 56121
rect 877 55997 917 56049
rect 969 55997 1041 56049
rect 1093 55997 1165 56049
rect 1217 55997 1289 56049
rect 1341 55997 1413 56049
rect 1465 55997 1537 56049
rect 1589 55997 1661 56049
rect 1713 55997 1785 56049
rect 1837 55997 1877 56049
rect 877 55925 1877 55997
rect 877 55873 917 55925
rect 969 55873 1041 55925
rect 1093 55873 1165 55925
rect 1217 55873 1289 55925
rect 1341 55873 1413 55925
rect 1465 55873 1537 55925
rect 1589 55873 1661 55925
rect 1713 55873 1785 55925
rect 1837 55873 1877 55925
rect 877 55801 1877 55873
rect 877 55749 917 55801
rect 969 55749 1041 55801
rect 1093 55749 1165 55801
rect 1217 55749 1289 55801
rect 1341 55749 1413 55801
rect 1465 55749 1537 55801
rect 1589 55749 1661 55801
rect 1713 55749 1785 55801
rect 1837 55749 1877 55801
rect 877 55677 1877 55749
rect 877 55625 917 55677
rect 969 55625 1041 55677
rect 1093 55625 1165 55677
rect 1217 55625 1289 55677
rect 1341 55625 1413 55677
rect 1465 55625 1537 55677
rect 1589 55625 1661 55677
rect 1713 55625 1785 55677
rect 1837 55625 1877 55677
rect 877 55553 1877 55625
rect 877 55501 917 55553
rect 969 55501 1041 55553
rect 1093 55501 1165 55553
rect 1217 55501 1289 55553
rect 1341 55501 1413 55553
rect 1465 55501 1537 55553
rect 1589 55501 1661 55553
rect 1713 55501 1785 55553
rect 1837 55501 1877 55553
rect 877 55429 1877 55501
rect 877 55377 917 55429
rect 969 55377 1041 55429
rect 1093 55377 1165 55429
rect 1217 55377 1289 55429
rect 1341 55377 1413 55429
rect 1465 55377 1537 55429
rect 1589 55377 1661 55429
rect 1713 55377 1785 55429
rect 1837 55377 1877 55429
rect 877 55305 1877 55377
rect 877 55253 917 55305
rect 969 55253 1041 55305
rect 1093 55253 1165 55305
rect 1217 55253 1289 55305
rect 1341 55253 1413 55305
rect 1465 55253 1537 55305
rect 1589 55253 1661 55305
rect 1713 55253 1785 55305
rect 1837 55253 1877 55305
rect 877 55181 1877 55253
rect 877 55129 917 55181
rect 969 55129 1041 55181
rect 1093 55129 1165 55181
rect 1217 55129 1289 55181
rect 1341 55129 1413 55181
rect 1465 55129 1537 55181
rect 1589 55129 1661 55181
rect 1713 55129 1785 55181
rect 1837 55129 1877 55181
rect 877 55057 1877 55129
rect 877 55005 917 55057
rect 969 55005 1041 55057
rect 1093 55005 1165 55057
rect 1217 55005 1289 55057
rect 1341 55005 1413 55057
rect 1465 55005 1537 55057
rect 1589 55005 1661 55057
rect 1713 55005 1785 55057
rect 1837 55005 1877 55057
rect 877 54933 1877 55005
rect 877 54881 917 54933
rect 969 54881 1041 54933
rect 1093 54881 1165 54933
rect 1217 54881 1289 54933
rect 1341 54881 1413 54933
rect 1465 54881 1537 54933
rect 1589 54881 1661 54933
rect 1713 54881 1785 54933
rect 1837 54881 1877 54933
rect 877 54809 1877 54881
rect 877 54757 917 54809
rect 969 54757 1041 54809
rect 1093 54757 1165 54809
rect 1217 54757 1289 54809
rect 1341 54757 1413 54809
rect 1465 54757 1537 54809
rect 1589 54757 1661 54809
rect 1713 54757 1785 54809
rect 1837 54757 1877 54809
rect 877 54685 1877 54757
rect 877 54633 917 54685
rect 969 54633 1041 54685
rect 1093 54633 1165 54685
rect 1217 54633 1289 54685
rect 1341 54633 1413 54685
rect 1465 54633 1537 54685
rect 1589 54633 1661 54685
rect 1713 54633 1785 54685
rect 1837 54633 1877 54685
rect 877 54561 1877 54633
rect 877 54509 917 54561
rect 969 54509 1041 54561
rect 1093 54509 1165 54561
rect 1217 54509 1289 54561
rect 1341 54509 1413 54561
rect 1465 54509 1537 54561
rect 1589 54509 1661 54561
rect 1713 54509 1785 54561
rect 1837 54509 1877 54561
rect 877 54437 1877 54509
rect 877 54385 917 54437
rect 969 54385 1041 54437
rect 1093 54385 1165 54437
rect 1217 54385 1289 54437
rect 1341 54385 1413 54437
rect 1465 54385 1537 54437
rect 1589 54385 1661 54437
rect 1713 54385 1785 54437
rect 1837 54385 1877 54437
rect 877 54313 1877 54385
rect 877 54261 917 54313
rect 969 54261 1041 54313
rect 1093 54261 1165 54313
rect 1217 54261 1289 54313
rect 1341 54261 1413 54313
rect 1465 54261 1537 54313
rect 1589 54261 1661 54313
rect 1713 54261 1785 54313
rect 1837 54261 1877 54313
rect 877 54189 1877 54261
rect 877 54137 917 54189
rect 969 54137 1041 54189
rect 1093 54137 1165 54189
rect 1217 54137 1289 54189
rect 1341 54137 1413 54189
rect 1465 54137 1537 54189
rect 1589 54137 1661 54189
rect 1713 54137 1785 54189
rect 1837 54137 1877 54189
rect 877 54065 1877 54137
rect 877 54013 917 54065
rect 969 54013 1041 54065
rect 1093 54013 1165 54065
rect 1217 54013 1289 54065
rect 1341 54013 1413 54065
rect 1465 54013 1537 54065
rect 1589 54013 1661 54065
rect 1713 54013 1785 54065
rect 1837 54013 1877 54065
rect 877 53941 1877 54013
rect 877 53889 917 53941
rect 969 53889 1041 53941
rect 1093 53889 1165 53941
rect 1217 53889 1289 53941
rect 1341 53889 1413 53941
rect 1465 53889 1537 53941
rect 1589 53889 1661 53941
rect 1713 53889 1785 53941
rect 1837 53889 1877 53941
rect 877 53817 1877 53889
rect 877 53765 917 53817
rect 969 53765 1041 53817
rect 1093 53765 1165 53817
rect 1217 53765 1289 53817
rect 1341 53765 1413 53817
rect 1465 53765 1537 53817
rect 1589 53765 1661 53817
rect 1713 53765 1785 53817
rect 1837 53765 1877 53817
rect 877 53693 1877 53765
rect 877 53641 917 53693
rect 969 53641 1041 53693
rect 1093 53641 1165 53693
rect 1217 53641 1289 53693
rect 1341 53641 1413 53693
rect 1465 53641 1537 53693
rect 1589 53641 1661 53693
rect 1713 53641 1785 53693
rect 1837 53641 1877 53693
rect 877 53633 1877 53641
rect 2793 56669 3793 56677
rect 2793 56617 2833 56669
rect 2885 56617 2957 56669
rect 3009 56617 3081 56669
rect 3133 56617 3205 56669
rect 3257 56617 3329 56669
rect 3381 56617 3453 56669
rect 3505 56617 3577 56669
rect 3629 56617 3701 56669
rect 3753 56617 3793 56669
rect 4313 56734 7229 56745
rect 4313 56688 4324 56734
rect 7218 56688 7229 56734
rect 4313 56677 7229 56688
rect 4313 56669 5313 56677
rect 2793 56545 3793 56617
rect 2793 56493 2833 56545
rect 2885 56493 2957 56545
rect 3009 56493 3081 56545
rect 3133 56493 3205 56545
rect 3257 56493 3329 56545
rect 3381 56493 3453 56545
rect 3505 56493 3577 56545
rect 3629 56493 3701 56545
rect 3753 56493 3793 56545
rect 2793 56421 3793 56493
rect 2793 56369 2833 56421
rect 2885 56369 2957 56421
rect 3009 56369 3081 56421
rect 3133 56369 3205 56421
rect 3257 56369 3329 56421
rect 3381 56369 3453 56421
rect 3505 56369 3577 56421
rect 3629 56369 3701 56421
rect 3753 56369 3793 56421
rect 2793 56297 3793 56369
rect 2793 56245 2833 56297
rect 2885 56245 2957 56297
rect 3009 56245 3081 56297
rect 3133 56245 3205 56297
rect 3257 56245 3329 56297
rect 3381 56245 3453 56297
rect 3505 56245 3577 56297
rect 3629 56245 3701 56297
rect 3753 56245 3793 56297
rect 2793 56173 3793 56245
rect 2793 56121 2833 56173
rect 2885 56121 2957 56173
rect 3009 56121 3081 56173
rect 3133 56121 3205 56173
rect 3257 56121 3329 56173
rect 3381 56121 3453 56173
rect 3505 56121 3577 56173
rect 3629 56121 3701 56173
rect 3753 56121 3793 56173
rect 2793 56049 3793 56121
rect 2793 55997 2833 56049
rect 2885 55997 2957 56049
rect 3009 55997 3081 56049
rect 3133 55997 3205 56049
rect 3257 55997 3329 56049
rect 3381 55997 3453 56049
rect 3505 55997 3577 56049
rect 3629 55997 3701 56049
rect 3753 55997 3793 56049
rect 2793 55925 3793 55997
rect 2793 55873 2833 55925
rect 2885 55873 2957 55925
rect 3009 55873 3081 55925
rect 3133 55873 3205 55925
rect 3257 55873 3329 55925
rect 3381 55873 3453 55925
rect 3505 55873 3577 55925
rect 3629 55873 3701 55925
rect 3753 55873 3793 55925
rect 2793 55801 3793 55873
rect 2793 55749 2833 55801
rect 2885 55749 2957 55801
rect 3009 55749 3081 55801
rect 3133 55749 3205 55801
rect 3257 55749 3329 55801
rect 3381 55749 3453 55801
rect 3505 55749 3577 55801
rect 3629 55749 3701 55801
rect 3753 55749 3793 55801
rect 2793 55677 3793 55749
rect 2793 55625 2833 55677
rect 2885 55625 2957 55677
rect 3009 55625 3081 55677
rect 3133 55625 3205 55677
rect 3257 55625 3329 55677
rect 3381 55625 3453 55677
rect 3505 55625 3577 55677
rect 3629 55625 3701 55677
rect 3753 55625 3793 55677
rect 2793 55553 3793 55625
rect 2793 55501 2833 55553
rect 2885 55501 2957 55553
rect 3009 55501 3081 55553
rect 3133 55501 3205 55553
rect 3257 55501 3329 55553
rect 3381 55501 3453 55553
rect 3505 55501 3577 55553
rect 3629 55501 3701 55553
rect 3753 55501 3793 55553
rect 2793 55429 3793 55501
rect 2793 55377 2833 55429
rect 2885 55377 2957 55429
rect 3009 55377 3081 55429
rect 3133 55377 3205 55429
rect 3257 55377 3329 55429
rect 3381 55377 3453 55429
rect 3505 55377 3577 55429
rect 3629 55377 3701 55429
rect 3753 55377 3793 55429
rect 2793 55305 3793 55377
rect 2793 55253 2833 55305
rect 2885 55253 2957 55305
rect 3009 55253 3081 55305
rect 3133 55253 3205 55305
rect 3257 55253 3329 55305
rect 3381 55253 3453 55305
rect 3505 55253 3577 55305
rect 3629 55253 3701 55305
rect 3753 55253 3793 55305
rect 2793 55181 3793 55253
rect 2793 55129 2833 55181
rect 2885 55129 2957 55181
rect 3009 55129 3081 55181
rect 3133 55129 3205 55181
rect 3257 55129 3329 55181
rect 3381 55129 3453 55181
rect 3505 55129 3577 55181
rect 3629 55129 3701 55181
rect 3753 55129 3793 55181
rect 2793 55057 3793 55129
rect 2793 55005 2833 55057
rect 2885 55005 2957 55057
rect 3009 55005 3081 55057
rect 3133 55005 3205 55057
rect 3257 55005 3329 55057
rect 3381 55005 3453 55057
rect 3505 55005 3577 55057
rect 3629 55005 3701 55057
rect 3753 55005 3793 55057
rect 2793 54933 3793 55005
rect 2793 54881 2833 54933
rect 2885 54881 2957 54933
rect 3009 54881 3081 54933
rect 3133 54881 3205 54933
rect 3257 54881 3329 54933
rect 3381 54881 3453 54933
rect 3505 54881 3577 54933
rect 3629 54881 3701 54933
rect 3753 54881 3793 54933
rect 2793 54809 3793 54881
rect 2793 54757 2833 54809
rect 2885 54757 2957 54809
rect 3009 54757 3081 54809
rect 3133 54757 3205 54809
rect 3257 54757 3329 54809
rect 3381 54757 3453 54809
rect 3505 54757 3577 54809
rect 3629 54757 3701 54809
rect 3753 54757 3793 54809
rect 2793 54685 3793 54757
rect 2793 54633 2833 54685
rect 2885 54633 2957 54685
rect 3009 54633 3081 54685
rect 3133 54633 3205 54685
rect 3257 54633 3329 54685
rect 3381 54633 3453 54685
rect 3505 54633 3577 54685
rect 3629 54633 3701 54685
rect 3753 54633 3793 54685
rect 2793 54561 3793 54633
rect 2793 54509 2833 54561
rect 2885 54509 2957 54561
rect 3009 54509 3081 54561
rect 3133 54509 3205 54561
rect 3257 54509 3329 54561
rect 3381 54509 3453 54561
rect 3505 54509 3577 54561
rect 3629 54509 3701 54561
rect 3753 54509 3793 54561
rect 2793 54437 3793 54509
rect 2793 54385 2833 54437
rect 2885 54385 2957 54437
rect 3009 54385 3081 54437
rect 3133 54385 3205 54437
rect 3257 54385 3329 54437
rect 3381 54385 3453 54437
rect 3505 54385 3577 54437
rect 3629 54385 3701 54437
rect 3753 54385 3793 54437
rect 2793 54313 3793 54385
rect 2793 54261 2833 54313
rect 2885 54261 2957 54313
rect 3009 54261 3081 54313
rect 3133 54261 3205 54313
rect 3257 54261 3329 54313
rect 3381 54261 3453 54313
rect 3505 54261 3577 54313
rect 3629 54261 3701 54313
rect 3753 54261 3793 54313
rect 2793 54189 3793 54261
rect 2793 54137 2833 54189
rect 2885 54137 2957 54189
rect 3009 54137 3081 54189
rect 3133 54137 3205 54189
rect 3257 54137 3329 54189
rect 3381 54137 3453 54189
rect 3505 54137 3577 54189
rect 3629 54137 3701 54189
rect 3753 54137 3793 54189
rect 2793 54065 3793 54137
rect 2793 54013 2833 54065
rect 2885 54013 2957 54065
rect 3009 54013 3081 54065
rect 3133 54013 3205 54065
rect 3257 54013 3329 54065
rect 3381 54013 3453 54065
rect 3505 54013 3577 54065
rect 3629 54013 3701 54065
rect 3753 54013 3793 54065
rect 2793 53941 3793 54013
rect 2793 53889 2833 53941
rect 2885 53889 2957 53941
rect 3009 53889 3081 53941
rect 3133 53889 3205 53941
rect 3257 53889 3329 53941
rect 3381 53889 3453 53941
rect 3505 53889 3577 53941
rect 3629 53889 3701 53941
rect 3753 53889 3793 53941
rect 2793 53817 3793 53889
rect 2793 53765 2833 53817
rect 2885 53765 2957 53817
rect 3009 53765 3081 53817
rect 3133 53765 3205 53817
rect 3257 53765 3329 53817
rect 3381 53765 3453 53817
rect 3505 53765 3577 53817
rect 3629 53765 3701 53817
rect 3753 53765 3793 53817
rect 2793 53693 3793 53765
rect 2793 53641 2833 53693
rect 2885 53641 2957 53693
rect 3009 53641 3081 53693
rect 3133 53641 3205 53693
rect 3257 53641 3329 53693
rect 3381 53641 3453 53693
rect 3505 53641 3577 53693
rect 3629 53641 3701 53693
rect 3753 53641 3793 53693
rect 2793 53633 3793 53641
rect 877 53622 3793 53633
rect 877 53576 888 53622
rect 3782 53576 3793 53622
rect 877 53565 3793 53576
rect 3853 56618 4253 56655
rect 3853 53692 3864 56618
rect 3910 53692 4196 56618
rect 4242 53692 4253 56618
rect 3853 53505 4253 53692
rect 4313 56617 4340 56669
rect 4392 56617 4464 56669
rect 4516 56617 4588 56669
rect 4640 56617 4712 56669
rect 4764 56617 5313 56669
rect 4313 56545 5313 56617
rect 4313 56493 4340 56545
rect 4392 56493 4464 56545
rect 4516 56493 4588 56545
rect 4640 56493 4712 56545
rect 4764 56493 5313 56545
rect 4313 56421 5313 56493
rect 4313 56369 4340 56421
rect 4392 56369 4464 56421
rect 4516 56369 4588 56421
rect 4640 56369 4712 56421
rect 4764 56369 5313 56421
rect 4313 56297 5313 56369
rect 4313 56245 4340 56297
rect 4392 56245 4464 56297
rect 4516 56245 4588 56297
rect 4640 56245 4712 56297
rect 4764 56245 5313 56297
rect 4313 56173 5313 56245
rect 4313 56121 4340 56173
rect 4392 56121 4464 56173
rect 4516 56121 4588 56173
rect 4640 56121 4712 56173
rect 4764 56121 5313 56173
rect 4313 56049 5313 56121
rect 4313 55997 4340 56049
rect 4392 55997 4464 56049
rect 4516 55997 4588 56049
rect 4640 55997 4712 56049
rect 4764 55997 5313 56049
rect 4313 55925 5313 55997
rect 4313 55873 4340 55925
rect 4392 55873 4464 55925
rect 4516 55873 4588 55925
rect 4640 55873 4712 55925
rect 4764 55873 5313 55925
rect 4313 55801 5313 55873
rect 4313 55749 4340 55801
rect 4392 55749 4464 55801
rect 4516 55749 4588 55801
rect 4640 55749 4712 55801
rect 4764 55749 5313 55801
rect 4313 55677 5313 55749
rect 4313 55625 4340 55677
rect 4392 55625 4464 55677
rect 4516 55625 4588 55677
rect 4640 55625 4712 55677
rect 4764 55625 5313 55677
rect 4313 55553 5313 55625
rect 4313 55501 4340 55553
rect 4392 55501 4464 55553
rect 4516 55501 4588 55553
rect 4640 55501 4712 55553
rect 4764 55501 5313 55553
rect 4313 55429 5313 55501
rect 4313 55377 4340 55429
rect 4392 55377 4464 55429
rect 4516 55377 4588 55429
rect 4640 55377 4712 55429
rect 4764 55377 5313 55429
rect 4313 55305 5313 55377
rect 4313 55253 4340 55305
rect 4392 55253 4464 55305
rect 4516 55253 4588 55305
rect 4640 55253 4712 55305
rect 4764 55253 5313 55305
rect 4313 55181 5313 55253
rect 4313 55129 4340 55181
rect 4392 55129 4464 55181
rect 4516 55129 4588 55181
rect 4640 55129 4712 55181
rect 4764 55129 5313 55181
rect 4313 55057 5313 55129
rect 4313 55005 4340 55057
rect 4392 55005 4464 55057
rect 4516 55005 4588 55057
rect 4640 55005 4712 55057
rect 4764 55005 5313 55057
rect 4313 54933 5313 55005
rect 4313 54881 4340 54933
rect 4392 54881 4464 54933
rect 4516 54881 4588 54933
rect 4640 54881 4712 54933
rect 4764 54881 5313 54933
rect 4313 54809 5313 54881
rect 4313 54757 4340 54809
rect 4392 54757 4464 54809
rect 4516 54757 4588 54809
rect 4640 54757 4712 54809
rect 4764 54757 5313 54809
rect 4313 54685 5313 54757
rect 4313 54633 4340 54685
rect 4392 54633 4464 54685
rect 4516 54633 4588 54685
rect 4640 54633 4712 54685
rect 4764 54633 5313 54685
rect 4313 54561 5313 54633
rect 4313 54509 4340 54561
rect 4392 54509 4464 54561
rect 4516 54509 4588 54561
rect 4640 54509 4712 54561
rect 4764 54509 5313 54561
rect 4313 54437 5313 54509
rect 4313 54385 4340 54437
rect 4392 54385 4464 54437
rect 4516 54385 4588 54437
rect 4640 54385 4712 54437
rect 4764 54385 5313 54437
rect 4313 54313 5313 54385
rect 4313 54261 4340 54313
rect 4392 54261 4464 54313
rect 4516 54261 4588 54313
rect 4640 54261 4712 54313
rect 4764 54261 5313 54313
rect 4313 54189 5313 54261
rect 4313 54137 4340 54189
rect 4392 54137 4464 54189
rect 4516 54137 4588 54189
rect 4640 54137 4712 54189
rect 4764 54137 5313 54189
rect 4313 54065 5313 54137
rect 4313 54013 4340 54065
rect 4392 54013 4464 54065
rect 4516 54013 4588 54065
rect 4640 54013 4712 54065
rect 4764 54013 5313 54065
rect 4313 53941 5313 54013
rect 4313 53889 4340 53941
rect 4392 53889 4464 53941
rect 4516 53889 4588 53941
rect 4640 53889 4712 53941
rect 4764 53889 5313 53941
rect 4313 53817 5313 53889
rect 4313 53765 4340 53817
rect 4392 53765 4464 53817
rect 4516 53765 4588 53817
rect 4640 53765 4712 53817
rect 4764 53765 5313 53817
rect 4313 53693 5313 53765
rect 4313 53641 4340 53693
rect 4392 53641 4464 53693
rect 4516 53641 4588 53693
rect 4640 53641 4712 53693
rect 4764 53641 5313 53693
rect 4313 53633 5313 53641
rect 6229 56669 7229 56677
rect 6229 56617 6297 56669
rect 6349 56617 6421 56669
rect 6473 56617 6545 56669
rect 6597 56617 6669 56669
rect 6721 56617 6793 56669
rect 6845 56617 6917 56669
rect 6969 56617 7041 56669
rect 7093 56617 7229 56669
rect 7749 56734 10665 56745
rect 7749 56688 7760 56734
rect 10654 56688 10665 56734
rect 7749 56677 10665 56688
rect 7749 56669 8749 56677
rect 6229 56545 7229 56617
rect 6229 56493 6297 56545
rect 6349 56493 6421 56545
rect 6473 56493 6545 56545
rect 6597 56493 6669 56545
rect 6721 56493 6793 56545
rect 6845 56493 6917 56545
rect 6969 56493 7041 56545
rect 7093 56493 7229 56545
rect 6229 56421 7229 56493
rect 6229 56369 6297 56421
rect 6349 56369 6421 56421
rect 6473 56369 6545 56421
rect 6597 56369 6669 56421
rect 6721 56369 6793 56421
rect 6845 56369 6917 56421
rect 6969 56369 7041 56421
rect 7093 56369 7229 56421
rect 6229 56297 7229 56369
rect 6229 56245 6297 56297
rect 6349 56245 6421 56297
rect 6473 56245 6545 56297
rect 6597 56245 6669 56297
rect 6721 56245 6793 56297
rect 6845 56245 6917 56297
rect 6969 56245 7041 56297
rect 7093 56245 7229 56297
rect 6229 56173 7229 56245
rect 6229 56121 6297 56173
rect 6349 56121 6421 56173
rect 6473 56121 6545 56173
rect 6597 56121 6669 56173
rect 6721 56121 6793 56173
rect 6845 56121 6917 56173
rect 6969 56121 7041 56173
rect 7093 56121 7229 56173
rect 6229 56049 7229 56121
rect 6229 55997 6297 56049
rect 6349 55997 6421 56049
rect 6473 55997 6545 56049
rect 6597 55997 6669 56049
rect 6721 55997 6793 56049
rect 6845 55997 6917 56049
rect 6969 55997 7041 56049
rect 7093 55997 7229 56049
rect 6229 55925 7229 55997
rect 6229 55873 6297 55925
rect 6349 55873 6421 55925
rect 6473 55873 6545 55925
rect 6597 55873 6669 55925
rect 6721 55873 6793 55925
rect 6845 55873 6917 55925
rect 6969 55873 7041 55925
rect 7093 55873 7229 55925
rect 6229 55801 7229 55873
rect 6229 55749 6297 55801
rect 6349 55749 6421 55801
rect 6473 55749 6545 55801
rect 6597 55749 6669 55801
rect 6721 55749 6793 55801
rect 6845 55749 6917 55801
rect 6969 55749 7041 55801
rect 7093 55749 7229 55801
rect 6229 55677 7229 55749
rect 6229 55625 6297 55677
rect 6349 55625 6421 55677
rect 6473 55625 6545 55677
rect 6597 55625 6669 55677
rect 6721 55625 6793 55677
rect 6845 55625 6917 55677
rect 6969 55625 7041 55677
rect 7093 55625 7229 55677
rect 6229 55553 7229 55625
rect 6229 55501 6297 55553
rect 6349 55501 6421 55553
rect 6473 55501 6545 55553
rect 6597 55501 6669 55553
rect 6721 55501 6793 55553
rect 6845 55501 6917 55553
rect 6969 55501 7041 55553
rect 7093 55501 7229 55553
rect 6229 55429 7229 55501
rect 6229 55377 6297 55429
rect 6349 55377 6421 55429
rect 6473 55377 6545 55429
rect 6597 55377 6669 55429
rect 6721 55377 6793 55429
rect 6845 55377 6917 55429
rect 6969 55377 7041 55429
rect 7093 55377 7229 55429
rect 6229 55305 7229 55377
rect 6229 55253 6297 55305
rect 6349 55253 6421 55305
rect 6473 55253 6545 55305
rect 6597 55253 6669 55305
rect 6721 55253 6793 55305
rect 6845 55253 6917 55305
rect 6969 55253 7041 55305
rect 7093 55253 7229 55305
rect 6229 55181 7229 55253
rect 6229 55129 6297 55181
rect 6349 55129 6421 55181
rect 6473 55129 6545 55181
rect 6597 55129 6669 55181
rect 6721 55129 6793 55181
rect 6845 55129 6917 55181
rect 6969 55129 7041 55181
rect 7093 55129 7229 55181
rect 6229 55057 7229 55129
rect 6229 55005 6297 55057
rect 6349 55005 6421 55057
rect 6473 55005 6545 55057
rect 6597 55005 6669 55057
rect 6721 55005 6793 55057
rect 6845 55005 6917 55057
rect 6969 55005 7041 55057
rect 7093 55005 7229 55057
rect 6229 54933 7229 55005
rect 6229 54881 6297 54933
rect 6349 54881 6421 54933
rect 6473 54881 6545 54933
rect 6597 54881 6669 54933
rect 6721 54881 6793 54933
rect 6845 54881 6917 54933
rect 6969 54881 7041 54933
rect 7093 54881 7229 54933
rect 6229 54809 7229 54881
rect 6229 54757 6297 54809
rect 6349 54757 6421 54809
rect 6473 54757 6545 54809
rect 6597 54757 6669 54809
rect 6721 54757 6793 54809
rect 6845 54757 6917 54809
rect 6969 54757 7041 54809
rect 7093 54757 7229 54809
rect 6229 54685 7229 54757
rect 6229 54633 6297 54685
rect 6349 54633 6421 54685
rect 6473 54633 6545 54685
rect 6597 54633 6669 54685
rect 6721 54633 6793 54685
rect 6845 54633 6917 54685
rect 6969 54633 7041 54685
rect 7093 54633 7229 54685
rect 6229 54561 7229 54633
rect 6229 54509 6297 54561
rect 6349 54509 6421 54561
rect 6473 54509 6545 54561
rect 6597 54509 6669 54561
rect 6721 54509 6793 54561
rect 6845 54509 6917 54561
rect 6969 54509 7041 54561
rect 7093 54509 7229 54561
rect 6229 54437 7229 54509
rect 6229 54385 6297 54437
rect 6349 54385 6421 54437
rect 6473 54385 6545 54437
rect 6597 54385 6669 54437
rect 6721 54385 6793 54437
rect 6845 54385 6917 54437
rect 6969 54385 7041 54437
rect 7093 54385 7229 54437
rect 6229 54313 7229 54385
rect 6229 54261 6297 54313
rect 6349 54261 6421 54313
rect 6473 54261 6545 54313
rect 6597 54261 6669 54313
rect 6721 54261 6793 54313
rect 6845 54261 6917 54313
rect 6969 54261 7041 54313
rect 7093 54261 7229 54313
rect 6229 54189 7229 54261
rect 6229 54137 6297 54189
rect 6349 54137 6421 54189
rect 6473 54137 6545 54189
rect 6597 54137 6669 54189
rect 6721 54137 6793 54189
rect 6845 54137 6917 54189
rect 6969 54137 7041 54189
rect 7093 54137 7229 54189
rect 6229 54065 7229 54137
rect 6229 54013 6297 54065
rect 6349 54013 6421 54065
rect 6473 54013 6545 54065
rect 6597 54013 6669 54065
rect 6721 54013 6793 54065
rect 6845 54013 6917 54065
rect 6969 54013 7041 54065
rect 7093 54013 7229 54065
rect 6229 53941 7229 54013
rect 6229 53889 6297 53941
rect 6349 53889 6421 53941
rect 6473 53889 6545 53941
rect 6597 53889 6669 53941
rect 6721 53889 6793 53941
rect 6845 53889 6917 53941
rect 6969 53889 7041 53941
rect 7093 53889 7229 53941
rect 6229 53817 7229 53889
rect 6229 53765 6297 53817
rect 6349 53765 6421 53817
rect 6473 53765 6545 53817
rect 6597 53765 6669 53817
rect 6721 53765 6793 53817
rect 6845 53765 6917 53817
rect 6969 53765 7041 53817
rect 7093 53765 7229 53817
rect 6229 53693 7229 53765
rect 6229 53641 6297 53693
rect 6349 53641 6421 53693
rect 6473 53641 6545 53693
rect 6597 53641 6669 53693
rect 6721 53641 6793 53693
rect 6845 53641 6917 53693
rect 6969 53641 7041 53693
rect 7093 53641 7229 53693
rect 6229 53633 7229 53641
rect 4313 53622 7229 53633
rect 4313 53576 4324 53622
rect 7218 53576 7229 53622
rect 4313 53565 7229 53576
rect 7289 56618 7689 56655
rect 7289 53692 7300 56618
rect 7346 53692 7632 56618
rect 7678 53692 7689 56618
rect 7289 53505 7689 53692
rect 7749 56617 7885 56669
rect 7937 56617 8009 56669
rect 8061 56617 8133 56669
rect 8185 56617 8257 56669
rect 8309 56617 8381 56669
rect 8433 56617 8505 56669
rect 8557 56617 8629 56669
rect 8681 56617 8749 56669
rect 7749 56545 8749 56617
rect 7749 56493 7885 56545
rect 7937 56493 8009 56545
rect 8061 56493 8133 56545
rect 8185 56493 8257 56545
rect 8309 56493 8381 56545
rect 8433 56493 8505 56545
rect 8557 56493 8629 56545
rect 8681 56493 8749 56545
rect 7749 56421 8749 56493
rect 7749 56369 7885 56421
rect 7937 56369 8009 56421
rect 8061 56369 8133 56421
rect 8185 56369 8257 56421
rect 8309 56369 8381 56421
rect 8433 56369 8505 56421
rect 8557 56369 8629 56421
rect 8681 56369 8749 56421
rect 7749 56297 8749 56369
rect 7749 56245 7885 56297
rect 7937 56245 8009 56297
rect 8061 56245 8133 56297
rect 8185 56245 8257 56297
rect 8309 56245 8381 56297
rect 8433 56245 8505 56297
rect 8557 56245 8629 56297
rect 8681 56245 8749 56297
rect 7749 56173 8749 56245
rect 7749 56121 7885 56173
rect 7937 56121 8009 56173
rect 8061 56121 8133 56173
rect 8185 56121 8257 56173
rect 8309 56121 8381 56173
rect 8433 56121 8505 56173
rect 8557 56121 8629 56173
rect 8681 56121 8749 56173
rect 7749 56049 8749 56121
rect 7749 55997 7885 56049
rect 7937 55997 8009 56049
rect 8061 55997 8133 56049
rect 8185 55997 8257 56049
rect 8309 55997 8381 56049
rect 8433 55997 8505 56049
rect 8557 55997 8629 56049
rect 8681 55997 8749 56049
rect 7749 55925 8749 55997
rect 7749 55873 7885 55925
rect 7937 55873 8009 55925
rect 8061 55873 8133 55925
rect 8185 55873 8257 55925
rect 8309 55873 8381 55925
rect 8433 55873 8505 55925
rect 8557 55873 8629 55925
rect 8681 55873 8749 55925
rect 7749 55801 8749 55873
rect 7749 55749 7885 55801
rect 7937 55749 8009 55801
rect 8061 55749 8133 55801
rect 8185 55749 8257 55801
rect 8309 55749 8381 55801
rect 8433 55749 8505 55801
rect 8557 55749 8629 55801
rect 8681 55749 8749 55801
rect 7749 55677 8749 55749
rect 7749 55625 7885 55677
rect 7937 55625 8009 55677
rect 8061 55625 8133 55677
rect 8185 55625 8257 55677
rect 8309 55625 8381 55677
rect 8433 55625 8505 55677
rect 8557 55625 8629 55677
rect 8681 55625 8749 55677
rect 7749 55553 8749 55625
rect 7749 55501 7885 55553
rect 7937 55501 8009 55553
rect 8061 55501 8133 55553
rect 8185 55501 8257 55553
rect 8309 55501 8381 55553
rect 8433 55501 8505 55553
rect 8557 55501 8629 55553
rect 8681 55501 8749 55553
rect 7749 55429 8749 55501
rect 7749 55377 7885 55429
rect 7937 55377 8009 55429
rect 8061 55377 8133 55429
rect 8185 55377 8257 55429
rect 8309 55377 8381 55429
rect 8433 55377 8505 55429
rect 8557 55377 8629 55429
rect 8681 55377 8749 55429
rect 7749 55305 8749 55377
rect 7749 55253 7885 55305
rect 7937 55253 8009 55305
rect 8061 55253 8133 55305
rect 8185 55253 8257 55305
rect 8309 55253 8381 55305
rect 8433 55253 8505 55305
rect 8557 55253 8629 55305
rect 8681 55253 8749 55305
rect 7749 55181 8749 55253
rect 7749 55129 7885 55181
rect 7937 55129 8009 55181
rect 8061 55129 8133 55181
rect 8185 55129 8257 55181
rect 8309 55129 8381 55181
rect 8433 55129 8505 55181
rect 8557 55129 8629 55181
rect 8681 55129 8749 55181
rect 7749 55057 8749 55129
rect 7749 55005 7885 55057
rect 7937 55005 8009 55057
rect 8061 55005 8133 55057
rect 8185 55005 8257 55057
rect 8309 55005 8381 55057
rect 8433 55005 8505 55057
rect 8557 55005 8629 55057
rect 8681 55005 8749 55057
rect 7749 54933 8749 55005
rect 7749 54881 7885 54933
rect 7937 54881 8009 54933
rect 8061 54881 8133 54933
rect 8185 54881 8257 54933
rect 8309 54881 8381 54933
rect 8433 54881 8505 54933
rect 8557 54881 8629 54933
rect 8681 54881 8749 54933
rect 7749 54809 8749 54881
rect 7749 54757 7885 54809
rect 7937 54757 8009 54809
rect 8061 54757 8133 54809
rect 8185 54757 8257 54809
rect 8309 54757 8381 54809
rect 8433 54757 8505 54809
rect 8557 54757 8629 54809
rect 8681 54757 8749 54809
rect 7749 54685 8749 54757
rect 7749 54633 7885 54685
rect 7937 54633 8009 54685
rect 8061 54633 8133 54685
rect 8185 54633 8257 54685
rect 8309 54633 8381 54685
rect 8433 54633 8505 54685
rect 8557 54633 8629 54685
rect 8681 54633 8749 54685
rect 7749 54561 8749 54633
rect 7749 54509 7885 54561
rect 7937 54509 8009 54561
rect 8061 54509 8133 54561
rect 8185 54509 8257 54561
rect 8309 54509 8381 54561
rect 8433 54509 8505 54561
rect 8557 54509 8629 54561
rect 8681 54509 8749 54561
rect 7749 54437 8749 54509
rect 7749 54385 7885 54437
rect 7937 54385 8009 54437
rect 8061 54385 8133 54437
rect 8185 54385 8257 54437
rect 8309 54385 8381 54437
rect 8433 54385 8505 54437
rect 8557 54385 8629 54437
rect 8681 54385 8749 54437
rect 7749 54313 8749 54385
rect 7749 54261 7885 54313
rect 7937 54261 8009 54313
rect 8061 54261 8133 54313
rect 8185 54261 8257 54313
rect 8309 54261 8381 54313
rect 8433 54261 8505 54313
rect 8557 54261 8629 54313
rect 8681 54261 8749 54313
rect 7749 54189 8749 54261
rect 7749 54137 7885 54189
rect 7937 54137 8009 54189
rect 8061 54137 8133 54189
rect 8185 54137 8257 54189
rect 8309 54137 8381 54189
rect 8433 54137 8505 54189
rect 8557 54137 8629 54189
rect 8681 54137 8749 54189
rect 7749 54065 8749 54137
rect 7749 54013 7885 54065
rect 7937 54013 8009 54065
rect 8061 54013 8133 54065
rect 8185 54013 8257 54065
rect 8309 54013 8381 54065
rect 8433 54013 8505 54065
rect 8557 54013 8629 54065
rect 8681 54013 8749 54065
rect 7749 53941 8749 54013
rect 7749 53889 7885 53941
rect 7937 53889 8009 53941
rect 8061 53889 8133 53941
rect 8185 53889 8257 53941
rect 8309 53889 8381 53941
rect 8433 53889 8505 53941
rect 8557 53889 8629 53941
rect 8681 53889 8749 53941
rect 7749 53817 8749 53889
rect 7749 53765 7885 53817
rect 7937 53765 8009 53817
rect 8061 53765 8133 53817
rect 8185 53765 8257 53817
rect 8309 53765 8381 53817
rect 8433 53765 8505 53817
rect 8557 53765 8629 53817
rect 8681 53765 8749 53817
rect 7749 53693 8749 53765
rect 7749 53641 7885 53693
rect 7937 53641 8009 53693
rect 8061 53641 8133 53693
rect 8185 53641 8257 53693
rect 8309 53641 8381 53693
rect 8433 53641 8505 53693
rect 8557 53641 8629 53693
rect 8681 53641 8749 53693
rect 7749 53633 8749 53641
rect 9665 56669 10665 56677
rect 9665 56617 10214 56669
rect 10266 56617 10338 56669
rect 10390 56617 10462 56669
rect 10514 56617 10586 56669
rect 10638 56617 10665 56669
rect 11185 56734 14101 56745
rect 11185 56688 11196 56734
rect 14090 56688 14101 56734
rect 11185 56677 14101 56688
rect 11185 56669 12185 56677
rect 9665 56545 10665 56617
rect 9665 56493 10214 56545
rect 10266 56493 10338 56545
rect 10390 56493 10462 56545
rect 10514 56493 10586 56545
rect 10638 56493 10665 56545
rect 9665 56421 10665 56493
rect 9665 56369 10214 56421
rect 10266 56369 10338 56421
rect 10390 56369 10462 56421
rect 10514 56369 10586 56421
rect 10638 56369 10665 56421
rect 9665 56297 10665 56369
rect 9665 56245 10214 56297
rect 10266 56245 10338 56297
rect 10390 56245 10462 56297
rect 10514 56245 10586 56297
rect 10638 56245 10665 56297
rect 9665 56173 10665 56245
rect 9665 56121 10214 56173
rect 10266 56121 10338 56173
rect 10390 56121 10462 56173
rect 10514 56121 10586 56173
rect 10638 56121 10665 56173
rect 9665 56049 10665 56121
rect 9665 55997 10214 56049
rect 10266 55997 10338 56049
rect 10390 55997 10462 56049
rect 10514 55997 10586 56049
rect 10638 55997 10665 56049
rect 9665 55925 10665 55997
rect 9665 55873 10214 55925
rect 10266 55873 10338 55925
rect 10390 55873 10462 55925
rect 10514 55873 10586 55925
rect 10638 55873 10665 55925
rect 9665 55801 10665 55873
rect 9665 55749 10214 55801
rect 10266 55749 10338 55801
rect 10390 55749 10462 55801
rect 10514 55749 10586 55801
rect 10638 55749 10665 55801
rect 9665 55677 10665 55749
rect 9665 55625 10214 55677
rect 10266 55625 10338 55677
rect 10390 55625 10462 55677
rect 10514 55625 10586 55677
rect 10638 55625 10665 55677
rect 9665 55553 10665 55625
rect 9665 55501 10214 55553
rect 10266 55501 10338 55553
rect 10390 55501 10462 55553
rect 10514 55501 10586 55553
rect 10638 55501 10665 55553
rect 9665 55429 10665 55501
rect 9665 55377 10214 55429
rect 10266 55377 10338 55429
rect 10390 55377 10462 55429
rect 10514 55377 10586 55429
rect 10638 55377 10665 55429
rect 9665 55305 10665 55377
rect 9665 55253 10214 55305
rect 10266 55253 10338 55305
rect 10390 55253 10462 55305
rect 10514 55253 10586 55305
rect 10638 55253 10665 55305
rect 9665 55181 10665 55253
rect 9665 55129 10214 55181
rect 10266 55129 10338 55181
rect 10390 55129 10462 55181
rect 10514 55129 10586 55181
rect 10638 55129 10665 55181
rect 9665 55057 10665 55129
rect 9665 55005 10214 55057
rect 10266 55005 10338 55057
rect 10390 55005 10462 55057
rect 10514 55005 10586 55057
rect 10638 55005 10665 55057
rect 9665 54933 10665 55005
rect 9665 54881 10214 54933
rect 10266 54881 10338 54933
rect 10390 54881 10462 54933
rect 10514 54881 10586 54933
rect 10638 54881 10665 54933
rect 9665 54809 10665 54881
rect 9665 54757 10214 54809
rect 10266 54757 10338 54809
rect 10390 54757 10462 54809
rect 10514 54757 10586 54809
rect 10638 54757 10665 54809
rect 9665 54685 10665 54757
rect 9665 54633 10214 54685
rect 10266 54633 10338 54685
rect 10390 54633 10462 54685
rect 10514 54633 10586 54685
rect 10638 54633 10665 54685
rect 9665 54561 10665 54633
rect 9665 54509 10214 54561
rect 10266 54509 10338 54561
rect 10390 54509 10462 54561
rect 10514 54509 10586 54561
rect 10638 54509 10665 54561
rect 9665 54437 10665 54509
rect 9665 54385 10214 54437
rect 10266 54385 10338 54437
rect 10390 54385 10462 54437
rect 10514 54385 10586 54437
rect 10638 54385 10665 54437
rect 9665 54313 10665 54385
rect 9665 54261 10214 54313
rect 10266 54261 10338 54313
rect 10390 54261 10462 54313
rect 10514 54261 10586 54313
rect 10638 54261 10665 54313
rect 9665 54189 10665 54261
rect 9665 54137 10214 54189
rect 10266 54137 10338 54189
rect 10390 54137 10462 54189
rect 10514 54137 10586 54189
rect 10638 54137 10665 54189
rect 9665 54065 10665 54137
rect 9665 54013 10214 54065
rect 10266 54013 10338 54065
rect 10390 54013 10462 54065
rect 10514 54013 10586 54065
rect 10638 54013 10665 54065
rect 9665 53941 10665 54013
rect 9665 53889 10214 53941
rect 10266 53889 10338 53941
rect 10390 53889 10462 53941
rect 10514 53889 10586 53941
rect 10638 53889 10665 53941
rect 9665 53817 10665 53889
rect 9665 53765 10214 53817
rect 10266 53765 10338 53817
rect 10390 53765 10462 53817
rect 10514 53765 10586 53817
rect 10638 53765 10665 53817
rect 9665 53693 10665 53765
rect 9665 53641 10214 53693
rect 10266 53641 10338 53693
rect 10390 53641 10462 53693
rect 10514 53641 10586 53693
rect 10638 53641 10665 53693
rect 9665 53633 10665 53641
rect 7749 53622 10665 53633
rect 7749 53576 7760 53622
rect 10654 53576 10665 53622
rect 7749 53565 10665 53576
rect 10725 56618 11125 56655
rect 10725 53692 10736 56618
rect 10782 53692 11068 56618
rect 11114 53692 11125 56618
rect 10725 53505 11125 53692
rect 11185 56617 11225 56669
rect 11277 56617 11349 56669
rect 11401 56617 11473 56669
rect 11525 56617 11597 56669
rect 11649 56617 11721 56669
rect 11773 56617 11845 56669
rect 11897 56617 11969 56669
rect 12021 56617 12093 56669
rect 12145 56617 12185 56669
rect 11185 56545 12185 56617
rect 11185 56493 11225 56545
rect 11277 56493 11349 56545
rect 11401 56493 11473 56545
rect 11525 56493 11597 56545
rect 11649 56493 11721 56545
rect 11773 56493 11845 56545
rect 11897 56493 11969 56545
rect 12021 56493 12093 56545
rect 12145 56493 12185 56545
rect 11185 56421 12185 56493
rect 11185 56369 11225 56421
rect 11277 56369 11349 56421
rect 11401 56369 11473 56421
rect 11525 56369 11597 56421
rect 11649 56369 11721 56421
rect 11773 56369 11845 56421
rect 11897 56369 11969 56421
rect 12021 56369 12093 56421
rect 12145 56369 12185 56421
rect 11185 56297 12185 56369
rect 11185 56245 11225 56297
rect 11277 56245 11349 56297
rect 11401 56245 11473 56297
rect 11525 56245 11597 56297
rect 11649 56245 11721 56297
rect 11773 56245 11845 56297
rect 11897 56245 11969 56297
rect 12021 56245 12093 56297
rect 12145 56245 12185 56297
rect 11185 56173 12185 56245
rect 11185 56121 11225 56173
rect 11277 56121 11349 56173
rect 11401 56121 11473 56173
rect 11525 56121 11597 56173
rect 11649 56121 11721 56173
rect 11773 56121 11845 56173
rect 11897 56121 11969 56173
rect 12021 56121 12093 56173
rect 12145 56121 12185 56173
rect 11185 56049 12185 56121
rect 11185 55997 11225 56049
rect 11277 55997 11349 56049
rect 11401 55997 11473 56049
rect 11525 55997 11597 56049
rect 11649 55997 11721 56049
rect 11773 55997 11845 56049
rect 11897 55997 11969 56049
rect 12021 55997 12093 56049
rect 12145 55997 12185 56049
rect 11185 55925 12185 55997
rect 11185 55873 11225 55925
rect 11277 55873 11349 55925
rect 11401 55873 11473 55925
rect 11525 55873 11597 55925
rect 11649 55873 11721 55925
rect 11773 55873 11845 55925
rect 11897 55873 11969 55925
rect 12021 55873 12093 55925
rect 12145 55873 12185 55925
rect 11185 55801 12185 55873
rect 11185 55749 11225 55801
rect 11277 55749 11349 55801
rect 11401 55749 11473 55801
rect 11525 55749 11597 55801
rect 11649 55749 11721 55801
rect 11773 55749 11845 55801
rect 11897 55749 11969 55801
rect 12021 55749 12093 55801
rect 12145 55749 12185 55801
rect 11185 55677 12185 55749
rect 11185 55625 11225 55677
rect 11277 55625 11349 55677
rect 11401 55625 11473 55677
rect 11525 55625 11597 55677
rect 11649 55625 11721 55677
rect 11773 55625 11845 55677
rect 11897 55625 11969 55677
rect 12021 55625 12093 55677
rect 12145 55625 12185 55677
rect 11185 55553 12185 55625
rect 11185 55501 11225 55553
rect 11277 55501 11349 55553
rect 11401 55501 11473 55553
rect 11525 55501 11597 55553
rect 11649 55501 11721 55553
rect 11773 55501 11845 55553
rect 11897 55501 11969 55553
rect 12021 55501 12093 55553
rect 12145 55501 12185 55553
rect 11185 55429 12185 55501
rect 11185 55377 11225 55429
rect 11277 55377 11349 55429
rect 11401 55377 11473 55429
rect 11525 55377 11597 55429
rect 11649 55377 11721 55429
rect 11773 55377 11845 55429
rect 11897 55377 11969 55429
rect 12021 55377 12093 55429
rect 12145 55377 12185 55429
rect 11185 55305 12185 55377
rect 11185 55253 11225 55305
rect 11277 55253 11349 55305
rect 11401 55253 11473 55305
rect 11525 55253 11597 55305
rect 11649 55253 11721 55305
rect 11773 55253 11845 55305
rect 11897 55253 11969 55305
rect 12021 55253 12093 55305
rect 12145 55253 12185 55305
rect 11185 55181 12185 55253
rect 11185 55129 11225 55181
rect 11277 55129 11349 55181
rect 11401 55129 11473 55181
rect 11525 55129 11597 55181
rect 11649 55129 11721 55181
rect 11773 55129 11845 55181
rect 11897 55129 11969 55181
rect 12021 55129 12093 55181
rect 12145 55129 12185 55181
rect 11185 55057 12185 55129
rect 11185 55005 11225 55057
rect 11277 55005 11349 55057
rect 11401 55005 11473 55057
rect 11525 55005 11597 55057
rect 11649 55005 11721 55057
rect 11773 55005 11845 55057
rect 11897 55005 11969 55057
rect 12021 55005 12093 55057
rect 12145 55005 12185 55057
rect 11185 54933 12185 55005
rect 11185 54881 11225 54933
rect 11277 54881 11349 54933
rect 11401 54881 11473 54933
rect 11525 54881 11597 54933
rect 11649 54881 11721 54933
rect 11773 54881 11845 54933
rect 11897 54881 11969 54933
rect 12021 54881 12093 54933
rect 12145 54881 12185 54933
rect 11185 54809 12185 54881
rect 11185 54757 11225 54809
rect 11277 54757 11349 54809
rect 11401 54757 11473 54809
rect 11525 54757 11597 54809
rect 11649 54757 11721 54809
rect 11773 54757 11845 54809
rect 11897 54757 11969 54809
rect 12021 54757 12093 54809
rect 12145 54757 12185 54809
rect 11185 54685 12185 54757
rect 11185 54633 11225 54685
rect 11277 54633 11349 54685
rect 11401 54633 11473 54685
rect 11525 54633 11597 54685
rect 11649 54633 11721 54685
rect 11773 54633 11845 54685
rect 11897 54633 11969 54685
rect 12021 54633 12093 54685
rect 12145 54633 12185 54685
rect 11185 54561 12185 54633
rect 11185 54509 11225 54561
rect 11277 54509 11349 54561
rect 11401 54509 11473 54561
rect 11525 54509 11597 54561
rect 11649 54509 11721 54561
rect 11773 54509 11845 54561
rect 11897 54509 11969 54561
rect 12021 54509 12093 54561
rect 12145 54509 12185 54561
rect 11185 54437 12185 54509
rect 11185 54385 11225 54437
rect 11277 54385 11349 54437
rect 11401 54385 11473 54437
rect 11525 54385 11597 54437
rect 11649 54385 11721 54437
rect 11773 54385 11845 54437
rect 11897 54385 11969 54437
rect 12021 54385 12093 54437
rect 12145 54385 12185 54437
rect 11185 54313 12185 54385
rect 11185 54261 11225 54313
rect 11277 54261 11349 54313
rect 11401 54261 11473 54313
rect 11525 54261 11597 54313
rect 11649 54261 11721 54313
rect 11773 54261 11845 54313
rect 11897 54261 11969 54313
rect 12021 54261 12093 54313
rect 12145 54261 12185 54313
rect 11185 54189 12185 54261
rect 11185 54137 11225 54189
rect 11277 54137 11349 54189
rect 11401 54137 11473 54189
rect 11525 54137 11597 54189
rect 11649 54137 11721 54189
rect 11773 54137 11845 54189
rect 11897 54137 11969 54189
rect 12021 54137 12093 54189
rect 12145 54137 12185 54189
rect 11185 54065 12185 54137
rect 11185 54013 11225 54065
rect 11277 54013 11349 54065
rect 11401 54013 11473 54065
rect 11525 54013 11597 54065
rect 11649 54013 11721 54065
rect 11773 54013 11845 54065
rect 11897 54013 11969 54065
rect 12021 54013 12093 54065
rect 12145 54013 12185 54065
rect 11185 53941 12185 54013
rect 11185 53889 11225 53941
rect 11277 53889 11349 53941
rect 11401 53889 11473 53941
rect 11525 53889 11597 53941
rect 11649 53889 11721 53941
rect 11773 53889 11845 53941
rect 11897 53889 11969 53941
rect 12021 53889 12093 53941
rect 12145 53889 12185 53941
rect 11185 53817 12185 53889
rect 11185 53765 11225 53817
rect 11277 53765 11349 53817
rect 11401 53765 11473 53817
rect 11525 53765 11597 53817
rect 11649 53765 11721 53817
rect 11773 53765 11845 53817
rect 11897 53765 11969 53817
rect 12021 53765 12093 53817
rect 12145 53765 12185 53817
rect 11185 53693 12185 53765
rect 11185 53641 11225 53693
rect 11277 53641 11349 53693
rect 11401 53641 11473 53693
rect 11525 53641 11597 53693
rect 11649 53641 11721 53693
rect 11773 53641 11845 53693
rect 11897 53641 11969 53693
rect 12021 53641 12093 53693
rect 12145 53641 12185 53693
rect 11185 53633 12185 53641
rect 13101 56669 14101 56677
rect 13101 56617 13141 56669
rect 13193 56617 13265 56669
rect 13317 56617 13389 56669
rect 13441 56617 13513 56669
rect 13565 56617 13637 56669
rect 13689 56617 13761 56669
rect 13813 56617 13885 56669
rect 13937 56617 14009 56669
rect 14061 56617 14101 56669
rect 14565 56655 14576 57048
rect 13101 56545 14101 56617
rect 13101 56493 13141 56545
rect 13193 56493 13265 56545
rect 13317 56493 13389 56545
rect 13441 56493 13513 56545
rect 13565 56493 13637 56545
rect 13689 56493 13761 56545
rect 13813 56493 13885 56545
rect 13937 56493 14009 56545
rect 14061 56493 14101 56545
rect 13101 56421 14101 56493
rect 13101 56369 13141 56421
rect 13193 56369 13265 56421
rect 13317 56369 13389 56421
rect 13441 56369 13513 56421
rect 13565 56369 13637 56421
rect 13689 56369 13761 56421
rect 13813 56369 13885 56421
rect 13937 56369 14009 56421
rect 14061 56369 14101 56421
rect 13101 56297 14101 56369
rect 13101 56245 13141 56297
rect 13193 56245 13265 56297
rect 13317 56245 13389 56297
rect 13441 56245 13513 56297
rect 13565 56245 13637 56297
rect 13689 56245 13761 56297
rect 13813 56245 13885 56297
rect 13937 56245 14009 56297
rect 14061 56245 14101 56297
rect 13101 56173 14101 56245
rect 13101 56121 13141 56173
rect 13193 56121 13265 56173
rect 13317 56121 13389 56173
rect 13441 56121 13513 56173
rect 13565 56121 13637 56173
rect 13689 56121 13761 56173
rect 13813 56121 13885 56173
rect 13937 56121 14009 56173
rect 14061 56121 14101 56173
rect 13101 56049 14101 56121
rect 13101 55997 13141 56049
rect 13193 55997 13265 56049
rect 13317 55997 13389 56049
rect 13441 55997 13513 56049
rect 13565 55997 13637 56049
rect 13689 55997 13761 56049
rect 13813 55997 13885 56049
rect 13937 55997 14009 56049
rect 14061 55997 14101 56049
rect 13101 55925 14101 55997
rect 13101 55873 13141 55925
rect 13193 55873 13265 55925
rect 13317 55873 13389 55925
rect 13441 55873 13513 55925
rect 13565 55873 13637 55925
rect 13689 55873 13761 55925
rect 13813 55873 13885 55925
rect 13937 55873 14009 55925
rect 14061 55873 14101 55925
rect 13101 55801 14101 55873
rect 13101 55749 13141 55801
rect 13193 55749 13265 55801
rect 13317 55749 13389 55801
rect 13441 55749 13513 55801
rect 13565 55749 13637 55801
rect 13689 55749 13761 55801
rect 13813 55749 13885 55801
rect 13937 55749 14009 55801
rect 14061 55749 14101 55801
rect 13101 55677 14101 55749
rect 13101 55625 13141 55677
rect 13193 55625 13265 55677
rect 13317 55625 13389 55677
rect 13441 55625 13513 55677
rect 13565 55625 13637 55677
rect 13689 55625 13761 55677
rect 13813 55625 13885 55677
rect 13937 55625 14009 55677
rect 14061 55625 14101 55677
rect 13101 55553 14101 55625
rect 13101 55501 13141 55553
rect 13193 55501 13265 55553
rect 13317 55501 13389 55553
rect 13441 55501 13513 55553
rect 13565 55501 13637 55553
rect 13689 55501 13761 55553
rect 13813 55501 13885 55553
rect 13937 55501 14009 55553
rect 14061 55501 14101 55553
rect 13101 55429 14101 55501
rect 13101 55377 13141 55429
rect 13193 55377 13265 55429
rect 13317 55377 13389 55429
rect 13441 55377 13513 55429
rect 13565 55377 13637 55429
rect 13689 55377 13761 55429
rect 13813 55377 13885 55429
rect 13937 55377 14009 55429
rect 14061 55377 14101 55429
rect 13101 55305 14101 55377
rect 13101 55253 13141 55305
rect 13193 55253 13265 55305
rect 13317 55253 13389 55305
rect 13441 55253 13513 55305
rect 13565 55253 13637 55305
rect 13689 55253 13761 55305
rect 13813 55253 13885 55305
rect 13937 55253 14009 55305
rect 14061 55253 14101 55305
rect 13101 55181 14101 55253
rect 13101 55129 13141 55181
rect 13193 55129 13265 55181
rect 13317 55129 13389 55181
rect 13441 55129 13513 55181
rect 13565 55129 13637 55181
rect 13689 55129 13761 55181
rect 13813 55129 13885 55181
rect 13937 55129 14009 55181
rect 14061 55129 14101 55181
rect 13101 55057 14101 55129
rect 13101 55005 13141 55057
rect 13193 55005 13265 55057
rect 13317 55005 13389 55057
rect 13441 55005 13513 55057
rect 13565 55005 13637 55057
rect 13689 55005 13761 55057
rect 13813 55005 13885 55057
rect 13937 55005 14009 55057
rect 14061 55005 14101 55057
rect 13101 54933 14101 55005
rect 13101 54881 13141 54933
rect 13193 54881 13265 54933
rect 13317 54881 13389 54933
rect 13441 54881 13513 54933
rect 13565 54881 13637 54933
rect 13689 54881 13761 54933
rect 13813 54881 13885 54933
rect 13937 54881 14009 54933
rect 14061 54881 14101 54933
rect 13101 54809 14101 54881
rect 13101 54757 13141 54809
rect 13193 54757 13265 54809
rect 13317 54757 13389 54809
rect 13441 54757 13513 54809
rect 13565 54757 13637 54809
rect 13689 54757 13761 54809
rect 13813 54757 13885 54809
rect 13937 54757 14009 54809
rect 14061 54757 14101 54809
rect 13101 54685 14101 54757
rect 13101 54633 13141 54685
rect 13193 54633 13265 54685
rect 13317 54633 13389 54685
rect 13441 54633 13513 54685
rect 13565 54633 13637 54685
rect 13689 54633 13761 54685
rect 13813 54633 13885 54685
rect 13937 54633 14009 54685
rect 14061 54633 14101 54685
rect 13101 54561 14101 54633
rect 13101 54509 13141 54561
rect 13193 54509 13265 54561
rect 13317 54509 13389 54561
rect 13441 54509 13513 54561
rect 13565 54509 13637 54561
rect 13689 54509 13761 54561
rect 13813 54509 13885 54561
rect 13937 54509 14009 54561
rect 14061 54509 14101 54561
rect 13101 54437 14101 54509
rect 13101 54385 13141 54437
rect 13193 54385 13265 54437
rect 13317 54385 13389 54437
rect 13441 54385 13513 54437
rect 13565 54385 13637 54437
rect 13689 54385 13761 54437
rect 13813 54385 13885 54437
rect 13937 54385 14009 54437
rect 14061 54385 14101 54437
rect 13101 54313 14101 54385
rect 13101 54261 13141 54313
rect 13193 54261 13265 54313
rect 13317 54261 13389 54313
rect 13441 54261 13513 54313
rect 13565 54261 13637 54313
rect 13689 54261 13761 54313
rect 13813 54261 13885 54313
rect 13937 54261 14009 54313
rect 14061 54261 14101 54313
rect 13101 54189 14101 54261
rect 13101 54137 13141 54189
rect 13193 54137 13265 54189
rect 13317 54137 13389 54189
rect 13441 54137 13513 54189
rect 13565 54137 13637 54189
rect 13689 54137 13761 54189
rect 13813 54137 13885 54189
rect 13937 54137 14009 54189
rect 14061 54137 14101 54189
rect 13101 54065 14101 54137
rect 13101 54013 13141 54065
rect 13193 54013 13265 54065
rect 13317 54013 13389 54065
rect 13441 54013 13513 54065
rect 13565 54013 13637 54065
rect 13689 54013 13761 54065
rect 13813 54013 13885 54065
rect 13937 54013 14009 54065
rect 14061 54013 14101 54065
rect 13101 53941 14101 54013
rect 13101 53889 13141 53941
rect 13193 53889 13265 53941
rect 13317 53889 13389 53941
rect 13441 53889 13513 53941
rect 13565 53889 13637 53941
rect 13689 53889 13761 53941
rect 13813 53889 13885 53941
rect 13937 53889 14009 53941
rect 14061 53889 14101 53941
rect 13101 53817 14101 53889
rect 13101 53765 13141 53817
rect 13193 53765 13265 53817
rect 13317 53765 13389 53817
rect 13441 53765 13513 53817
rect 13565 53765 13637 53817
rect 13689 53765 13761 53817
rect 13813 53765 13885 53817
rect 13937 53765 14009 53817
rect 14061 53765 14101 53817
rect 13101 53693 14101 53765
rect 13101 53641 13141 53693
rect 13193 53641 13265 53693
rect 13317 53641 13389 53693
rect 13441 53641 13513 53693
rect 13565 53641 13637 53693
rect 13689 53641 13761 53693
rect 13813 53641 13885 53693
rect 13937 53641 14009 53693
rect 14061 53641 14101 53693
rect 13101 53633 14101 53641
rect 11185 53622 14101 53633
rect 11185 53576 11196 53622
rect 14090 53576 14101 53622
rect 11185 53565 14101 53576
rect 14161 56618 14576 56655
rect 14161 53692 14172 56618
rect 14218 53692 14576 56618
rect 14161 53505 14576 53692
rect 402 53484 14576 53505
rect 402 53432 2501 53484
rect 2553 53432 2609 53484
rect 2661 53432 4871 53484
rect 4923 53432 4979 53484
rect 5031 53432 7247 53484
rect 7299 53432 7355 53484
rect 7407 53432 7463 53484
rect 7515 53432 7571 53484
rect 7623 53432 7679 53484
rect 7731 53432 9947 53484
rect 9999 53432 10055 53484
rect 10107 53432 12317 53484
rect 12369 53432 12425 53484
rect 12477 53432 14576 53484
rect 402 53376 14576 53432
rect 402 53324 2501 53376
rect 2553 53324 2609 53376
rect 2661 53324 4871 53376
rect 4923 53324 4979 53376
rect 5031 53324 7247 53376
rect 7299 53324 7355 53376
rect 7407 53324 7463 53376
rect 7515 53324 7571 53376
rect 7623 53324 7679 53376
rect 7731 53324 9947 53376
rect 9999 53324 10055 53376
rect 10107 53324 12317 53376
rect 12369 53324 12425 53376
rect 12477 53324 14576 53376
rect 402 53268 14576 53324
rect 402 53251 2501 53268
rect 2553 53251 2609 53268
rect 2661 53251 4871 53268
rect 4923 53251 4979 53268
rect 5031 53251 7247 53268
rect 7299 53251 7355 53268
rect 7407 53251 7463 53268
rect 7515 53251 7571 53268
rect 7623 53251 7679 53268
rect 7731 53251 9947 53268
rect 9999 53251 10055 53268
rect 10107 53251 12317 53268
rect 12369 53251 12425 53268
rect 12477 53251 14576 53268
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14633 57105
rect 345 53194 14633 53205
rect 71 52611 2225 52622
rect 71 52586 268 52611
rect 10 52574 268 52586
rect 10 52522 22 52574
rect 74 52522 268 52574
rect 10 52466 268 52522
rect 10 52414 22 52466
rect 74 52414 268 52466
rect 10 52358 268 52414
rect 10 52306 22 52358
rect 74 52306 268 52358
rect 10 52250 268 52306
rect 10 52198 22 52250
rect 74 52198 268 52250
rect 10 52142 268 52198
rect 10 52090 22 52142
rect 74 52090 268 52142
rect 10 52034 268 52090
rect 10 51982 22 52034
rect 74 51982 268 52034
rect 10 51926 268 51982
rect 10 51874 22 51926
rect 74 51874 268 51926
rect 10 51818 268 51874
rect 10 51766 22 51818
rect 74 51766 268 51818
rect 10 51710 268 51766
rect 10 51658 22 51710
rect 74 51658 268 51710
rect 10 51622 268 51658
rect 10 51602 86 51622
rect 10 51550 22 51602
rect 74 51550 86 51602
rect 10 51494 86 51550
rect 10 51442 22 51494
rect 74 51442 86 51494
rect 10 51422 86 51442
rect 257 51422 268 51622
rect 10 51386 268 51422
rect 10 51334 22 51386
rect 74 51334 268 51386
rect 10 51278 268 51334
rect 10 51226 22 51278
rect 74 51226 268 51278
rect 10 51214 268 51226
rect 71 50422 268 51214
rect 257 49854 268 50422
rect 71 48854 268 49854
rect 257 48654 268 48854
rect 71 47665 268 48654
rect 2214 47665 2225 52611
rect 71 47654 2225 47665
rect 2551 52611 12427 52622
rect 2551 47665 2562 52611
rect 2908 52588 3016 52611
rect 11962 52588 12070 52611
rect 2908 52536 2934 52588
rect 2986 52536 3016 52588
rect 11962 52536 11992 52588
rect 12044 52536 12070 52588
rect 2908 52464 3016 52536
rect 11962 52464 12070 52536
rect 2908 52412 2934 52464
rect 2986 52412 3016 52464
rect 11962 52412 11992 52464
rect 12044 52412 12070 52464
rect 2908 52340 3016 52412
rect 11962 52340 12070 52412
rect 2908 52288 2934 52340
rect 2986 52288 3016 52340
rect 11962 52288 11992 52340
rect 12044 52288 12070 52340
rect 2908 52265 3016 52288
rect 11962 52265 12070 52288
rect 2908 52254 12070 52265
rect 2908 48022 2919 52254
rect 3105 52029 11873 52040
rect 3105 51983 3142 52029
rect 11836 51983 11873 52029
rect 3105 51965 4863 51983
rect 4915 51965 4987 51983
rect 5039 51965 7277 51983
rect 7329 51965 7401 51983
rect 7453 51965 7525 51983
rect 7577 51965 7649 51983
rect 7701 51965 9939 51983
rect 9991 51965 10063 51983
rect 10115 51965 11873 51983
rect 3105 51900 11873 51965
rect 3105 48376 3116 51900
rect 3162 51893 11816 51900
rect 3162 51875 4863 51893
rect 4915 51875 4987 51893
rect 5039 51875 7277 51893
rect 7329 51875 7401 51893
rect 7453 51875 7525 51893
rect 7577 51875 7649 51893
rect 7701 51875 9939 51893
rect 9991 51875 10063 51893
rect 10115 51875 11816 51893
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51818 11662 51829
rect 3316 51260 3327 51818
rect 3489 51627 11489 51639
rect 3489 51626 3559 51627
rect 3611 51626 3683 51627
rect 3735 51626 3807 51627
rect 3859 51626 3931 51627
rect 3983 51626 4055 51627
rect 4107 51626 4179 51627
rect 4231 51626 4303 51627
rect 4355 51626 4427 51627
rect 4479 51626 4551 51627
rect 4603 51626 4675 51627
rect 4727 51626 5180 51627
rect 5232 51626 5304 51627
rect 5356 51626 5428 51627
rect 5480 51626 5552 51627
rect 5604 51626 5676 51627
rect 5728 51626 5800 51627
rect 5852 51626 5924 51627
rect 5976 51626 6048 51627
rect 6100 51626 6172 51627
rect 6224 51626 6296 51627
rect 6348 51626 6420 51627
rect 6472 51626 6544 51627
rect 6596 51626 6668 51627
rect 6720 51626 6792 51627
rect 6844 51626 6916 51627
rect 6968 51626 7040 51627
rect 7092 51626 7886 51627
rect 7938 51626 8010 51627
rect 8062 51626 8134 51627
rect 8186 51626 8258 51627
rect 8310 51626 8382 51627
rect 8434 51626 8506 51627
rect 8558 51626 8630 51627
rect 8682 51626 8754 51627
rect 8806 51626 8878 51627
rect 8930 51626 9002 51627
rect 9054 51626 9126 51627
rect 9178 51626 9250 51627
rect 9302 51626 9374 51627
rect 9426 51626 9498 51627
rect 9550 51626 9622 51627
rect 9674 51626 9746 51627
rect 9798 51626 10251 51627
rect 10303 51626 10375 51627
rect 10427 51626 10499 51627
rect 10551 51626 10623 51627
rect 10675 51626 10747 51627
rect 10799 51626 10871 51627
rect 10923 51626 10995 51627
rect 11047 51626 11119 51627
rect 11171 51626 11243 51627
rect 11295 51626 11367 51627
rect 11419 51626 11489 51627
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51575 3559 51580
rect 3611 51575 3683 51580
rect 3735 51575 3807 51580
rect 3859 51575 3931 51580
rect 3983 51575 4055 51580
rect 4107 51575 4179 51580
rect 4231 51575 4303 51580
rect 4355 51575 4427 51580
rect 4479 51575 4551 51580
rect 4603 51575 4675 51580
rect 4727 51575 5180 51580
rect 5232 51575 5304 51580
rect 5356 51575 5428 51580
rect 5480 51575 5552 51580
rect 5604 51575 5676 51580
rect 5728 51575 5800 51580
rect 5852 51575 5924 51580
rect 5976 51575 6048 51580
rect 6100 51575 6172 51580
rect 6224 51575 6296 51580
rect 6348 51575 6420 51580
rect 6472 51575 6544 51580
rect 6596 51575 6668 51580
rect 6720 51575 6792 51580
rect 6844 51575 6916 51580
rect 6968 51575 7040 51580
rect 7092 51575 7886 51580
rect 7938 51575 8010 51580
rect 8062 51575 8134 51580
rect 8186 51575 8258 51580
rect 8310 51575 8382 51580
rect 8434 51575 8506 51580
rect 8558 51575 8630 51580
rect 8682 51575 8754 51580
rect 8806 51575 8878 51580
rect 8930 51575 9002 51580
rect 9054 51575 9126 51580
rect 9178 51575 9250 51580
rect 9302 51575 9374 51580
rect 9426 51575 9498 51580
rect 9550 51575 9622 51580
rect 9674 51575 9746 51580
rect 9798 51575 10251 51580
rect 10303 51575 10375 51580
rect 10427 51575 10499 51580
rect 10551 51575 10623 51580
rect 10675 51575 10747 51580
rect 10799 51575 10871 51580
rect 10923 51575 10995 51580
rect 11047 51575 11119 51580
rect 11171 51575 11243 51580
rect 11295 51575 11367 51580
rect 11419 51575 11489 51580
rect 3489 51503 11489 51575
rect 3489 51498 3559 51503
rect 3611 51498 3683 51503
rect 3735 51498 3807 51503
rect 3859 51498 3931 51503
rect 3983 51498 4055 51503
rect 4107 51498 4179 51503
rect 4231 51498 4303 51503
rect 4355 51498 4427 51503
rect 4479 51498 4551 51503
rect 4603 51498 4675 51503
rect 4727 51498 5180 51503
rect 5232 51498 5304 51503
rect 5356 51498 5428 51503
rect 5480 51498 5552 51503
rect 5604 51498 5676 51503
rect 5728 51498 5800 51503
rect 5852 51498 5924 51503
rect 5976 51498 6048 51503
rect 6100 51498 6172 51503
rect 6224 51498 6296 51503
rect 6348 51498 6420 51503
rect 6472 51498 6544 51503
rect 6596 51498 6668 51503
rect 6720 51498 6792 51503
rect 6844 51498 6916 51503
rect 6968 51498 7040 51503
rect 7092 51498 7886 51503
rect 7938 51498 8010 51503
rect 8062 51498 8134 51503
rect 8186 51498 8258 51503
rect 8310 51498 8382 51503
rect 8434 51498 8506 51503
rect 8558 51498 8630 51503
rect 8682 51498 8754 51503
rect 8806 51498 8878 51503
rect 8930 51498 9002 51503
rect 9054 51498 9126 51503
rect 9178 51498 9250 51503
rect 9302 51498 9374 51503
rect 9426 51498 9498 51503
rect 9550 51498 9622 51503
rect 9674 51498 9746 51503
rect 9798 51498 10251 51503
rect 10303 51498 10375 51503
rect 10427 51498 10499 51503
rect 10551 51498 10623 51503
rect 10675 51498 10747 51503
rect 10799 51498 10871 51503
rect 10923 51498 10995 51503
rect 11047 51498 11119 51503
rect 11171 51498 11243 51503
rect 11295 51498 11367 51503
rect 11419 51498 11489 51503
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51451 3559 51452
rect 3611 51451 3683 51452
rect 3735 51451 3807 51452
rect 3859 51451 3931 51452
rect 3983 51451 4055 51452
rect 4107 51451 4179 51452
rect 4231 51451 4303 51452
rect 4355 51451 4427 51452
rect 4479 51451 4551 51452
rect 4603 51451 4675 51452
rect 4727 51451 5180 51452
rect 5232 51451 5304 51452
rect 5356 51451 5428 51452
rect 5480 51451 5552 51452
rect 5604 51451 5676 51452
rect 5728 51451 5800 51452
rect 5852 51451 5924 51452
rect 5976 51451 6048 51452
rect 6100 51451 6172 51452
rect 6224 51451 6296 51452
rect 6348 51451 6420 51452
rect 6472 51451 6544 51452
rect 6596 51451 6668 51452
rect 6720 51451 6792 51452
rect 6844 51451 6916 51452
rect 6968 51451 7040 51452
rect 7092 51451 7886 51452
rect 7938 51451 8010 51452
rect 8062 51451 8134 51452
rect 8186 51451 8258 51452
rect 8310 51451 8382 51452
rect 8434 51451 8506 51452
rect 8558 51451 8630 51452
rect 8682 51451 8754 51452
rect 8806 51451 8878 51452
rect 8930 51451 9002 51452
rect 9054 51451 9126 51452
rect 9178 51451 9250 51452
rect 9302 51451 9374 51452
rect 9426 51451 9498 51452
rect 9550 51451 9622 51452
rect 9674 51451 9746 51452
rect 9798 51451 10251 51452
rect 10303 51451 10375 51452
rect 10427 51451 10499 51452
rect 10551 51451 10623 51452
rect 10675 51451 10747 51452
rect 10799 51451 10871 51452
rect 10923 51451 10995 51452
rect 11047 51451 11119 51452
rect 11171 51451 11243 51452
rect 11295 51451 11367 51452
rect 11419 51451 11489 51452
rect 3489 51439 11489 51451
rect 11651 51260 11662 51818
rect 3316 51249 11662 51260
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51170 4863 51203
rect 4915 51170 4987 51203
rect 5039 51170 7277 51203
rect 7329 51170 7401 51203
rect 7453 51170 7525 51203
rect 7577 51170 7649 51203
rect 7701 51170 9939 51203
rect 9991 51170 10063 51203
rect 10115 51170 11816 51203
rect 3162 51098 11816 51170
rect 3162 51095 4863 51098
rect 4915 51095 4987 51098
rect 5039 51095 7277 51098
rect 7329 51095 7401 51098
rect 7453 51095 7525 51098
rect 7577 51095 7649 51098
rect 7701 51095 9939 51098
rect 9991 51095 10063 51098
rect 10115 51095 11816 51098
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 51046 4863 51049
rect 4915 51046 4987 51049
rect 5039 51046 7277 51049
rect 7329 51046 7401 51049
rect 7453 51046 7525 51049
rect 7577 51046 7649 51049
rect 7701 51046 9939 51049
rect 9991 51046 10063 51049
rect 10115 51046 11816 51049
rect 3162 50974 11816 51046
rect 3162 50941 4863 50974
rect 4915 50941 4987 50974
rect 5039 50941 7277 50974
rect 7329 50941 7401 50974
rect 7453 50941 7525 50974
rect 7577 50941 7649 50974
rect 7701 50941 9939 50974
rect 9991 50941 10063 50974
rect 10115 50941 11816 50974
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50884 11662 50895
rect 3316 50326 3327 50884
rect 3489 50693 11489 50705
rect 3489 50692 3559 50693
rect 3611 50692 3683 50693
rect 3735 50692 3807 50693
rect 3859 50692 3931 50693
rect 3983 50692 4055 50693
rect 4107 50692 4179 50693
rect 4231 50692 4303 50693
rect 4355 50692 4427 50693
rect 4479 50692 4551 50693
rect 4603 50692 4675 50693
rect 4727 50692 5180 50693
rect 5232 50692 5304 50693
rect 5356 50692 5428 50693
rect 5480 50692 5552 50693
rect 5604 50692 5676 50693
rect 5728 50692 5800 50693
rect 5852 50692 5924 50693
rect 5976 50692 6048 50693
rect 6100 50692 6172 50693
rect 6224 50692 6296 50693
rect 6348 50692 6420 50693
rect 6472 50692 6544 50693
rect 6596 50692 6668 50693
rect 6720 50692 6792 50693
rect 6844 50692 6916 50693
rect 6968 50692 7040 50693
rect 7092 50692 7886 50693
rect 7938 50692 8010 50693
rect 8062 50692 8134 50693
rect 8186 50692 8258 50693
rect 8310 50692 8382 50693
rect 8434 50692 8506 50693
rect 8558 50692 8630 50693
rect 8682 50692 8754 50693
rect 8806 50692 8878 50693
rect 8930 50692 9002 50693
rect 9054 50692 9126 50693
rect 9178 50692 9250 50693
rect 9302 50692 9374 50693
rect 9426 50692 9498 50693
rect 9550 50692 9622 50693
rect 9674 50692 9746 50693
rect 9798 50692 10251 50693
rect 10303 50692 10375 50693
rect 10427 50692 10499 50693
rect 10551 50692 10623 50693
rect 10675 50692 10747 50693
rect 10799 50692 10871 50693
rect 10923 50692 10995 50693
rect 11047 50692 11119 50693
rect 11171 50692 11243 50693
rect 11295 50692 11367 50693
rect 11419 50692 11489 50693
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50641 3559 50646
rect 3611 50641 3683 50646
rect 3735 50641 3807 50646
rect 3859 50641 3931 50646
rect 3983 50641 4055 50646
rect 4107 50641 4179 50646
rect 4231 50641 4303 50646
rect 4355 50641 4427 50646
rect 4479 50641 4551 50646
rect 4603 50641 4675 50646
rect 4727 50641 5180 50646
rect 5232 50641 5304 50646
rect 5356 50641 5428 50646
rect 5480 50641 5552 50646
rect 5604 50641 5676 50646
rect 5728 50641 5800 50646
rect 5852 50641 5924 50646
rect 5976 50641 6048 50646
rect 6100 50641 6172 50646
rect 6224 50641 6296 50646
rect 6348 50641 6420 50646
rect 6472 50641 6544 50646
rect 6596 50641 6668 50646
rect 6720 50641 6792 50646
rect 6844 50641 6916 50646
rect 6968 50641 7040 50646
rect 7092 50641 7886 50646
rect 7938 50641 8010 50646
rect 8062 50641 8134 50646
rect 8186 50641 8258 50646
rect 8310 50641 8382 50646
rect 8434 50641 8506 50646
rect 8558 50641 8630 50646
rect 8682 50641 8754 50646
rect 8806 50641 8878 50646
rect 8930 50641 9002 50646
rect 9054 50641 9126 50646
rect 9178 50641 9250 50646
rect 9302 50641 9374 50646
rect 9426 50641 9498 50646
rect 9550 50641 9622 50646
rect 9674 50641 9746 50646
rect 9798 50641 10251 50646
rect 10303 50641 10375 50646
rect 10427 50641 10499 50646
rect 10551 50641 10623 50646
rect 10675 50641 10747 50646
rect 10799 50641 10871 50646
rect 10923 50641 10995 50646
rect 11047 50641 11119 50646
rect 11171 50641 11243 50646
rect 11295 50641 11367 50646
rect 11419 50641 11489 50646
rect 3489 50569 11489 50641
rect 3489 50564 3559 50569
rect 3611 50564 3683 50569
rect 3735 50564 3807 50569
rect 3859 50564 3931 50569
rect 3983 50564 4055 50569
rect 4107 50564 4179 50569
rect 4231 50564 4303 50569
rect 4355 50564 4427 50569
rect 4479 50564 4551 50569
rect 4603 50564 4675 50569
rect 4727 50564 5180 50569
rect 5232 50564 5304 50569
rect 5356 50564 5428 50569
rect 5480 50564 5552 50569
rect 5604 50564 5676 50569
rect 5728 50564 5800 50569
rect 5852 50564 5924 50569
rect 5976 50564 6048 50569
rect 6100 50564 6172 50569
rect 6224 50564 6296 50569
rect 6348 50564 6420 50569
rect 6472 50564 6544 50569
rect 6596 50564 6668 50569
rect 6720 50564 6792 50569
rect 6844 50564 6916 50569
rect 6968 50564 7040 50569
rect 7092 50564 7886 50569
rect 7938 50564 8010 50569
rect 8062 50564 8134 50569
rect 8186 50564 8258 50569
rect 8310 50564 8382 50569
rect 8434 50564 8506 50569
rect 8558 50564 8630 50569
rect 8682 50564 8754 50569
rect 8806 50564 8878 50569
rect 8930 50564 9002 50569
rect 9054 50564 9126 50569
rect 9178 50564 9250 50569
rect 9302 50564 9374 50569
rect 9426 50564 9498 50569
rect 9550 50564 9622 50569
rect 9674 50564 9746 50569
rect 9798 50564 10251 50569
rect 10303 50564 10375 50569
rect 10427 50564 10499 50569
rect 10551 50564 10623 50569
rect 10675 50564 10747 50569
rect 10799 50564 10871 50569
rect 10923 50564 10995 50569
rect 11047 50564 11119 50569
rect 11171 50564 11243 50569
rect 11295 50564 11367 50569
rect 11419 50564 11489 50569
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50517 3559 50518
rect 3611 50517 3683 50518
rect 3735 50517 3807 50518
rect 3859 50517 3931 50518
rect 3983 50517 4055 50518
rect 4107 50517 4179 50518
rect 4231 50517 4303 50518
rect 4355 50517 4427 50518
rect 4479 50517 4551 50518
rect 4603 50517 4675 50518
rect 4727 50517 5180 50518
rect 5232 50517 5304 50518
rect 5356 50517 5428 50518
rect 5480 50517 5552 50518
rect 5604 50517 5676 50518
rect 5728 50517 5800 50518
rect 5852 50517 5924 50518
rect 5976 50517 6048 50518
rect 6100 50517 6172 50518
rect 6224 50517 6296 50518
rect 6348 50517 6420 50518
rect 6472 50517 6544 50518
rect 6596 50517 6668 50518
rect 6720 50517 6792 50518
rect 6844 50517 6916 50518
rect 6968 50517 7040 50518
rect 7092 50517 7886 50518
rect 7938 50517 8010 50518
rect 8062 50517 8134 50518
rect 8186 50517 8258 50518
rect 8310 50517 8382 50518
rect 8434 50517 8506 50518
rect 8558 50517 8630 50518
rect 8682 50517 8754 50518
rect 8806 50517 8878 50518
rect 8930 50517 9002 50518
rect 9054 50517 9126 50518
rect 9178 50517 9250 50518
rect 9302 50517 9374 50518
rect 9426 50517 9498 50518
rect 9550 50517 9622 50518
rect 9674 50517 9746 50518
rect 9798 50517 10251 50518
rect 10303 50517 10375 50518
rect 10427 50517 10499 50518
rect 10551 50517 10623 50518
rect 10675 50517 10747 50518
rect 10799 50517 10871 50518
rect 10923 50517 10995 50518
rect 11047 50517 11119 50518
rect 11171 50517 11243 50518
rect 11295 50517 11367 50518
rect 11419 50517 11489 50518
rect 3489 50505 11489 50517
rect 11651 50326 11662 50884
rect 3316 50315 11662 50326
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50236 4863 50269
rect 4915 50236 4987 50269
rect 5039 50236 7277 50269
rect 7329 50236 7401 50269
rect 7453 50236 7525 50269
rect 7577 50236 7649 50269
rect 7701 50236 9939 50269
rect 9991 50236 10063 50269
rect 10115 50236 11816 50269
rect 3162 50164 11816 50236
rect 3162 50161 4863 50164
rect 4915 50161 4987 50164
rect 5039 50161 7277 50164
rect 7329 50161 7401 50164
rect 7453 50161 7525 50164
rect 7577 50161 7649 50164
rect 7701 50161 9939 50164
rect 9991 50161 10063 50164
rect 10115 50161 11816 50164
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50112 4863 50115
rect 4915 50112 4987 50115
rect 5039 50112 7277 50115
rect 7329 50112 7401 50115
rect 7453 50112 7525 50115
rect 7577 50112 7649 50115
rect 7701 50112 9939 50115
rect 9991 50112 10063 50115
rect 10115 50112 11816 50115
rect 3162 50040 11816 50112
rect 3162 50007 4863 50040
rect 4915 50007 4987 50040
rect 5039 50007 7277 50040
rect 7329 50007 7401 50040
rect 7453 50007 7525 50040
rect 7577 50007 7649 50040
rect 7701 50007 9939 50040
rect 9991 50007 10063 50040
rect 10115 50007 11816 50040
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49950 11662 49961
rect 3316 49392 3327 49950
rect 3489 49759 11489 49771
rect 3489 49758 3559 49759
rect 3611 49758 3683 49759
rect 3735 49758 3807 49759
rect 3859 49758 3931 49759
rect 3983 49758 4055 49759
rect 4107 49758 4179 49759
rect 4231 49758 4303 49759
rect 4355 49758 4427 49759
rect 4479 49758 4551 49759
rect 4603 49758 4675 49759
rect 4727 49758 5180 49759
rect 5232 49758 5304 49759
rect 5356 49758 5428 49759
rect 5480 49758 5552 49759
rect 5604 49758 5676 49759
rect 5728 49758 5800 49759
rect 5852 49758 5924 49759
rect 5976 49758 6048 49759
rect 6100 49758 6172 49759
rect 6224 49758 6296 49759
rect 6348 49758 6420 49759
rect 6472 49758 6544 49759
rect 6596 49758 6668 49759
rect 6720 49758 6792 49759
rect 6844 49758 6916 49759
rect 6968 49758 7040 49759
rect 7092 49758 7886 49759
rect 7938 49758 8010 49759
rect 8062 49758 8134 49759
rect 8186 49758 8258 49759
rect 8310 49758 8382 49759
rect 8434 49758 8506 49759
rect 8558 49758 8630 49759
rect 8682 49758 8754 49759
rect 8806 49758 8878 49759
rect 8930 49758 9002 49759
rect 9054 49758 9126 49759
rect 9178 49758 9250 49759
rect 9302 49758 9374 49759
rect 9426 49758 9498 49759
rect 9550 49758 9622 49759
rect 9674 49758 9746 49759
rect 9798 49758 10251 49759
rect 10303 49758 10375 49759
rect 10427 49758 10499 49759
rect 10551 49758 10623 49759
rect 10675 49758 10747 49759
rect 10799 49758 10871 49759
rect 10923 49758 10995 49759
rect 11047 49758 11119 49759
rect 11171 49758 11243 49759
rect 11295 49758 11367 49759
rect 11419 49758 11489 49759
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49707 3559 49712
rect 3611 49707 3683 49712
rect 3735 49707 3807 49712
rect 3859 49707 3931 49712
rect 3983 49707 4055 49712
rect 4107 49707 4179 49712
rect 4231 49707 4303 49712
rect 4355 49707 4427 49712
rect 4479 49707 4551 49712
rect 4603 49707 4675 49712
rect 4727 49707 5180 49712
rect 5232 49707 5304 49712
rect 5356 49707 5428 49712
rect 5480 49707 5552 49712
rect 5604 49707 5676 49712
rect 5728 49707 5800 49712
rect 5852 49707 5924 49712
rect 5976 49707 6048 49712
rect 6100 49707 6172 49712
rect 6224 49707 6296 49712
rect 6348 49707 6420 49712
rect 6472 49707 6544 49712
rect 6596 49707 6668 49712
rect 6720 49707 6792 49712
rect 6844 49707 6916 49712
rect 6968 49707 7040 49712
rect 7092 49707 7886 49712
rect 7938 49707 8010 49712
rect 8062 49707 8134 49712
rect 8186 49707 8258 49712
rect 8310 49707 8382 49712
rect 8434 49707 8506 49712
rect 8558 49707 8630 49712
rect 8682 49707 8754 49712
rect 8806 49707 8878 49712
rect 8930 49707 9002 49712
rect 9054 49707 9126 49712
rect 9178 49707 9250 49712
rect 9302 49707 9374 49712
rect 9426 49707 9498 49712
rect 9550 49707 9622 49712
rect 9674 49707 9746 49712
rect 9798 49707 10251 49712
rect 10303 49707 10375 49712
rect 10427 49707 10499 49712
rect 10551 49707 10623 49712
rect 10675 49707 10747 49712
rect 10799 49707 10871 49712
rect 10923 49707 10995 49712
rect 11047 49707 11119 49712
rect 11171 49707 11243 49712
rect 11295 49707 11367 49712
rect 11419 49707 11489 49712
rect 3489 49635 11489 49707
rect 3489 49630 3559 49635
rect 3611 49630 3683 49635
rect 3735 49630 3807 49635
rect 3859 49630 3931 49635
rect 3983 49630 4055 49635
rect 4107 49630 4179 49635
rect 4231 49630 4303 49635
rect 4355 49630 4427 49635
rect 4479 49630 4551 49635
rect 4603 49630 4675 49635
rect 4727 49630 5180 49635
rect 5232 49630 5304 49635
rect 5356 49630 5428 49635
rect 5480 49630 5552 49635
rect 5604 49630 5676 49635
rect 5728 49630 5800 49635
rect 5852 49630 5924 49635
rect 5976 49630 6048 49635
rect 6100 49630 6172 49635
rect 6224 49630 6296 49635
rect 6348 49630 6420 49635
rect 6472 49630 6544 49635
rect 6596 49630 6668 49635
rect 6720 49630 6792 49635
rect 6844 49630 6916 49635
rect 6968 49630 7040 49635
rect 7092 49630 7886 49635
rect 7938 49630 8010 49635
rect 8062 49630 8134 49635
rect 8186 49630 8258 49635
rect 8310 49630 8382 49635
rect 8434 49630 8506 49635
rect 8558 49630 8630 49635
rect 8682 49630 8754 49635
rect 8806 49630 8878 49635
rect 8930 49630 9002 49635
rect 9054 49630 9126 49635
rect 9178 49630 9250 49635
rect 9302 49630 9374 49635
rect 9426 49630 9498 49635
rect 9550 49630 9622 49635
rect 9674 49630 9746 49635
rect 9798 49630 10251 49635
rect 10303 49630 10375 49635
rect 10427 49630 10499 49635
rect 10551 49630 10623 49635
rect 10675 49630 10747 49635
rect 10799 49630 10871 49635
rect 10923 49630 10995 49635
rect 11047 49630 11119 49635
rect 11171 49630 11243 49635
rect 11295 49630 11367 49635
rect 11419 49630 11489 49635
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49583 3559 49584
rect 3611 49583 3683 49584
rect 3735 49583 3807 49584
rect 3859 49583 3931 49584
rect 3983 49583 4055 49584
rect 4107 49583 4179 49584
rect 4231 49583 4303 49584
rect 4355 49583 4427 49584
rect 4479 49583 4551 49584
rect 4603 49583 4675 49584
rect 4727 49583 5180 49584
rect 5232 49583 5304 49584
rect 5356 49583 5428 49584
rect 5480 49583 5552 49584
rect 5604 49583 5676 49584
rect 5728 49583 5800 49584
rect 5852 49583 5924 49584
rect 5976 49583 6048 49584
rect 6100 49583 6172 49584
rect 6224 49583 6296 49584
rect 6348 49583 6420 49584
rect 6472 49583 6544 49584
rect 6596 49583 6668 49584
rect 6720 49583 6792 49584
rect 6844 49583 6916 49584
rect 6968 49583 7040 49584
rect 7092 49583 7886 49584
rect 7938 49583 8010 49584
rect 8062 49583 8134 49584
rect 8186 49583 8258 49584
rect 8310 49583 8382 49584
rect 8434 49583 8506 49584
rect 8558 49583 8630 49584
rect 8682 49583 8754 49584
rect 8806 49583 8878 49584
rect 8930 49583 9002 49584
rect 9054 49583 9126 49584
rect 9178 49583 9250 49584
rect 9302 49583 9374 49584
rect 9426 49583 9498 49584
rect 9550 49583 9622 49584
rect 9674 49583 9746 49584
rect 9798 49583 10251 49584
rect 10303 49583 10375 49584
rect 10427 49583 10499 49584
rect 10551 49583 10623 49584
rect 10675 49583 10747 49584
rect 10799 49583 10871 49584
rect 10923 49583 10995 49584
rect 11047 49583 11119 49584
rect 11171 49583 11243 49584
rect 11295 49583 11367 49584
rect 11419 49583 11489 49584
rect 3489 49571 11489 49583
rect 11651 49392 11662 49950
rect 3316 49381 11662 49392
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49302 4863 49335
rect 4915 49302 4987 49335
rect 5039 49302 7277 49335
rect 7329 49302 7401 49335
rect 7453 49302 7525 49335
rect 7577 49302 7649 49335
rect 7701 49302 9939 49335
rect 9991 49302 10063 49335
rect 10115 49302 11816 49335
rect 3162 49230 11816 49302
rect 3162 49227 4863 49230
rect 4915 49227 4987 49230
rect 5039 49227 7277 49230
rect 7329 49227 7401 49230
rect 7453 49227 7525 49230
rect 7577 49227 7649 49230
rect 7701 49227 9939 49230
rect 9991 49227 10063 49230
rect 10115 49227 11816 49230
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49178 4863 49181
rect 4915 49178 4987 49181
rect 5039 49178 7277 49181
rect 7329 49178 7401 49181
rect 7453 49178 7525 49181
rect 7577 49178 7649 49181
rect 7701 49178 9939 49181
rect 9991 49178 10063 49181
rect 10115 49178 11816 49181
rect 3162 49106 11816 49178
rect 3162 49073 4863 49106
rect 4915 49073 4987 49106
rect 5039 49073 7277 49106
rect 7329 49073 7401 49106
rect 7453 49073 7525 49106
rect 7577 49073 7649 49106
rect 7701 49073 9939 49106
rect 9991 49073 10063 49106
rect 10115 49073 11816 49106
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49016 11662 49027
rect 3316 48458 3327 49016
rect 3489 48825 11489 48837
rect 3489 48824 3559 48825
rect 3611 48824 3683 48825
rect 3735 48824 3807 48825
rect 3859 48824 3931 48825
rect 3983 48824 4055 48825
rect 4107 48824 4179 48825
rect 4231 48824 4303 48825
rect 4355 48824 4427 48825
rect 4479 48824 4551 48825
rect 4603 48824 4675 48825
rect 4727 48824 5180 48825
rect 5232 48824 5304 48825
rect 5356 48824 5428 48825
rect 5480 48824 5552 48825
rect 5604 48824 5676 48825
rect 5728 48824 5800 48825
rect 5852 48824 5924 48825
rect 5976 48824 6048 48825
rect 6100 48824 6172 48825
rect 6224 48824 6296 48825
rect 6348 48824 6420 48825
rect 6472 48824 6544 48825
rect 6596 48824 6668 48825
rect 6720 48824 6792 48825
rect 6844 48824 6916 48825
rect 6968 48824 7040 48825
rect 7092 48824 7886 48825
rect 7938 48824 8010 48825
rect 8062 48824 8134 48825
rect 8186 48824 8258 48825
rect 8310 48824 8382 48825
rect 8434 48824 8506 48825
rect 8558 48824 8630 48825
rect 8682 48824 8754 48825
rect 8806 48824 8878 48825
rect 8930 48824 9002 48825
rect 9054 48824 9126 48825
rect 9178 48824 9250 48825
rect 9302 48824 9374 48825
rect 9426 48824 9498 48825
rect 9550 48824 9622 48825
rect 9674 48824 9746 48825
rect 9798 48824 10251 48825
rect 10303 48824 10375 48825
rect 10427 48824 10499 48825
rect 10551 48824 10623 48825
rect 10675 48824 10747 48825
rect 10799 48824 10871 48825
rect 10923 48824 10995 48825
rect 11047 48824 11119 48825
rect 11171 48824 11243 48825
rect 11295 48824 11367 48825
rect 11419 48824 11489 48825
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48773 3559 48778
rect 3611 48773 3683 48778
rect 3735 48773 3807 48778
rect 3859 48773 3931 48778
rect 3983 48773 4055 48778
rect 4107 48773 4179 48778
rect 4231 48773 4303 48778
rect 4355 48773 4427 48778
rect 4479 48773 4551 48778
rect 4603 48773 4675 48778
rect 4727 48773 5180 48778
rect 5232 48773 5304 48778
rect 5356 48773 5428 48778
rect 5480 48773 5552 48778
rect 5604 48773 5676 48778
rect 5728 48773 5800 48778
rect 5852 48773 5924 48778
rect 5976 48773 6048 48778
rect 6100 48773 6172 48778
rect 6224 48773 6296 48778
rect 6348 48773 6420 48778
rect 6472 48773 6544 48778
rect 6596 48773 6668 48778
rect 6720 48773 6792 48778
rect 6844 48773 6916 48778
rect 6968 48773 7040 48778
rect 7092 48773 7886 48778
rect 7938 48773 8010 48778
rect 8062 48773 8134 48778
rect 8186 48773 8258 48778
rect 8310 48773 8382 48778
rect 8434 48773 8506 48778
rect 8558 48773 8630 48778
rect 8682 48773 8754 48778
rect 8806 48773 8878 48778
rect 8930 48773 9002 48778
rect 9054 48773 9126 48778
rect 9178 48773 9250 48778
rect 9302 48773 9374 48778
rect 9426 48773 9498 48778
rect 9550 48773 9622 48778
rect 9674 48773 9746 48778
rect 9798 48773 10251 48778
rect 10303 48773 10375 48778
rect 10427 48773 10499 48778
rect 10551 48773 10623 48778
rect 10675 48773 10747 48778
rect 10799 48773 10871 48778
rect 10923 48773 10995 48778
rect 11047 48773 11119 48778
rect 11171 48773 11243 48778
rect 11295 48773 11367 48778
rect 11419 48773 11489 48778
rect 3489 48701 11489 48773
rect 3489 48696 3559 48701
rect 3611 48696 3683 48701
rect 3735 48696 3807 48701
rect 3859 48696 3931 48701
rect 3983 48696 4055 48701
rect 4107 48696 4179 48701
rect 4231 48696 4303 48701
rect 4355 48696 4427 48701
rect 4479 48696 4551 48701
rect 4603 48696 4675 48701
rect 4727 48696 5180 48701
rect 5232 48696 5304 48701
rect 5356 48696 5428 48701
rect 5480 48696 5552 48701
rect 5604 48696 5676 48701
rect 5728 48696 5800 48701
rect 5852 48696 5924 48701
rect 5976 48696 6048 48701
rect 6100 48696 6172 48701
rect 6224 48696 6296 48701
rect 6348 48696 6420 48701
rect 6472 48696 6544 48701
rect 6596 48696 6668 48701
rect 6720 48696 6792 48701
rect 6844 48696 6916 48701
rect 6968 48696 7040 48701
rect 7092 48696 7886 48701
rect 7938 48696 8010 48701
rect 8062 48696 8134 48701
rect 8186 48696 8258 48701
rect 8310 48696 8382 48701
rect 8434 48696 8506 48701
rect 8558 48696 8630 48701
rect 8682 48696 8754 48701
rect 8806 48696 8878 48701
rect 8930 48696 9002 48701
rect 9054 48696 9126 48701
rect 9178 48696 9250 48701
rect 9302 48696 9374 48701
rect 9426 48696 9498 48701
rect 9550 48696 9622 48701
rect 9674 48696 9746 48701
rect 9798 48696 10251 48701
rect 10303 48696 10375 48701
rect 10427 48696 10499 48701
rect 10551 48696 10623 48701
rect 10675 48696 10747 48701
rect 10799 48696 10871 48701
rect 10923 48696 10995 48701
rect 11047 48696 11119 48701
rect 11171 48696 11243 48701
rect 11295 48696 11367 48701
rect 11419 48696 11489 48701
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48649 3559 48650
rect 3611 48649 3683 48650
rect 3735 48649 3807 48650
rect 3859 48649 3931 48650
rect 3983 48649 4055 48650
rect 4107 48649 4179 48650
rect 4231 48649 4303 48650
rect 4355 48649 4427 48650
rect 4479 48649 4551 48650
rect 4603 48649 4675 48650
rect 4727 48649 5180 48650
rect 5232 48649 5304 48650
rect 5356 48649 5428 48650
rect 5480 48649 5552 48650
rect 5604 48649 5676 48650
rect 5728 48649 5800 48650
rect 5852 48649 5924 48650
rect 5976 48649 6048 48650
rect 6100 48649 6172 48650
rect 6224 48649 6296 48650
rect 6348 48649 6420 48650
rect 6472 48649 6544 48650
rect 6596 48649 6668 48650
rect 6720 48649 6792 48650
rect 6844 48649 6916 48650
rect 6968 48649 7040 48650
rect 7092 48649 7886 48650
rect 7938 48649 8010 48650
rect 8062 48649 8134 48650
rect 8186 48649 8258 48650
rect 8310 48649 8382 48650
rect 8434 48649 8506 48650
rect 8558 48649 8630 48650
rect 8682 48649 8754 48650
rect 8806 48649 8878 48650
rect 8930 48649 9002 48650
rect 9054 48649 9126 48650
rect 9178 48649 9250 48650
rect 9302 48649 9374 48650
rect 9426 48649 9498 48650
rect 9550 48649 9622 48650
rect 9674 48649 9746 48650
rect 9798 48649 10251 48650
rect 10303 48649 10375 48650
rect 10427 48649 10499 48650
rect 10551 48649 10623 48650
rect 10675 48649 10747 48650
rect 10799 48649 10871 48650
rect 10923 48649 10995 48650
rect 11047 48649 11119 48650
rect 11171 48649 11243 48650
rect 11295 48649 11367 48650
rect 11419 48649 11489 48650
rect 3489 48637 11489 48649
rect 11651 48458 11662 49016
rect 3316 48447 11662 48458
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48383 4863 48401
rect 4915 48383 4987 48401
rect 5039 48383 7277 48401
rect 7329 48383 7401 48401
rect 7453 48383 7525 48401
rect 7577 48383 7649 48401
rect 7701 48383 9939 48401
rect 9991 48383 10063 48401
rect 10115 48383 11816 48401
rect 3162 48376 11816 48383
rect 11862 48376 11873 51900
rect 3105 48311 11873 48376
rect 3105 48293 4863 48311
rect 4915 48293 4987 48311
rect 5039 48293 7277 48311
rect 7329 48293 7401 48311
rect 7453 48293 7525 48311
rect 7577 48293 7649 48311
rect 7701 48293 9939 48311
rect 9991 48293 10063 48311
rect 10115 48293 11873 48311
rect 3105 48247 3142 48293
rect 11836 48247 11873 48293
rect 3105 48236 11873 48247
rect 12059 48022 12070 52254
rect 2908 48011 12070 48022
rect 2908 47988 3016 48011
rect 11962 47988 12070 48011
rect 2908 47936 2934 47988
rect 2986 47936 3016 47988
rect 11962 47936 11992 47988
rect 12044 47936 12070 47988
rect 2908 47864 3016 47936
rect 11962 47864 12070 47936
rect 2908 47812 2934 47864
rect 2986 47812 3016 47864
rect 11962 47812 11992 47864
rect 12044 47812 12070 47864
rect 2908 47740 3016 47812
rect 11962 47740 12070 47812
rect 2908 47688 2934 47740
rect 2986 47688 3016 47740
rect 11962 47688 11992 47740
rect 12044 47688 12070 47740
rect 2908 47665 3016 47688
rect 11962 47665 12070 47688
rect 12416 47665 12427 52611
rect 2551 47654 12427 47665
rect 12753 52611 14907 52622
rect 12753 47665 12764 52611
rect 14710 52586 14907 52611
rect 14710 52574 14968 52586
rect 14710 52522 14904 52574
rect 14956 52522 14968 52574
rect 14710 52466 14968 52522
rect 14710 52414 14904 52466
rect 14956 52414 14968 52466
rect 14710 52358 14968 52414
rect 14710 52306 14904 52358
rect 14956 52306 14968 52358
rect 14710 52250 14968 52306
rect 14710 52198 14904 52250
rect 14956 52198 14968 52250
rect 14710 52142 14968 52198
rect 14710 52090 14904 52142
rect 14956 52090 14968 52142
rect 14710 52034 14968 52090
rect 14710 51982 14904 52034
rect 14956 51982 14968 52034
rect 14710 51926 14968 51982
rect 14710 51874 14904 51926
rect 14956 51874 14968 51926
rect 14710 51818 14968 51874
rect 14710 51766 14904 51818
rect 14956 51766 14968 51818
rect 14710 51710 14968 51766
rect 14710 51658 14904 51710
rect 14956 51658 14968 51710
rect 14710 51622 14968 51658
rect 14710 51422 14721 51622
rect 14892 51602 14968 51622
rect 14892 51550 14904 51602
rect 14956 51550 14968 51602
rect 14892 51494 14968 51550
rect 14892 51442 14904 51494
rect 14956 51442 14968 51494
rect 14892 51422 14968 51442
rect 14710 51386 14968 51422
rect 14710 51334 14904 51386
rect 14956 51334 14968 51386
rect 14710 51278 14968 51334
rect 14710 51226 14904 51278
rect 14956 51226 14968 51278
rect 14710 51214 14968 51226
rect 14710 50422 14907 51214
rect 14710 49854 14721 50422
rect 14710 48854 14907 49854
rect 14710 48654 14721 48854
rect 14710 47665 14907 48654
rect 12753 47654 14907 47665
rect 71 42647 725 42658
rect 71 41658 268 42647
rect 257 41458 268 41658
rect 71 40458 268 41458
rect 257 40258 268 40458
rect 71 39258 268 40258
rect 257 39058 268 39258
rect 71 38186 268 39058
rect 10 38174 268 38186
rect 10 38122 22 38174
rect 74 38122 268 38174
rect 10 38066 268 38122
rect 10 38014 22 38066
rect 74 38058 268 38066
rect 74 38014 86 38058
rect 10 37958 86 38014
rect 10 37906 22 37958
rect 74 37906 86 37958
rect 10 37858 86 37906
rect 257 37858 268 38058
rect 10 37850 268 37858
rect 10 37798 22 37850
rect 74 37798 268 37850
rect 10 37742 268 37798
rect 10 37690 22 37742
rect 74 37690 268 37742
rect 10 37634 268 37690
rect 10 37582 22 37634
rect 74 37582 268 37634
rect 10 37526 268 37582
rect 10 37474 22 37526
rect 74 37474 268 37526
rect 10 37418 268 37474
rect 10 37366 22 37418
rect 74 37366 268 37418
rect 10 37310 268 37366
rect 10 37258 22 37310
rect 74 37258 268 37310
rect 10 37202 268 37258
rect 10 37150 22 37202
rect 74 37150 268 37202
rect 10 37094 268 37150
rect 10 37042 22 37094
rect 74 37042 268 37094
rect 10 36986 268 37042
rect 10 36934 22 36986
rect 74 36934 268 36986
rect 10 36878 268 36934
rect 10 36826 22 36878
rect 74 36858 268 36878
rect 74 36826 86 36858
rect 10 36814 86 36826
rect 257 36658 268 36858
rect 71 35658 268 36658
rect 257 35458 268 35658
rect 71 34458 268 35458
rect 257 34258 268 34458
rect 71 33258 268 34258
rect 257 33058 268 33258
rect 71 32058 268 33058
rect 257 31858 268 32058
rect 71 30858 268 31858
rect 257 30658 268 30858
rect 71 29658 268 30658
rect 257 29458 268 29658
rect 71 28458 268 29458
rect 257 28258 268 28458
rect 71 27258 268 28258
rect 257 27058 268 27258
rect 71 26058 268 27058
rect 257 25858 268 26058
rect 71 24858 268 25858
rect 257 24658 268 24858
rect 71 23658 268 24658
rect 257 23458 268 23658
rect 71 22458 268 23458
rect 257 21390 268 22458
rect 71 20390 268 21390
rect 257 20190 268 20390
rect 71 19190 268 20190
rect 257 18990 268 19190
rect 71 17990 268 18990
rect 257 17790 268 17990
rect 71 16790 268 17790
rect 257 16590 268 16790
rect 71 15590 268 16590
rect 257 15390 268 15590
rect 71 14390 268 15390
rect 257 14190 268 14390
rect 71 13190 268 14190
rect 257 12990 268 13190
rect 71 11990 268 12990
rect 257 11790 268 11990
rect 71 10790 268 11790
rect 257 10590 268 10790
rect 71 9590 268 10590
rect 257 9390 268 9590
rect 71 8390 268 9390
rect 257 8190 268 8390
rect 71 7190 268 8190
rect 257 6990 268 7190
rect 71 5990 268 6990
rect 257 5790 268 5990
rect 71 4790 268 5790
rect 257 4590 268 4790
rect 71 3590 268 4590
rect 257 3390 268 3590
rect 71 2390 268 3390
rect 257 2190 268 2390
rect 71 1201 268 2190
rect 714 1201 725 42647
rect 13012 42647 14907 42658
rect 13012 27201 13023 42647
rect 13969 41658 14264 42647
rect 13969 41458 13980 41658
rect 14253 41458 14264 41658
rect 13969 40458 14264 41458
rect 13969 40258 13980 40458
rect 14253 40258 14264 40458
rect 13969 39258 14264 40258
rect 13969 39058 13980 39258
rect 14253 39058 14264 39258
rect 13969 38058 14264 39058
rect 13969 37858 13980 38058
rect 14253 37858 14264 38058
rect 13969 36858 14264 37858
rect 13969 36658 13980 36858
rect 14253 36658 14264 36858
rect 13969 35658 14264 36658
rect 13969 35458 13980 35658
rect 14253 35458 14264 35658
rect 13969 34458 14264 35458
rect 13969 34258 13980 34458
rect 14253 34258 14264 34458
rect 13969 33258 14264 34258
rect 13969 33058 13980 33258
rect 14253 33058 14264 33258
rect 13969 32058 14264 33058
rect 13969 31858 13980 32058
rect 14253 31858 14264 32058
rect 13969 30858 14264 31858
rect 13969 30658 13980 30858
rect 14253 30658 14264 30858
rect 13969 29658 14264 30658
rect 13969 29458 13980 29658
rect 14253 29458 14264 29658
rect 13969 28458 14264 29458
rect 13969 28190 13980 28458
rect 14253 28190 14264 28458
rect 13969 27201 14264 28190
rect 13012 27190 14264 27201
rect 71 1190 725 1201
rect 14253 1201 14264 27190
rect 14710 41658 14907 42647
rect 14710 41458 14721 41658
rect 14710 40458 14907 41458
rect 14710 40258 14721 40458
rect 14710 39258 14907 40258
rect 14710 39058 14721 39258
rect 14710 38186 14907 39058
rect 14710 38174 14968 38186
rect 14710 38122 14904 38174
rect 14956 38122 14968 38174
rect 14710 38066 14968 38122
rect 14710 38058 14904 38066
rect 14710 37858 14721 38058
rect 14892 38014 14904 38058
rect 14956 38014 14968 38066
rect 14892 37958 14968 38014
rect 14892 37906 14904 37958
rect 14956 37906 14968 37958
rect 14892 37858 14968 37906
rect 14710 37850 14968 37858
rect 14710 37798 14904 37850
rect 14956 37798 14968 37850
rect 14710 37742 14968 37798
rect 14710 37690 14904 37742
rect 14956 37690 14968 37742
rect 14710 37634 14968 37690
rect 14710 37582 14904 37634
rect 14956 37582 14968 37634
rect 14710 37526 14968 37582
rect 14710 37474 14904 37526
rect 14956 37474 14968 37526
rect 14710 37418 14968 37474
rect 14710 37366 14904 37418
rect 14956 37366 14968 37418
rect 14710 37310 14968 37366
rect 14710 37258 14904 37310
rect 14956 37258 14968 37310
rect 14710 37202 14968 37258
rect 14710 37150 14904 37202
rect 14956 37150 14968 37202
rect 14710 37094 14968 37150
rect 14710 37042 14904 37094
rect 14956 37042 14968 37094
rect 14710 36986 14968 37042
rect 14710 36934 14904 36986
rect 14956 36934 14968 36986
rect 14710 36878 14968 36934
rect 14710 36858 14904 36878
rect 14710 36658 14721 36858
rect 14892 36826 14904 36858
rect 14956 36826 14968 36878
rect 14892 36814 14968 36826
rect 14710 35658 14907 36658
rect 14710 35458 14721 35658
rect 14710 34458 14907 35458
rect 14710 34258 14721 34458
rect 14710 33258 14907 34258
rect 14710 33058 14721 33258
rect 14710 32058 14907 33058
rect 14710 31858 14721 32058
rect 14710 30858 14907 31858
rect 14710 30658 14721 30858
rect 14710 29658 14907 30658
rect 14710 29458 14721 29658
rect 14710 28458 14907 29458
rect 14710 28258 14721 28458
rect 14710 27258 14907 28258
rect 14710 27058 14721 27258
rect 14710 26058 14907 27058
rect 14710 25858 14721 26058
rect 14710 24858 14907 25858
rect 14710 24658 14721 24858
rect 14710 23658 14907 24658
rect 14710 23458 14721 23658
rect 14710 22458 14907 23458
rect 14710 21390 14721 22458
rect 14710 20390 14907 21390
rect 14710 20190 14721 20390
rect 14710 19190 14907 20190
rect 14710 18990 14721 19190
rect 14710 17990 14907 18990
rect 14710 17790 14721 17990
rect 14710 16790 14907 17790
rect 14710 16590 14721 16790
rect 14710 15590 14907 16590
rect 14710 15390 14721 15590
rect 14710 14390 14907 15390
rect 14710 14190 14721 14390
rect 14710 13190 14907 14190
rect 14710 12990 14721 13190
rect 14710 11990 14907 12990
rect 14710 11790 14721 11990
rect 14710 10790 14907 11790
rect 14710 10590 14721 10790
rect 14710 9590 14907 10590
rect 14710 9390 14721 9590
rect 14710 8390 14907 9390
rect 14710 8190 14721 8390
rect 14710 7190 14907 8190
rect 14710 6990 14721 7190
rect 14710 5990 14907 6990
rect 14710 5790 14721 5990
rect 14710 4790 14907 5790
rect 14710 4590 14721 4790
rect 14710 3590 14907 4590
rect 14710 3390 14721 3590
rect 14710 2390 14907 3390
rect 14710 2190 14721 2390
rect 14710 1201 14907 2190
rect 14253 1190 14907 1201
<< via1 >>
rect 2501 57105 2553 57108
rect 2609 57105 2661 57108
rect 4871 57105 4923 57108
rect 4979 57105 5031 57108
rect 7247 57105 7299 57108
rect 7355 57105 7407 57108
rect 7463 57105 7515 57108
rect 7571 57105 7623 57108
rect 7679 57105 7731 57108
rect 9947 57105 9999 57108
rect 10055 57105 10107 57108
rect 12317 57105 12369 57108
rect 12425 57105 12477 57108
rect 2501 57059 2553 57105
rect 2609 57059 2661 57105
rect 4871 57059 4923 57105
rect 4979 57059 5031 57105
rect 7247 57059 7299 57105
rect 7355 57059 7407 57105
rect 7463 57059 7515 57105
rect 7571 57059 7623 57105
rect 7679 57059 7731 57105
rect 9947 57059 9999 57105
rect 10055 57059 10107 57105
rect 12317 57059 12369 57105
rect 12425 57059 12477 57105
rect 2501 57056 2553 57059
rect 2609 57056 2661 57059
rect 4871 57056 4923 57059
rect 4979 57056 5031 57059
rect 7247 57056 7299 57059
rect 7355 57056 7407 57059
rect 7463 57056 7515 57059
rect 7571 57056 7623 57059
rect 7679 57056 7731 57059
rect 9947 57056 9999 57059
rect 10055 57056 10107 57059
rect 12317 57056 12369 57059
rect 12425 57056 12477 57059
rect 917 56617 969 56669
rect 1041 56617 1093 56669
rect 1165 56617 1217 56669
rect 1289 56617 1341 56669
rect 1413 56617 1465 56669
rect 1537 56617 1589 56669
rect 1661 56617 1713 56669
rect 1785 56617 1837 56669
rect 917 56493 969 56545
rect 1041 56493 1093 56545
rect 1165 56493 1217 56545
rect 1289 56493 1341 56545
rect 1413 56493 1465 56545
rect 1537 56493 1589 56545
rect 1661 56493 1713 56545
rect 1785 56493 1837 56545
rect 917 56369 969 56421
rect 1041 56369 1093 56421
rect 1165 56369 1217 56421
rect 1289 56369 1341 56421
rect 1413 56369 1465 56421
rect 1537 56369 1589 56421
rect 1661 56369 1713 56421
rect 1785 56369 1837 56421
rect 917 56245 969 56297
rect 1041 56245 1093 56297
rect 1165 56245 1217 56297
rect 1289 56245 1341 56297
rect 1413 56245 1465 56297
rect 1537 56245 1589 56297
rect 1661 56245 1713 56297
rect 1785 56245 1837 56297
rect 917 56121 969 56173
rect 1041 56121 1093 56173
rect 1165 56121 1217 56173
rect 1289 56121 1341 56173
rect 1413 56121 1465 56173
rect 1537 56121 1589 56173
rect 1661 56121 1713 56173
rect 1785 56121 1837 56173
rect 917 55997 969 56049
rect 1041 55997 1093 56049
rect 1165 55997 1217 56049
rect 1289 55997 1341 56049
rect 1413 55997 1465 56049
rect 1537 55997 1589 56049
rect 1661 55997 1713 56049
rect 1785 55997 1837 56049
rect 917 55873 969 55925
rect 1041 55873 1093 55925
rect 1165 55873 1217 55925
rect 1289 55873 1341 55925
rect 1413 55873 1465 55925
rect 1537 55873 1589 55925
rect 1661 55873 1713 55925
rect 1785 55873 1837 55925
rect 917 55749 969 55801
rect 1041 55749 1093 55801
rect 1165 55749 1217 55801
rect 1289 55749 1341 55801
rect 1413 55749 1465 55801
rect 1537 55749 1589 55801
rect 1661 55749 1713 55801
rect 1785 55749 1837 55801
rect 917 55625 969 55677
rect 1041 55625 1093 55677
rect 1165 55625 1217 55677
rect 1289 55625 1341 55677
rect 1413 55625 1465 55677
rect 1537 55625 1589 55677
rect 1661 55625 1713 55677
rect 1785 55625 1837 55677
rect 917 55501 969 55553
rect 1041 55501 1093 55553
rect 1165 55501 1217 55553
rect 1289 55501 1341 55553
rect 1413 55501 1465 55553
rect 1537 55501 1589 55553
rect 1661 55501 1713 55553
rect 1785 55501 1837 55553
rect 917 55377 969 55429
rect 1041 55377 1093 55429
rect 1165 55377 1217 55429
rect 1289 55377 1341 55429
rect 1413 55377 1465 55429
rect 1537 55377 1589 55429
rect 1661 55377 1713 55429
rect 1785 55377 1837 55429
rect 917 55253 969 55305
rect 1041 55253 1093 55305
rect 1165 55253 1217 55305
rect 1289 55253 1341 55305
rect 1413 55253 1465 55305
rect 1537 55253 1589 55305
rect 1661 55253 1713 55305
rect 1785 55253 1837 55305
rect 917 55129 969 55181
rect 1041 55129 1093 55181
rect 1165 55129 1217 55181
rect 1289 55129 1341 55181
rect 1413 55129 1465 55181
rect 1537 55129 1589 55181
rect 1661 55129 1713 55181
rect 1785 55129 1837 55181
rect 917 55005 969 55057
rect 1041 55005 1093 55057
rect 1165 55005 1217 55057
rect 1289 55005 1341 55057
rect 1413 55005 1465 55057
rect 1537 55005 1589 55057
rect 1661 55005 1713 55057
rect 1785 55005 1837 55057
rect 917 54881 969 54933
rect 1041 54881 1093 54933
rect 1165 54881 1217 54933
rect 1289 54881 1341 54933
rect 1413 54881 1465 54933
rect 1537 54881 1589 54933
rect 1661 54881 1713 54933
rect 1785 54881 1837 54933
rect 917 54757 969 54809
rect 1041 54757 1093 54809
rect 1165 54757 1217 54809
rect 1289 54757 1341 54809
rect 1413 54757 1465 54809
rect 1537 54757 1589 54809
rect 1661 54757 1713 54809
rect 1785 54757 1837 54809
rect 917 54633 969 54685
rect 1041 54633 1093 54685
rect 1165 54633 1217 54685
rect 1289 54633 1341 54685
rect 1413 54633 1465 54685
rect 1537 54633 1589 54685
rect 1661 54633 1713 54685
rect 1785 54633 1837 54685
rect 917 54509 969 54561
rect 1041 54509 1093 54561
rect 1165 54509 1217 54561
rect 1289 54509 1341 54561
rect 1413 54509 1465 54561
rect 1537 54509 1589 54561
rect 1661 54509 1713 54561
rect 1785 54509 1837 54561
rect 917 54385 969 54437
rect 1041 54385 1093 54437
rect 1165 54385 1217 54437
rect 1289 54385 1341 54437
rect 1413 54385 1465 54437
rect 1537 54385 1589 54437
rect 1661 54385 1713 54437
rect 1785 54385 1837 54437
rect 917 54261 969 54313
rect 1041 54261 1093 54313
rect 1165 54261 1217 54313
rect 1289 54261 1341 54313
rect 1413 54261 1465 54313
rect 1537 54261 1589 54313
rect 1661 54261 1713 54313
rect 1785 54261 1837 54313
rect 917 54137 969 54189
rect 1041 54137 1093 54189
rect 1165 54137 1217 54189
rect 1289 54137 1341 54189
rect 1413 54137 1465 54189
rect 1537 54137 1589 54189
rect 1661 54137 1713 54189
rect 1785 54137 1837 54189
rect 917 54013 969 54065
rect 1041 54013 1093 54065
rect 1165 54013 1217 54065
rect 1289 54013 1341 54065
rect 1413 54013 1465 54065
rect 1537 54013 1589 54065
rect 1661 54013 1713 54065
rect 1785 54013 1837 54065
rect 917 53889 969 53941
rect 1041 53889 1093 53941
rect 1165 53889 1217 53941
rect 1289 53889 1341 53941
rect 1413 53889 1465 53941
rect 1537 53889 1589 53941
rect 1661 53889 1713 53941
rect 1785 53889 1837 53941
rect 917 53765 969 53817
rect 1041 53765 1093 53817
rect 1165 53765 1217 53817
rect 1289 53765 1341 53817
rect 1413 53765 1465 53817
rect 1537 53765 1589 53817
rect 1661 53765 1713 53817
rect 1785 53765 1837 53817
rect 917 53641 969 53693
rect 1041 53641 1093 53693
rect 1165 53641 1217 53693
rect 1289 53641 1341 53693
rect 1413 53641 1465 53693
rect 1537 53641 1589 53693
rect 1661 53641 1713 53693
rect 1785 53641 1837 53693
rect 2833 56617 2885 56669
rect 2957 56617 3009 56669
rect 3081 56617 3133 56669
rect 3205 56617 3257 56669
rect 3329 56617 3381 56669
rect 3453 56617 3505 56669
rect 3577 56617 3629 56669
rect 3701 56617 3753 56669
rect 2833 56493 2885 56545
rect 2957 56493 3009 56545
rect 3081 56493 3133 56545
rect 3205 56493 3257 56545
rect 3329 56493 3381 56545
rect 3453 56493 3505 56545
rect 3577 56493 3629 56545
rect 3701 56493 3753 56545
rect 2833 56369 2885 56421
rect 2957 56369 3009 56421
rect 3081 56369 3133 56421
rect 3205 56369 3257 56421
rect 3329 56369 3381 56421
rect 3453 56369 3505 56421
rect 3577 56369 3629 56421
rect 3701 56369 3753 56421
rect 2833 56245 2885 56297
rect 2957 56245 3009 56297
rect 3081 56245 3133 56297
rect 3205 56245 3257 56297
rect 3329 56245 3381 56297
rect 3453 56245 3505 56297
rect 3577 56245 3629 56297
rect 3701 56245 3753 56297
rect 2833 56121 2885 56173
rect 2957 56121 3009 56173
rect 3081 56121 3133 56173
rect 3205 56121 3257 56173
rect 3329 56121 3381 56173
rect 3453 56121 3505 56173
rect 3577 56121 3629 56173
rect 3701 56121 3753 56173
rect 2833 55997 2885 56049
rect 2957 55997 3009 56049
rect 3081 55997 3133 56049
rect 3205 55997 3257 56049
rect 3329 55997 3381 56049
rect 3453 55997 3505 56049
rect 3577 55997 3629 56049
rect 3701 55997 3753 56049
rect 2833 55873 2885 55925
rect 2957 55873 3009 55925
rect 3081 55873 3133 55925
rect 3205 55873 3257 55925
rect 3329 55873 3381 55925
rect 3453 55873 3505 55925
rect 3577 55873 3629 55925
rect 3701 55873 3753 55925
rect 2833 55749 2885 55801
rect 2957 55749 3009 55801
rect 3081 55749 3133 55801
rect 3205 55749 3257 55801
rect 3329 55749 3381 55801
rect 3453 55749 3505 55801
rect 3577 55749 3629 55801
rect 3701 55749 3753 55801
rect 2833 55625 2885 55677
rect 2957 55625 3009 55677
rect 3081 55625 3133 55677
rect 3205 55625 3257 55677
rect 3329 55625 3381 55677
rect 3453 55625 3505 55677
rect 3577 55625 3629 55677
rect 3701 55625 3753 55677
rect 2833 55501 2885 55553
rect 2957 55501 3009 55553
rect 3081 55501 3133 55553
rect 3205 55501 3257 55553
rect 3329 55501 3381 55553
rect 3453 55501 3505 55553
rect 3577 55501 3629 55553
rect 3701 55501 3753 55553
rect 2833 55377 2885 55429
rect 2957 55377 3009 55429
rect 3081 55377 3133 55429
rect 3205 55377 3257 55429
rect 3329 55377 3381 55429
rect 3453 55377 3505 55429
rect 3577 55377 3629 55429
rect 3701 55377 3753 55429
rect 2833 55253 2885 55305
rect 2957 55253 3009 55305
rect 3081 55253 3133 55305
rect 3205 55253 3257 55305
rect 3329 55253 3381 55305
rect 3453 55253 3505 55305
rect 3577 55253 3629 55305
rect 3701 55253 3753 55305
rect 2833 55129 2885 55181
rect 2957 55129 3009 55181
rect 3081 55129 3133 55181
rect 3205 55129 3257 55181
rect 3329 55129 3381 55181
rect 3453 55129 3505 55181
rect 3577 55129 3629 55181
rect 3701 55129 3753 55181
rect 2833 55005 2885 55057
rect 2957 55005 3009 55057
rect 3081 55005 3133 55057
rect 3205 55005 3257 55057
rect 3329 55005 3381 55057
rect 3453 55005 3505 55057
rect 3577 55005 3629 55057
rect 3701 55005 3753 55057
rect 2833 54881 2885 54933
rect 2957 54881 3009 54933
rect 3081 54881 3133 54933
rect 3205 54881 3257 54933
rect 3329 54881 3381 54933
rect 3453 54881 3505 54933
rect 3577 54881 3629 54933
rect 3701 54881 3753 54933
rect 2833 54757 2885 54809
rect 2957 54757 3009 54809
rect 3081 54757 3133 54809
rect 3205 54757 3257 54809
rect 3329 54757 3381 54809
rect 3453 54757 3505 54809
rect 3577 54757 3629 54809
rect 3701 54757 3753 54809
rect 2833 54633 2885 54685
rect 2957 54633 3009 54685
rect 3081 54633 3133 54685
rect 3205 54633 3257 54685
rect 3329 54633 3381 54685
rect 3453 54633 3505 54685
rect 3577 54633 3629 54685
rect 3701 54633 3753 54685
rect 2833 54509 2885 54561
rect 2957 54509 3009 54561
rect 3081 54509 3133 54561
rect 3205 54509 3257 54561
rect 3329 54509 3381 54561
rect 3453 54509 3505 54561
rect 3577 54509 3629 54561
rect 3701 54509 3753 54561
rect 2833 54385 2885 54437
rect 2957 54385 3009 54437
rect 3081 54385 3133 54437
rect 3205 54385 3257 54437
rect 3329 54385 3381 54437
rect 3453 54385 3505 54437
rect 3577 54385 3629 54437
rect 3701 54385 3753 54437
rect 2833 54261 2885 54313
rect 2957 54261 3009 54313
rect 3081 54261 3133 54313
rect 3205 54261 3257 54313
rect 3329 54261 3381 54313
rect 3453 54261 3505 54313
rect 3577 54261 3629 54313
rect 3701 54261 3753 54313
rect 2833 54137 2885 54189
rect 2957 54137 3009 54189
rect 3081 54137 3133 54189
rect 3205 54137 3257 54189
rect 3329 54137 3381 54189
rect 3453 54137 3505 54189
rect 3577 54137 3629 54189
rect 3701 54137 3753 54189
rect 2833 54013 2885 54065
rect 2957 54013 3009 54065
rect 3081 54013 3133 54065
rect 3205 54013 3257 54065
rect 3329 54013 3381 54065
rect 3453 54013 3505 54065
rect 3577 54013 3629 54065
rect 3701 54013 3753 54065
rect 2833 53889 2885 53941
rect 2957 53889 3009 53941
rect 3081 53889 3133 53941
rect 3205 53889 3257 53941
rect 3329 53889 3381 53941
rect 3453 53889 3505 53941
rect 3577 53889 3629 53941
rect 3701 53889 3753 53941
rect 2833 53765 2885 53817
rect 2957 53765 3009 53817
rect 3081 53765 3133 53817
rect 3205 53765 3257 53817
rect 3329 53765 3381 53817
rect 3453 53765 3505 53817
rect 3577 53765 3629 53817
rect 3701 53765 3753 53817
rect 2833 53641 2885 53693
rect 2957 53641 3009 53693
rect 3081 53641 3133 53693
rect 3205 53641 3257 53693
rect 3329 53641 3381 53693
rect 3453 53641 3505 53693
rect 3577 53641 3629 53693
rect 3701 53641 3753 53693
rect 4340 56617 4392 56669
rect 4464 56617 4516 56669
rect 4588 56617 4640 56669
rect 4712 56617 4764 56669
rect 4340 56493 4392 56545
rect 4464 56493 4516 56545
rect 4588 56493 4640 56545
rect 4712 56493 4764 56545
rect 4340 56369 4392 56421
rect 4464 56369 4516 56421
rect 4588 56369 4640 56421
rect 4712 56369 4764 56421
rect 4340 56245 4392 56297
rect 4464 56245 4516 56297
rect 4588 56245 4640 56297
rect 4712 56245 4764 56297
rect 4340 56121 4392 56173
rect 4464 56121 4516 56173
rect 4588 56121 4640 56173
rect 4712 56121 4764 56173
rect 4340 55997 4392 56049
rect 4464 55997 4516 56049
rect 4588 55997 4640 56049
rect 4712 55997 4764 56049
rect 4340 55873 4392 55925
rect 4464 55873 4516 55925
rect 4588 55873 4640 55925
rect 4712 55873 4764 55925
rect 4340 55749 4392 55801
rect 4464 55749 4516 55801
rect 4588 55749 4640 55801
rect 4712 55749 4764 55801
rect 4340 55625 4392 55677
rect 4464 55625 4516 55677
rect 4588 55625 4640 55677
rect 4712 55625 4764 55677
rect 4340 55501 4392 55553
rect 4464 55501 4516 55553
rect 4588 55501 4640 55553
rect 4712 55501 4764 55553
rect 4340 55377 4392 55429
rect 4464 55377 4516 55429
rect 4588 55377 4640 55429
rect 4712 55377 4764 55429
rect 4340 55253 4392 55305
rect 4464 55253 4516 55305
rect 4588 55253 4640 55305
rect 4712 55253 4764 55305
rect 4340 55129 4392 55181
rect 4464 55129 4516 55181
rect 4588 55129 4640 55181
rect 4712 55129 4764 55181
rect 4340 55005 4392 55057
rect 4464 55005 4516 55057
rect 4588 55005 4640 55057
rect 4712 55005 4764 55057
rect 4340 54881 4392 54933
rect 4464 54881 4516 54933
rect 4588 54881 4640 54933
rect 4712 54881 4764 54933
rect 4340 54757 4392 54809
rect 4464 54757 4516 54809
rect 4588 54757 4640 54809
rect 4712 54757 4764 54809
rect 4340 54633 4392 54685
rect 4464 54633 4516 54685
rect 4588 54633 4640 54685
rect 4712 54633 4764 54685
rect 4340 54509 4392 54561
rect 4464 54509 4516 54561
rect 4588 54509 4640 54561
rect 4712 54509 4764 54561
rect 4340 54385 4392 54437
rect 4464 54385 4516 54437
rect 4588 54385 4640 54437
rect 4712 54385 4764 54437
rect 4340 54261 4392 54313
rect 4464 54261 4516 54313
rect 4588 54261 4640 54313
rect 4712 54261 4764 54313
rect 4340 54137 4392 54189
rect 4464 54137 4516 54189
rect 4588 54137 4640 54189
rect 4712 54137 4764 54189
rect 4340 54013 4392 54065
rect 4464 54013 4516 54065
rect 4588 54013 4640 54065
rect 4712 54013 4764 54065
rect 4340 53889 4392 53941
rect 4464 53889 4516 53941
rect 4588 53889 4640 53941
rect 4712 53889 4764 53941
rect 4340 53765 4392 53817
rect 4464 53765 4516 53817
rect 4588 53765 4640 53817
rect 4712 53765 4764 53817
rect 4340 53641 4392 53693
rect 4464 53641 4516 53693
rect 4588 53641 4640 53693
rect 4712 53641 4764 53693
rect 6297 56617 6349 56669
rect 6421 56617 6473 56669
rect 6545 56617 6597 56669
rect 6669 56617 6721 56669
rect 6793 56617 6845 56669
rect 6917 56617 6969 56669
rect 7041 56617 7093 56669
rect 6297 56493 6349 56545
rect 6421 56493 6473 56545
rect 6545 56493 6597 56545
rect 6669 56493 6721 56545
rect 6793 56493 6845 56545
rect 6917 56493 6969 56545
rect 7041 56493 7093 56545
rect 6297 56369 6349 56421
rect 6421 56369 6473 56421
rect 6545 56369 6597 56421
rect 6669 56369 6721 56421
rect 6793 56369 6845 56421
rect 6917 56369 6969 56421
rect 7041 56369 7093 56421
rect 6297 56245 6349 56297
rect 6421 56245 6473 56297
rect 6545 56245 6597 56297
rect 6669 56245 6721 56297
rect 6793 56245 6845 56297
rect 6917 56245 6969 56297
rect 7041 56245 7093 56297
rect 6297 56121 6349 56173
rect 6421 56121 6473 56173
rect 6545 56121 6597 56173
rect 6669 56121 6721 56173
rect 6793 56121 6845 56173
rect 6917 56121 6969 56173
rect 7041 56121 7093 56173
rect 6297 55997 6349 56049
rect 6421 55997 6473 56049
rect 6545 55997 6597 56049
rect 6669 55997 6721 56049
rect 6793 55997 6845 56049
rect 6917 55997 6969 56049
rect 7041 55997 7093 56049
rect 6297 55873 6349 55925
rect 6421 55873 6473 55925
rect 6545 55873 6597 55925
rect 6669 55873 6721 55925
rect 6793 55873 6845 55925
rect 6917 55873 6969 55925
rect 7041 55873 7093 55925
rect 6297 55749 6349 55801
rect 6421 55749 6473 55801
rect 6545 55749 6597 55801
rect 6669 55749 6721 55801
rect 6793 55749 6845 55801
rect 6917 55749 6969 55801
rect 7041 55749 7093 55801
rect 6297 55625 6349 55677
rect 6421 55625 6473 55677
rect 6545 55625 6597 55677
rect 6669 55625 6721 55677
rect 6793 55625 6845 55677
rect 6917 55625 6969 55677
rect 7041 55625 7093 55677
rect 6297 55501 6349 55553
rect 6421 55501 6473 55553
rect 6545 55501 6597 55553
rect 6669 55501 6721 55553
rect 6793 55501 6845 55553
rect 6917 55501 6969 55553
rect 7041 55501 7093 55553
rect 6297 55377 6349 55429
rect 6421 55377 6473 55429
rect 6545 55377 6597 55429
rect 6669 55377 6721 55429
rect 6793 55377 6845 55429
rect 6917 55377 6969 55429
rect 7041 55377 7093 55429
rect 6297 55253 6349 55305
rect 6421 55253 6473 55305
rect 6545 55253 6597 55305
rect 6669 55253 6721 55305
rect 6793 55253 6845 55305
rect 6917 55253 6969 55305
rect 7041 55253 7093 55305
rect 6297 55129 6349 55181
rect 6421 55129 6473 55181
rect 6545 55129 6597 55181
rect 6669 55129 6721 55181
rect 6793 55129 6845 55181
rect 6917 55129 6969 55181
rect 7041 55129 7093 55181
rect 6297 55005 6349 55057
rect 6421 55005 6473 55057
rect 6545 55005 6597 55057
rect 6669 55005 6721 55057
rect 6793 55005 6845 55057
rect 6917 55005 6969 55057
rect 7041 55005 7093 55057
rect 6297 54881 6349 54933
rect 6421 54881 6473 54933
rect 6545 54881 6597 54933
rect 6669 54881 6721 54933
rect 6793 54881 6845 54933
rect 6917 54881 6969 54933
rect 7041 54881 7093 54933
rect 6297 54757 6349 54809
rect 6421 54757 6473 54809
rect 6545 54757 6597 54809
rect 6669 54757 6721 54809
rect 6793 54757 6845 54809
rect 6917 54757 6969 54809
rect 7041 54757 7093 54809
rect 6297 54633 6349 54685
rect 6421 54633 6473 54685
rect 6545 54633 6597 54685
rect 6669 54633 6721 54685
rect 6793 54633 6845 54685
rect 6917 54633 6969 54685
rect 7041 54633 7093 54685
rect 6297 54509 6349 54561
rect 6421 54509 6473 54561
rect 6545 54509 6597 54561
rect 6669 54509 6721 54561
rect 6793 54509 6845 54561
rect 6917 54509 6969 54561
rect 7041 54509 7093 54561
rect 6297 54385 6349 54437
rect 6421 54385 6473 54437
rect 6545 54385 6597 54437
rect 6669 54385 6721 54437
rect 6793 54385 6845 54437
rect 6917 54385 6969 54437
rect 7041 54385 7093 54437
rect 6297 54261 6349 54313
rect 6421 54261 6473 54313
rect 6545 54261 6597 54313
rect 6669 54261 6721 54313
rect 6793 54261 6845 54313
rect 6917 54261 6969 54313
rect 7041 54261 7093 54313
rect 6297 54137 6349 54189
rect 6421 54137 6473 54189
rect 6545 54137 6597 54189
rect 6669 54137 6721 54189
rect 6793 54137 6845 54189
rect 6917 54137 6969 54189
rect 7041 54137 7093 54189
rect 6297 54013 6349 54065
rect 6421 54013 6473 54065
rect 6545 54013 6597 54065
rect 6669 54013 6721 54065
rect 6793 54013 6845 54065
rect 6917 54013 6969 54065
rect 7041 54013 7093 54065
rect 6297 53889 6349 53941
rect 6421 53889 6473 53941
rect 6545 53889 6597 53941
rect 6669 53889 6721 53941
rect 6793 53889 6845 53941
rect 6917 53889 6969 53941
rect 7041 53889 7093 53941
rect 6297 53765 6349 53817
rect 6421 53765 6473 53817
rect 6545 53765 6597 53817
rect 6669 53765 6721 53817
rect 6793 53765 6845 53817
rect 6917 53765 6969 53817
rect 7041 53765 7093 53817
rect 6297 53641 6349 53693
rect 6421 53641 6473 53693
rect 6545 53641 6597 53693
rect 6669 53641 6721 53693
rect 6793 53641 6845 53693
rect 6917 53641 6969 53693
rect 7041 53641 7093 53693
rect 7885 56617 7937 56669
rect 8009 56617 8061 56669
rect 8133 56617 8185 56669
rect 8257 56617 8309 56669
rect 8381 56617 8433 56669
rect 8505 56617 8557 56669
rect 8629 56617 8681 56669
rect 7885 56493 7937 56545
rect 8009 56493 8061 56545
rect 8133 56493 8185 56545
rect 8257 56493 8309 56545
rect 8381 56493 8433 56545
rect 8505 56493 8557 56545
rect 8629 56493 8681 56545
rect 7885 56369 7937 56421
rect 8009 56369 8061 56421
rect 8133 56369 8185 56421
rect 8257 56369 8309 56421
rect 8381 56369 8433 56421
rect 8505 56369 8557 56421
rect 8629 56369 8681 56421
rect 7885 56245 7937 56297
rect 8009 56245 8061 56297
rect 8133 56245 8185 56297
rect 8257 56245 8309 56297
rect 8381 56245 8433 56297
rect 8505 56245 8557 56297
rect 8629 56245 8681 56297
rect 7885 56121 7937 56173
rect 8009 56121 8061 56173
rect 8133 56121 8185 56173
rect 8257 56121 8309 56173
rect 8381 56121 8433 56173
rect 8505 56121 8557 56173
rect 8629 56121 8681 56173
rect 7885 55997 7937 56049
rect 8009 55997 8061 56049
rect 8133 55997 8185 56049
rect 8257 55997 8309 56049
rect 8381 55997 8433 56049
rect 8505 55997 8557 56049
rect 8629 55997 8681 56049
rect 7885 55873 7937 55925
rect 8009 55873 8061 55925
rect 8133 55873 8185 55925
rect 8257 55873 8309 55925
rect 8381 55873 8433 55925
rect 8505 55873 8557 55925
rect 8629 55873 8681 55925
rect 7885 55749 7937 55801
rect 8009 55749 8061 55801
rect 8133 55749 8185 55801
rect 8257 55749 8309 55801
rect 8381 55749 8433 55801
rect 8505 55749 8557 55801
rect 8629 55749 8681 55801
rect 7885 55625 7937 55677
rect 8009 55625 8061 55677
rect 8133 55625 8185 55677
rect 8257 55625 8309 55677
rect 8381 55625 8433 55677
rect 8505 55625 8557 55677
rect 8629 55625 8681 55677
rect 7885 55501 7937 55553
rect 8009 55501 8061 55553
rect 8133 55501 8185 55553
rect 8257 55501 8309 55553
rect 8381 55501 8433 55553
rect 8505 55501 8557 55553
rect 8629 55501 8681 55553
rect 7885 55377 7937 55429
rect 8009 55377 8061 55429
rect 8133 55377 8185 55429
rect 8257 55377 8309 55429
rect 8381 55377 8433 55429
rect 8505 55377 8557 55429
rect 8629 55377 8681 55429
rect 7885 55253 7937 55305
rect 8009 55253 8061 55305
rect 8133 55253 8185 55305
rect 8257 55253 8309 55305
rect 8381 55253 8433 55305
rect 8505 55253 8557 55305
rect 8629 55253 8681 55305
rect 7885 55129 7937 55181
rect 8009 55129 8061 55181
rect 8133 55129 8185 55181
rect 8257 55129 8309 55181
rect 8381 55129 8433 55181
rect 8505 55129 8557 55181
rect 8629 55129 8681 55181
rect 7885 55005 7937 55057
rect 8009 55005 8061 55057
rect 8133 55005 8185 55057
rect 8257 55005 8309 55057
rect 8381 55005 8433 55057
rect 8505 55005 8557 55057
rect 8629 55005 8681 55057
rect 7885 54881 7937 54933
rect 8009 54881 8061 54933
rect 8133 54881 8185 54933
rect 8257 54881 8309 54933
rect 8381 54881 8433 54933
rect 8505 54881 8557 54933
rect 8629 54881 8681 54933
rect 7885 54757 7937 54809
rect 8009 54757 8061 54809
rect 8133 54757 8185 54809
rect 8257 54757 8309 54809
rect 8381 54757 8433 54809
rect 8505 54757 8557 54809
rect 8629 54757 8681 54809
rect 7885 54633 7937 54685
rect 8009 54633 8061 54685
rect 8133 54633 8185 54685
rect 8257 54633 8309 54685
rect 8381 54633 8433 54685
rect 8505 54633 8557 54685
rect 8629 54633 8681 54685
rect 7885 54509 7937 54561
rect 8009 54509 8061 54561
rect 8133 54509 8185 54561
rect 8257 54509 8309 54561
rect 8381 54509 8433 54561
rect 8505 54509 8557 54561
rect 8629 54509 8681 54561
rect 7885 54385 7937 54437
rect 8009 54385 8061 54437
rect 8133 54385 8185 54437
rect 8257 54385 8309 54437
rect 8381 54385 8433 54437
rect 8505 54385 8557 54437
rect 8629 54385 8681 54437
rect 7885 54261 7937 54313
rect 8009 54261 8061 54313
rect 8133 54261 8185 54313
rect 8257 54261 8309 54313
rect 8381 54261 8433 54313
rect 8505 54261 8557 54313
rect 8629 54261 8681 54313
rect 7885 54137 7937 54189
rect 8009 54137 8061 54189
rect 8133 54137 8185 54189
rect 8257 54137 8309 54189
rect 8381 54137 8433 54189
rect 8505 54137 8557 54189
rect 8629 54137 8681 54189
rect 7885 54013 7937 54065
rect 8009 54013 8061 54065
rect 8133 54013 8185 54065
rect 8257 54013 8309 54065
rect 8381 54013 8433 54065
rect 8505 54013 8557 54065
rect 8629 54013 8681 54065
rect 7885 53889 7937 53941
rect 8009 53889 8061 53941
rect 8133 53889 8185 53941
rect 8257 53889 8309 53941
rect 8381 53889 8433 53941
rect 8505 53889 8557 53941
rect 8629 53889 8681 53941
rect 7885 53765 7937 53817
rect 8009 53765 8061 53817
rect 8133 53765 8185 53817
rect 8257 53765 8309 53817
rect 8381 53765 8433 53817
rect 8505 53765 8557 53817
rect 8629 53765 8681 53817
rect 7885 53641 7937 53693
rect 8009 53641 8061 53693
rect 8133 53641 8185 53693
rect 8257 53641 8309 53693
rect 8381 53641 8433 53693
rect 8505 53641 8557 53693
rect 8629 53641 8681 53693
rect 10214 56617 10266 56669
rect 10338 56617 10390 56669
rect 10462 56617 10514 56669
rect 10586 56617 10638 56669
rect 10214 56493 10266 56545
rect 10338 56493 10390 56545
rect 10462 56493 10514 56545
rect 10586 56493 10638 56545
rect 10214 56369 10266 56421
rect 10338 56369 10390 56421
rect 10462 56369 10514 56421
rect 10586 56369 10638 56421
rect 10214 56245 10266 56297
rect 10338 56245 10390 56297
rect 10462 56245 10514 56297
rect 10586 56245 10638 56297
rect 10214 56121 10266 56173
rect 10338 56121 10390 56173
rect 10462 56121 10514 56173
rect 10586 56121 10638 56173
rect 10214 55997 10266 56049
rect 10338 55997 10390 56049
rect 10462 55997 10514 56049
rect 10586 55997 10638 56049
rect 10214 55873 10266 55925
rect 10338 55873 10390 55925
rect 10462 55873 10514 55925
rect 10586 55873 10638 55925
rect 10214 55749 10266 55801
rect 10338 55749 10390 55801
rect 10462 55749 10514 55801
rect 10586 55749 10638 55801
rect 10214 55625 10266 55677
rect 10338 55625 10390 55677
rect 10462 55625 10514 55677
rect 10586 55625 10638 55677
rect 10214 55501 10266 55553
rect 10338 55501 10390 55553
rect 10462 55501 10514 55553
rect 10586 55501 10638 55553
rect 10214 55377 10266 55429
rect 10338 55377 10390 55429
rect 10462 55377 10514 55429
rect 10586 55377 10638 55429
rect 10214 55253 10266 55305
rect 10338 55253 10390 55305
rect 10462 55253 10514 55305
rect 10586 55253 10638 55305
rect 10214 55129 10266 55181
rect 10338 55129 10390 55181
rect 10462 55129 10514 55181
rect 10586 55129 10638 55181
rect 10214 55005 10266 55057
rect 10338 55005 10390 55057
rect 10462 55005 10514 55057
rect 10586 55005 10638 55057
rect 10214 54881 10266 54933
rect 10338 54881 10390 54933
rect 10462 54881 10514 54933
rect 10586 54881 10638 54933
rect 10214 54757 10266 54809
rect 10338 54757 10390 54809
rect 10462 54757 10514 54809
rect 10586 54757 10638 54809
rect 10214 54633 10266 54685
rect 10338 54633 10390 54685
rect 10462 54633 10514 54685
rect 10586 54633 10638 54685
rect 10214 54509 10266 54561
rect 10338 54509 10390 54561
rect 10462 54509 10514 54561
rect 10586 54509 10638 54561
rect 10214 54385 10266 54437
rect 10338 54385 10390 54437
rect 10462 54385 10514 54437
rect 10586 54385 10638 54437
rect 10214 54261 10266 54313
rect 10338 54261 10390 54313
rect 10462 54261 10514 54313
rect 10586 54261 10638 54313
rect 10214 54137 10266 54189
rect 10338 54137 10390 54189
rect 10462 54137 10514 54189
rect 10586 54137 10638 54189
rect 10214 54013 10266 54065
rect 10338 54013 10390 54065
rect 10462 54013 10514 54065
rect 10586 54013 10638 54065
rect 10214 53889 10266 53941
rect 10338 53889 10390 53941
rect 10462 53889 10514 53941
rect 10586 53889 10638 53941
rect 10214 53765 10266 53817
rect 10338 53765 10390 53817
rect 10462 53765 10514 53817
rect 10586 53765 10638 53817
rect 10214 53641 10266 53693
rect 10338 53641 10390 53693
rect 10462 53641 10514 53693
rect 10586 53641 10638 53693
rect 11225 56617 11277 56669
rect 11349 56617 11401 56669
rect 11473 56617 11525 56669
rect 11597 56617 11649 56669
rect 11721 56617 11773 56669
rect 11845 56617 11897 56669
rect 11969 56617 12021 56669
rect 12093 56617 12145 56669
rect 11225 56493 11277 56545
rect 11349 56493 11401 56545
rect 11473 56493 11525 56545
rect 11597 56493 11649 56545
rect 11721 56493 11773 56545
rect 11845 56493 11897 56545
rect 11969 56493 12021 56545
rect 12093 56493 12145 56545
rect 11225 56369 11277 56421
rect 11349 56369 11401 56421
rect 11473 56369 11525 56421
rect 11597 56369 11649 56421
rect 11721 56369 11773 56421
rect 11845 56369 11897 56421
rect 11969 56369 12021 56421
rect 12093 56369 12145 56421
rect 11225 56245 11277 56297
rect 11349 56245 11401 56297
rect 11473 56245 11525 56297
rect 11597 56245 11649 56297
rect 11721 56245 11773 56297
rect 11845 56245 11897 56297
rect 11969 56245 12021 56297
rect 12093 56245 12145 56297
rect 11225 56121 11277 56173
rect 11349 56121 11401 56173
rect 11473 56121 11525 56173
rect 11597 56121 11649 56173
rect 11721 56121 11773 56173
rect 11845 56121 11897 56173
rect 11969 56121 12021 56173
rect 12093 56121 12145 56173
rect 11225 55997 11277 56049
rect 11349 55997 11401 56049
rect 11473 55997 11525 56049
rect 11597 55997 11649 56049
rect 11721 55997 11773 56049
rect 11845 55997 11897 56049
rect 11969 55997 12021 56049
rect 12093 55997 12145 56049
rect 11225 55873 11277 55925
rect 11349 55873 11401 55925
rect 11473 55873 11525 55925
rect 11597 55873 11649 55925
rect 11721 55873 11773 55925
rect 11845 55873 11897 55925
rect 11969 55873 12021 55925
rect 12093 55873 12145 55925
rect 11225 55749 11277 55801
rect 11349 55749 11401 55801
rect 11473 55749 11525 55801
rect 11597 55749 11649 55801
rect 11721 55749 11773 55801
rect 11845 55749 11897 55801
rect 11969 55749 12021 55801
rect 12093 55749 12145 55801
rect 11225 55625 11277 55677
rect 11349 55625 11401 55677
rect 11473 55625 11525 55677
rect 11597 55625 11649 55677
rect 11721 55625 11773 55677
rect 11845 55625 11897 55677
rect 11969 55625 12021 55677
rect 12093 55625 12145 55677
rect 11225 55501 11277 55553
rect 11349 55501 11401 55553
rect 11473 55501 11525 55553
rect 11597 55501 11649 55553
rect 11721 55501 11773 55553
rect 11845 55501 11897 55553
rect 11969 55501 12021 55553
rect 12093 55501 12145 55553
rect 11225 55377 11277 55429
rect 11349 55377 11401 55429
rect 11473 55377 11525 55429
rect 11597 55377 11649 55429
rect 11721 55377 11773 55429
rect 11845 55377 11897 55429
rect 11969 55377 12021 55429
rect 12093 55377 12145 55429
rect 11225 55253 11277 55305
rect 11349 55253 11401 55305
rect 11473 55253 11525 55305
rect 11597 55253 11649 55305
rect 11721 55253 11773 55305
rect 11845 55253 11897 55305
rect 11969 55253 12021 55305
rect 12093 55253 12145 55305
rect 11225 55129 11277 55181
rect 11349 55129 11401 55181
rect 11473 55129 11525 55181
rect 11597 55129 11649 55181
rect 11721 55129 11773 55181
rect 11845 55129 11897 55181
rect 11969 55129 12021 55181
rect 12093 55129 12145 55181
rect 11225 55005 11277 55057
rect 11349 55005 11401 55057
rect 11473 55005 11525 55057
rect 11597 55005 11649 55057
rect 11721 55005 11773 55057
rect 11845 55005 11897 55057
rect 11969 55005 12021 55057
rect 12093 55005 12145 55057
rect 11225 54881 11277 54933
rect 11349 54881 11401 54933
rect 11473 54881 11525 54933
rect 11597 54881 11649 54933
rect 11721 54881 11773 54933
rect 11845 54881 11897 54933
rect 11969 54881 12021 54933
rect 12093 54881 12145 54933
rect 11225 54757 11277 54809
rect 11349 54757 11401 54809
rect 11473 54757 11525 54809
rect 11597 54757 11649 54809
rect 11721 54757 11773 54809
rect 11845 54757 11897 54809
rect 11969 54757 12021 54809
rect 12093 54757 12145 54809
rect 11225 54633 11277 54685
rect 11349 54633 11401 54685
rect 11473 54633 11525 54685
rect 11597 54633 11649 54685
rect 11721 54633 11773 54685
rect 11845 54633 11897 54685
rect 11969 54633 12021 54685
rect 12093 54633 12145 54685
rect 11225 54509 11277 54561
rect 11349 54509 11401 54561
rect 11473 54509 11525 54561
rect 11597 54509 11649 54561
rect 11721 54509 11773 54561
rect 11845 54509 11897 54561
rect 11969 54509 12021 54561
rect 12093 54509 12145 54561
rect 11225 54385 11277 54437
rect 11349 54385 11401 54437
rect 11473 54385 11525 54437
rect 11597 54385 11649 54437
rect 11721 54385 11773 54437
rect 11845 54385 11897 54437
rect 11969 54385 12021 54437
rect 12093 54385 12145 54437
rect 11225 54261 11277 54313
rect 11349 54261 11401 54313
rect 11473 54261 11525 54313
rect 11597 54261 11649 54313
rect 11721 54261 11773 54313
rect 11845 54261 11897 54313
rect 11969 54261 12021 54313
rect 12093 54261 12145 54313
rect 11225 54137 11277 54189
rect 11349 54137 11401 54189
rect 11473 54137 11525 54189
rect 11597 54137 11649 54189
rect 11721 54137 11773 54189
rect 11845 54137 11897 54189
rect 11969 54137 12021 54189
rect 12093 54137 12145 54189
rect 11225 54013 11277 54065
rect 11349 54013 11401 54065
rect 11473 54013 11525 54065
rect 11597 54013 11649 54065
rect 11721 54013 11773 54065
rect 11845 54013 11897 54065
rect 11969 54013 12021 54065
rect 12093 54013 12145 54065
rect 11225 53889 11277 53941
rect 11349 53889 11401 53941
rect 11473 53889 11525 53941
rect 11597 53889 11649 53941
rect 11721 53889 11773 53941
rect 11845 53889 11897 53941
rect 11969 53889 12021 53941
rect 12093 53889 12145 53941
rect 11225 53765 11277 53817
rect 11349 53765 11401 53817
rect 11473 53765 11525 53817
rect 11597 53765 11649 53817
rect 11721 53765 11773 53817
rect 11845 53765 11897 53817
rect 11969 53765 12021 53817
rect 12093 53765 12145 53817
rect 11225 53641 11277 53693
rect 11349 53641 11401 53693
rect 11473 53641 11525 53693
rect 11597 53641 11649 53693
rect 11721 53641 11773 53693
rect 11845 53641 11897 53693
rect 11969 53641 12021 53693
rect 12093 53641 12145 53693
rect 13141 56617 13193 56669
rect 13265 56617 13317 56669
rect 13389 56617 13441 56669
rect 13513 56617 13565 56669
rect 13637 56617 13689 56669
rect 13761 56617 13813 56669
rect 13885 56617 13937 56669
rect 14009 56617 14061 56669
rect 13141 56493 13193 56545
rect 13265 56493 13317 56545
rect 13389 56493 13441 56545
rect 13513 56493 13565 56545
rect 13637 56493 13689 56545
rect 13761 56493 13813 56545
rect 13885 56493 13937 56545
rect 14009 56493 14061 56545
rect 13141 56369 13193 56421
rect 13265 56369 13317 56421
rect 13389 56369 13441 56421
rect 13513 56369 13565 56421
rect 13637 56369 13689 56421
rect 13761 56369 13813 56421
rect 13885 56369 13937 56421
rect 14009 56369 14061 56421
rect 13141 56245 13193 56297
rect 13265 56245 13317 56297
rect 13389 56245 13441 56297
rect 13513 56245 13565 56297
rect 13637 56245 13689 56297
rect 13761 56245 13813 56297
rect 13885 56245 13937 56297
rect 14009 56245 14061 56297
rect 13141 56121 13193 56173
rect 13265 56121 13317 56173
rect 13389 56121 13441 56173
rect 13513 56121 13565 56173
rect 13637 56121 13689 56173
rect 13761 56121 13813 56173
rect 13885 56121 13937 56173
rect 14009 56121 14061 56173
rect 13141 55997 13193 56049
rect 13265 55997 13317 56049
rect 13389 55997 13441 56049
rect 13513 55997 13565 56049
rect 13637 55997 13689 56049
rect 13761 55997 13813 56049
rect 13885 55997 13937 56049
rect 14009 55997 14061 56049
rect 13141 55873 13193 55925
rect 13265 55873 13317 55925
rect 13389 55873 13441 55925
rect 13513 55873 13565 55925
rect 13637 55873 13689 55925
rect 13761 55873 13813 55925
rect 13885 55873 13937 55925
rect 14009 55873 14061 55925
rect 13141 55749 13193 55801
rect 13265 55749 13317 55801
rect 13389 55749 13441 55801
rect 13513 55749 13565 55801
rect 13637 55749 13689 55801
rect 13761 55749 13813 55801
rect 13885 55749 13937 55801
rect 14009 55749 14061 55801
rect 13141 55625 13193 55677
rect 13265 55625 13317 55677
rect 13389 55625 13441 55677
rect 13513 55625 13565 55677
rect 13637 55625 13689 55677
rect 13761 55625 13813 55677
rect 13885 55625 13937 55677
rect 14009 55625 14061 55677
rect 13141 55501 13193 55553
rect 13265 55501 13317 55553
rect 13389 55501 13441 55553
rect 13513 55501 13565 55553
rect 13637 55501 13689 55553
rect 13761 55501 13813 55553
rect 13885 55501 13937 55553
rect 14009 55501 14061 55553
rect 13141 55377 13193 55429
rect 13265 55377 13317 55429
rect 13389 55377 13441 55429
rect 13513 55377 13565 55429
rect 13637 55377 13689 55429
rect 13761 55377 13813 55429
rect 13885 55377 13937 55429
rect 14009 55377 14061 55429
rect 13141 55253 13193 55305
rect 13265 55253 13317 55305
rect 13389 55253 13441 55305
rect 13513 55253 13565 55305
rect 13637 55253 13689 55305
rect 13761 55253 13813 55305
rect 13885 55253 13937 55305
rect 14009 55253 14061 55305
rect 13141 55129 13193 55181
rect 13265 55129 13317 55181
rect 13389 55129 13441 55181
rect 13513 55129 13565 55181
rect 13637 55129 13689 55181
rect 13761 55129 13813 55181
rect 13885 55129 13937 55181
rect 14009 55129 14061 55181
rect 13141 55005 13193 55057
rect 13265 55005 13317 55057
rect 13389 55005 13441 55057
rect 13513 55005 13565 55057
rect 13637 55005 13689 55057
rect 13761 55005 13813 55057
rect 13885 55005 13937 55057
rect 14009 55005 14061 55057
rect 13141 54881 13193 54933
rect 13265 54881 13317 54933
rect 13389 54881 13441 54933
rect 13513 54881 13565 54933
rect 13637 54881 13689 54933
rect 13761 54881 13813 54933
rect 13885 54881 13937 54933
rect 14009 54881 14061 54933
rect 13141 54757 13193 54809
rect 13265 54757 13317 54809
rect 13389 54757 13441 54809
rect 13513 54757 13565 54809
rect 13637 54757 13689 54809
rect 13761 54757 13813 54809
rect 13885 54757 13937 54809
rect 14009 54757 14061 54809
rect 13141 54633 13193 54685
rect 13265 54633 13317 54685
rect 13389 54633 13441 54685
rect 13513 54633 13565 54685
rect 13637 54633 13689 54685
rect 13761 54633 13813 54685
rect 13885 54633 13937 54685
rect 14009 54633 14061 54685
rect 13141 54509 13193 54561
rect 13265 54509 13317 54561
rect 13389 54509 13441 54561
rect 13513 54509 13565 54561
rect 13637 54509 13689 54561
rect 13761 54509 13813 54561
rect 13885 54509 13937 54561
rect 14009 54509 14061 54561
rect 13141 54385 13193 54437
rect 13265 54385 13317 54437
rect 13389 54385 13441 54437
rect 13513 54385 13565 54437
rect 13637 54385 13689 54437
rect 13761 54385 13813 54437
rect 13885 54385 13937 54437
rect 14009 54385 14061 54437
rect 13141 54261 13193 54313
rect 13265 54261 13317 54313
rect 13389 54261 13441 54313
rect 13513 54261 13565 54313
rect 13637 54261 13689 54313
rect 13761 54261 13813 54313
rect 13885 54261 13937 54313
rect 14009 54261 14061 54313
rect 13141 54137 13193 54189
rect 13265 54137 13317 54189
rect 13389 54137 13441 54189
rect 13513 54137 13565 54189
rect 13637 54137 13689 54189
rect 13761 54137 13813 54189
rect 13885 54137 13937 54189
rect 14009 54137 14061 54189
rect 13141 54013 13193 54065
rect 13265 54013 13317 54065
rect 13389 54013 13441 54065
rect 13513 54013 13565 54065
rect 13637 54013 13689 54065
rect 13761 54013 13813 54065
rect 13885 54013 13937 54065
rect 14009 54013 14061 54065
rect 13141 53889 13193 53941
rect 13265 53889 13317 53941
rect 13389 53889 13441 53941
rect 13513 53889 13565 53941
rect 13637 53889 13689 53941
rect 13761 53889 13813 53941
rect 13885 53889 13937 53941
rect 14009 53889 14061 53941
rect 13141 53765 13193 53817
rect 13265 53765 13317 53817
rect 13389 53765 13441 53817
rect 13513 53765 13565 53817
rect 13637 53765 13689 53817
rect 13761 53765 13813 53817
rect 13885 53765 13937 53817
rect 14009 53765 14061 53817
rect 13141 53641 13193 53693
rect 13265 53641 13317 53693
rect 13389 53641 13441 53693
rect 13513 53641 13565 53693
rect 13637 53641 13689 53693
rect 13761 53641 13813 53693
rect 13885 53641 13937 53693
rect 14009 53641 14061 53693
rect 2501 53432 2553 53484
rect 2609 53432 2661 53484
rect 4871 53432 4923 53484
rect 4979 53432 5031 53484
rect 7247 53432 7299 53484
rect 7355 53432 7407 53484
rect 7463 53432 7515 53484
rect 7571 53432 7623 53484
rect 7679 53432 7731 53484
rect 9947 53432 9999 53484
rect 10055 53432 10107 53484
rect 12317 53432 12369 53484
rect 12425 53432 12477 53484
rect 2501 53324 2553 53376
rect 2609 53324 2661 53376
rect 4871 53324 4923 53376
rect 4979 53324 5031 53376
rect 7247 53324 7299 53376
rect 7355 53324 7407 53376
rect 7463 53324 7515 53376
rect 7571 53324 7623 53376
rect 7679 53324 7731 53376
rect 9947 53324 9999 53376
rect 10055 53324 10107 53376
rect 12317 53324 12369 53376
rect 12425 53324 12477 53376
rect 2501 53251 2553 53268
rect 2609 53251 2661 53268
rect 4871 53251 4923 53268
rect 4979 53251 5031 53268
rect 7247 53251 7299 53268
rect 7355 53251 7407 53268
rect 7463 53251 7515 53268
rect 7571 53251 7623 53268
rect 7679 53251 7731 53268
rect 9947 53251 9999 53268
rect 10055 53251 10107 53268
rect 12317 53251 12369 53268
rect 12425 53251 12477 53268
rect 2501 53216 2553 53251
rect 2609 53216 2661 53251
rect 4871 53216 4923 53251
rect 4979 53216 5031 53251
rect 7247 53216 7299 53251
rect 7355 53216 7407 53251
rect 7463 53216 7515 53251
rect 7571 53216 7623 53251
rect 7679 53216 7731 53251
rect 9947 53216 9999 53251
rect 10055 53216 10107 53251
rect 12317 53216 12369 53251
rect 12425 53216 12477 53251
rect 22 52522 74 52574
rect 22 52414 74 52466
rect 22 52306 74 52358
rect 22 52198 74 52250
rect 22 52090 74 52142
rect 22 51982 74 52034
rect 22 51874 74 51926
rect 22 51766 74 51818
rect 22 51658 74 51710
rect 22 51550 74 51602
rect 22 51442 74 51494
rect 22 51334 74 51386
rect 22 51226 74 51278
rect 2810 52536 2862 52588
rect 2934 52536 2986 52588
rect 3058 52536 3110 52588
rect 3182 52536 3234 52588
rect 3306 52536 3358 52588
rect 3430 52536 3482 52588
rect 3554 52536 3606 52588
rect 3678 52536 3730 52588
rect 3802 52536 3854 52588
rect 3926 52536 3978 52588
rect 4050 52536 4102 52588
rect 4174 52536 4226 52588
rect 4298 52536 4350 52588
rect 4422 52536 4474 52588
rect 4546 52536 4598 52588
rect 4670 52536 4722 52588
rect 5180 52536 5232 52588
rect 5304 52536 5356 52588
rect 5428 52536 5480 52588
rect 5552 52536 5604 52588
rect 5676 52536 5728 52588
rect 5800 52536 5852 52588
rect 5924 52536 5976 52588
rect 6048 52536 6100 52588
rect 6172 52536 6224 52588
rect 6296 52536 6348 52588
rect 6420 52536 6472 52588
rect 6544 52536 6596 52588
rect 6668 52536 6720 52588
rect 6792 52536 6844 52588
rect 6916 52536 6968 52588
rect 7040 52536 7092 52588
rect 7886 52536 7938 52588
rect 8010 52536 8062 52588
rect 8134 52536 8186 52588
rect 8258 52536 8310 52588
rect 8382 52536 8434 52588
rect 8506 52536 8558 52588
rect 8630 52536 8682 52588
rect 8754 52536 8806 52588
rect 8878 52536 8930 52588
rect 9002 52536 9054 52588
rect 9126 52536 9178 52588
rect 9250 52536 9302 52588
rect 9374 52536 9426 52588
rect 9498 52536 9550 52588
rect 9622 52536 9674 52588
rect 9746 52536 9798 52588
rect 10256 52536 10308 52588
rect 10380 52536 10432 52588
rect 10504 52536 10556 52588
rect 10628 52536 10680 52588
rect 10752 52536 10804 52588
rect 10876 52536 10928 52588
rect 11000 52536 11052 52588
rect 11124 52536 11176 52588
rect 11248 52536 11300 52588
rect 11372 52536 11424 52588
rect 11496 52536 11548 52588
rect 11620 52536 11672 52588
rect 11744 52536 11796 52588
rect 11868 52536 11920 52588
rect 11992 52536 12044 52588
rect 12116 52536 12168 52588
rect 2810 52412 2862 52464
rect 2934 52412 2986 52464
rect 3058 52412 3110 52464
rect 3182 52412 3234 52464
rect 3306 52412 3358 52464
rect 3430 52412 3482 52464
rect 3554 52412 3606 52464
rect 3678 52412 3730 52464
rect 3802 52412 3854 52464
rect 3926 52412 3978 52464
rect 4050 52412 4102 52464
rect 4174 52412 4226 52464
rect 4298 52412 4350 52464
rect 4422 52412 4474 52464
rect 4546 52412 4598 52464
rect 4670 52412 4722 52464
rect 5180 52412 5232 52464
rect 5304 52412 5356 52464
rect 5428 52412 5480 52464
rect 5552 52412 5604 52464
rect 5676 52412 5728 52464
rect 5800 52412 5852 52464
rect 5924 52412 5976 52464
rect 6048 52412 6100 52464
rect 6172 52412 6224 52464
rect 6296 52412 6348 52464
rect 6420 52412 6472 52464
rect 6544 52412 6596 52464
rect 6668 52412 6720 52464
rect 6792 52412 6844 52464
rect 6916 52412 6968 52464
rect 7040 52412 7092 52464
rect 7886 52412 7938 52464
rect 8010 52412 8062 52464
rect 8134 52412 8186 52464
rect 8258 52412 8310 52464
rect 8382 52412 8434 52464
rect 8506 52412 8558 52464
rect 8630 52412 8682 52464
rect 8754 52412 8806 52464
rect 8878 52412 8930 52464
rect 9002 52412 9054 52464
rect 9126 52412 9178 52464
rect 9250 52412 9302 52464
rect 9374 52412 9426 52464
rect 9498 52412 9550 52464
rect 9622 52412 9674 52464
rect 9746 52412 9798 52464
rect 10256 52412 10308 52464
rect 10380 52412 10432 52464
rect 10504 52412 10556 52464
rect 10628 52412 10680 52464
rect 10752 52412 10804 52464
rect 10876 52412 10928 52464
rect 11000 52412 11052 52464
rect 11124 52412 11176 52464
rect 11248 52412 11300 52464
rect 11372 52412 11424 52464
rect 11496 52412 11548 52464
rect 11620 52412 11672 52464
rect 11744 52412 11796 52464
rect 11868 52412 11920 52464
rect 11992 52412 12044 52464
rect 12116 52412 12168 52464
rect 2810 52288 2862 52340
rect 2934 52288 2986 52340
rect 3058 52288 3110 52340
rect 3182 52288 3234 52340
rect 3306 52288 3358 52340
rect 3430 52288 3482 52340
rect 3554 52288 3606 52340
rect 3678 52288 3730 52340
rect 3802 52288 3854 52340
rect 3926 52288 3978 52340
rect 4050 52288 4102 52340
rect 4174 52288 4226 52340
rect 4298 52288 4350 52340
rect 4422 52288 4474 52340
rect 4546 52288 4598 52340
rect 4670 52288 4722 52340
rect 5180 52288 5232 52340
rect 5304 52288 5356 52340
rect 5428 52288 5480 52340
rect 5552 52288 5604 52340
rect 5676 52288 5728 52340
rect 5800 52288 5852 52340
rect 5924 52288 5976 52340
rect 6048 52288 6100 52340
rect 6172 52288 6224 52340
rect 6296 52288 6348 52340
rect 6420 52288 6472 52340
rect 6544 52288 6596 52340
rect 6668 52288 6720 52340
rect 6792 52288 6844 52340
rect 6916 52288 6968 52340
rect 7040 52288 7092 52340
rect 7886 52288 7938 52340
rect 8010 52288 8062 52340
rect 8134 52288 8186 52340
rect 8258 52288 8310 52340
rect 8382 52288 8434 52340
rect 8506 52288 8558 52340
rect 8630 52288 8682 52340
rect 8754 52288 8806 52340
rect 8878 52288 8930 52340
rect 9002 52288 9054 52340
rect 9126 52288 9178 52340
rect 9250 52288 9302 52340
rect 9374 52288 9426 52340
rect 9498 52288 9550 52340
rect 9622 52288 9674 52340
rect 9746 52288 9798 52340
rect 10256 52288 10308 52340
rect 10380 52288 10432 52340
rect 10504 52288 10556 52340
rect 10628 52288 10680 52340
rect 10752 52288 10804 52340
rect 10876 52288 10928 52340
rect 11000 52288 11052 52340
rect 11124 52288 11176 52340
rect 11248 52288 11300 52340
rect 11372 52288 11424 52340
rect 11496 52288 11548 52340
rect 11620 52288 11672 52340
rect 11744 52288 11796 52340
rect 11868 52288 11920 52340
rect 11992 52288 12044 52340
rect 12116 52288 12168 52340
rect 4863 51983 4915 52017
rect 4987 51983 5039 52017
rect 7277 51983 7329 52017
rect 7401 51983 7453 52017
rect 7525 51983 7577 52017
rect 7649 51983 7701 52017
rect 9939 51983 9991 52017
rect 10063 51983 10115 52017
rect 4863 51965 4915 51983
rect 4987 51965 5039 51983
rect 7277 51965 7329 51983
rect 7401 51965 7453 51983
rect 7525 51965 7577 51983
rect 7649 51965 7701 51983
rect 9939 51965 9991 51983
rect 10063 51965 10115 51983
rect 4863 51875 4915 51893
rect 4987 51875 5039 51893
rect 7277 51875 7329 51893
rect 7401 51875 7453 51893
rect 7525 51875 7577 51893
rect 7649 51875 7701 51893
rect 9939 51875 9991 51893
rect 10063 51875 10115 51893
rect 4863 51841 4915 51875
rect 4987 51841 5039 51875
rect 7277 51841 7329 51875
rect 7401 51841 7453 51875
rect 7525 51841 7577 51875
rect 7649 51841 7701 51875
rect 9939 51841 9991 51875
rect 10063 51841 10115 51875
rect 3559 51626 3611 51627
rect 3683 51626 3735 51627
rect 3807 51626 3859 51627
rect 3931 51626 3983 51627
rect 4055 51626 4107 51627
rect 4179 51626 4231 51627
rect 4303 51626 4355 51627
rect 4427 51626 4479 51627
rect 4551 51626 4603 51627
rect 4675 51626 4727 51627
rect 5180 51626 5232 51627
rect 5304 51626 5356 51627
rect 5428 51626 5480 51627
rect 5552 51626 5604 51627
rect 5676 51626 5728 51627
rect 5800 51626 5852 51627
rect 5924 51626 5976 51627
rect 6048 51626 6100 51627
rect 6172 51626 6224 51627
rect 6296 51626 6348 51627
rect 6420 51626 6472 51627
rect 6544 51626 6596 51627
rect 6668 51626 6720 51627
rect 6792 51626 6844 51627
rect 6916 51626 6968 51627
rect 7040 51626 7092 51627
rect 7886 51626 7938 51627
rect 8010 51626 8062 51627
rect 8134 51626 8186 51627
rect 8258 51626 8310 51627
rect 8382 51626 8434 51627
rect 8506 51626 8558 51627
rect 8630 51626 8682 51627
rect 8754 51626 8806 51627
rect 8878 51626 8930 51627
rect 9002 51626 9054 51627
rect 9126 51626 9178 51627
rect 9250 51626 9302 51627
rect 9374 51626 9426 51627
rect 9498 51626 9550 51627
rect 9622 51626 9674 51627
rect 9746 51626 9798 51627
rect 10251 51626 10303 51627
rect 10375 51626 10427 51627
rect 10499 51626 10551 51627
rect 10623 51626 10675 51627
rect 10747 51626 10799 51627
rect 10871 51626 10923 51627
rect 10995 51626 11047 51627
rect 11119 51626 11171 51627
rect 11243 51626 11295 51627
rect 11367 51626 11419 51627
rect 3559 51580 3611 51626
rect 3683 51580 3735 51626
rect 3807 51580 3859 51626
rect 3931 51580 3983 51626
rect 4055 51580 4107 51626
rect 4179 51580 4231 51626
rect 4303 51580 4355 51626
rect 4427 51580 4479 51626
rect 4551 51580 4603 51626
rect 4675 51580 4727 51626
rect 5180 51580 5232 51626
rect 5304 51580 5356 51626
rect 5428 51580 5480 51626
rect 5552 51580 5604 51626
rect 5676 51580 5728 51626
rect 5800 51580 5852 51626
rect 5924 51580 5976 51626
rect 6048 51580 6100 51626
rect 6172 51580 6224 51626
rect 6296 51580 6348 51626
rect 6420 51580 6472 51626
rect 6544 51580 6596 51626
rect 6668 51580 6720 51626
rect 6792 51580 6844 51626
rect 6916 51580 6968 51626
rect 7040 51580 7092 51626
rect 7886 51580 7938 51626
rect 8010 51580 8062 51626
rect 8134 51580 8186 51626
rect 8258 51580 8310 51626
rect 8382 51580 8434 51626
rect 8506 51580 8558 51626
rect 8630 51580 8682 51626
rect 8754 51580 8806 51626
rect 8878 51580 8930 51626
rect 9002 51580 9054 51626
rect 9126 51580 9178 51626
rect 9250 51580 9302 51626
rect 9374 51580 9426 51626
rect 9498 51580 9550 51626
rect 9622 51580 9674 51626
rect 9746 51580 9798 51626
rect 10251 51580 10303 51626
rect 10375 51580 10427 51626
rect 10499 51580 10551 51626
rect 10623 51580 10675 51626
rect 10747 51580 10799 51626
rect 10871 51580 10923 51626
rect 10995 51580 11047 51626
rect 11119 51580 11171 51626
rect 11243 51580 11295 51626
rect 11367 51580 11419 51626
rect 3559 51575 3611 51580
rect 3683 51575 3735 51580
rect 3807 51575 3859 51580
rect 3931 51575 3983 51580
rect 4055 51575 4107 51580
rect 4179 51575 4231 51580
rect 4303 51575 4355 51580
rect 4427 51575 4479 51580
rect 4551 51575 4603 51580
rect 4675 51575 4727 51580
rect 5180 51575 5232 51580
rect 5304 51575 5356 51580
rect 5428 51575 5480 51580
rect 5552 51575 5604 51580
rect 5676 51575 5728 51580
rect 5800 51575 5852 51580
rect 5924 51575 5976 51580
rect 6048 51575 6100 51580
rect 6172 51575 6224 51580
rect 6296 51575 6348 51580
rect 6420 51575 6472 51580
rect 6544 51575 6596 51580
rect 6668 51575 6720 51580
rect 6792 51575 6844 51580
rect 6916 51575 6968 51580
rect 7040 51575 7092 51580
rect 7886 51575 7938 51580
rect 8010 51575 8062 51580
rect 8134 51575 8186 51580
rect 8258 51575 8310 51580
rect 8382 51575 8434 51580
rect 8506 51575 8558 51580
rect 8630 51575 8682 51580
rect 8754 51575 8806 51580
rect 8878 51575 8930 51580
rect 9002 51575 9054 51580
rect 9126 51575 9178 51580
rect 9250 51575 9302 51580
rect 9374 51575 9426 51580
rect 9498 51575 9550 51580
rect 9622 51575 9674 51580
rect 9746 51575 9798 51580
rect 10251 51575 10303 51580
rect 10375 51575 10427 51580
rect 10499 51575 10551 51580
rect 10623 51575 10675 51580
rect 10747 51575 10799 51580
rect 10871 51575 10923 51580
rect 10995 51575 11047 51580
rect 11119 51575 11171 51580
rect 11243 51575 11295 51580
rect 11367 51575 11419 51580
rect 3559 51498 3611 51503
rect 3683 51498 3735 51503
rect 3807 51498 3859 51503
rect 3931 51498 3983 51503
rect 4055 51498 4107 51503
rect 4179 51498 4231 51503
rect 4303 51498 4355 51503
rect 4427 51498 4479 51503
rect 4551 51498 4603 51503
rect 4675 51498 4727 51503
rect 5180 51498 5232 51503
rect 5304 51498 5356 51503
rect 5428 51498 5480 51503
rect 5552 51498 5604 51503
rect 5676 51498 5728 51503
rect 5800 51498 5852 51503
rect 5924 51498 5976 51503
rect 6048 51498 6100 51503
rect 6172 51498 6224 51503
rect 6296 51498 6348 51503
rect 6420 51498 6472 51503
rect 6544 51498 6596 51503
rect 6668 51498 6720 51503
rect 6792 51498 6844 51503
rect 6916 51498 6968 51503
rect 7040 51498 7092 51503
rect 7886 51498 7938 51503
rect 8010 51498 8062 51503
rect 8134 51498 8186 51503
rect 8258 51498 8310 51503
rect 8382 51498 8434 51503
rect 8506 51498 8558 51503
rect 8630 51498 8682 51503
rect 8754 51498 8806 51503
rect 8878 51498 8930 51503
rect 9002 51498 9054 51503
rect 9126 51498 9178 51503
rect 9250 51498 9302 51503
rect 9374 51498 9426 51503
rect 9498 51498 9550 51503
rect 9622 51498 9674 51503
rect 9746 51498 9798 51503
rect 10251 51498 10303 51503
rect 10375 51498 10427 51503
rect 10499 51498 10551 51503
rect 10623 51498 10675 51503
rect 10747 51498 10799 51503
rect 10871 51498 10923 51503
rect 10995 51498 11047 51503
rect 11119 51498 11171 51503
rect 11243 51498 11295 51503
rect 11367 51498 11419 51503
rect 3559 51452 3611 51498
rect 3683 51452 3735 51498
rect 3807 51452 3859 51498
rect 3931 51452 3983 51498
rect 4055 51452 4107 51498
rect 4179 51452 4231 51498
rect 4303 51452 4355 51498
rect 4427 51452 4479 51498
rect 4551 51452 4603 51498
rect 4675 51452 4727 51498
rect 5180 51452 5232 51498
rect 5304 51452 5356 51498
rect 5428 51452 5480 51498
rect 5552 51452 5604 51498
rect 5676 51452 5728 51498
rect 5800 51452 5852 51498
rect 5924 51452 5976 51498
rect 6048 51452 6100 51498
rect 6172 51452 6224 51498
rect 6296 51452 6348 51498
rect 6420 51452 6472 51498
rect 6544 51452 6596 51498
rect 6668 51452 6720 51498
rect 6792 51452 6844 51498
rect 6916 51452 6968 51498
rect 7040 51452 7092 51498
rect 7886 51452 7938 51498
rect 8010 51452 8062 51498
rect 8134 51452 8186 51498
rect 8258 51452 8310 51498
rect 8382 51452 8434 51498
rect 8506 51452 8558 51498
rect 8630 51452 8682 51498
rect 8754 51452 8806 51498
rect 8878 51452 8930 51498
rect 9002 51452 9054 51498
rect 9126 51452 9178 51498
rect 9250 51452 9302 51498
rect 9374 51452 9426 51498
rect 9498 51452 9550 51498
rect 9622 51452 9674 51498
rect 9746 51452 9798 51498
rect 10251 51452 10303 51498
rect 10375 51452 10427 51498
rect 10499 51452 10551 51498
rect 10623 51452 10675 51498
rect 10747 51452 10799 51498
rect 10871 51452 10923 51498
rect 10995 51452 11047 51498
rect 11119 51452 11171 51498
rect 11243 51452 11295 51498
rect 11367 51452 11419 51498
rect 3559 51451 3611 51452
rect 3683 51451 3735 51452
rect 3807 51451 3859 51452
rect 3931 51451 3983 51452
rect 4055 51451 4107 51452
rect 4179 51451 4231 51452
rect 4303 51451 4355 51452
rect 4427 51451 4479 51452
rect 4551 51451 4603 51452
rect 4675 51451 4727 51452
rect 5180 51451 5232 51452
rect 5304 51451 5356 51452
rect 5428 51451 5480 51452
rect 5552 51451 5604 51452
rect 5676 51451 5728 51452
rect 5800 51451 5852 51452
rect 5924 51451 5976 51452
rect 6048 51451 6100 51452
rect 6172 51451 6224 51452
rect 6296 51451 6348 51452
rect 6420 51451 6472 51452
rect 6544 51451 6596 51452
rect 6668 51451 6720 51452
rect 6792 51451 6844 51452
rect 6916 51451 6968 51452
rect 7040 51451 7092 51452
rect 7886 51451 7938 51452
rect 8010 51451 8062 51452
rect 8134 51451 8186 51452
rect 8258 51451 8310 51452
rect 8382 51451 8434 51452
rect 8506 51451 8558 51452
rect 8630 51451 8682 51452
rect 8754 51451 8806 51452
rect 8878 51451 8930 51452
rect 9002 51451 9054 51452
rect 9126 51451 9178 51452
rect 9250 51451 9302 51452
rect 9374 51451 9426 51452
rect 9498 51451 9550 51452
rect 9622 51451 9674 51452
rect 9746 51451 9798 51452
rect 10251 51451 10303 51452
rect 10375 51451 10427 51452
rect 10499 51451 10551 51452
rect 10623 51451 10675 51452
rect 10747 51451 10799 51452
rect 10871 51451 10923 51452
rect 10995 51451 11047 51452
rect 11119 51451 11171 51452
rect 11243 51451 11295 51452
rect 11367 51451 11419 51452
rect 4863 51203 4915 51222
rect 4987 51203 5039 51222
rect 7277 51203 7329 51222
rect 7401 51203 7453 51222
rect 7525 51203 7577 51222
rect 7649 51203 7701 51222
rect 9939 51203 9991 51222
rect 10063 51203 10115 51222
rect 4863 51170 4915 51203
rect 4987 51170 5039 51203
rect 7277 51170 7329 51203
rect 7401 51170 7453 51203
rect 7525 51170 7577 51203
rect 7649 51170 7701 51203
rect 9939 51170 9991 51203
rect 10063 51170 10115 51203
rect 4863 51095 4915 51098
rect 4987 51095 5039 51098
rect 7277 51095 7329 51098
rect 7401 51095 7453 51098
rect 7525 51095 7577 51098
rect 7649 51095 7701 51098
rect 9939 51095 9991 51098
rect 10063 51095 10115 51098
rect 4863 51049 4915 51095
rect 4987 51049 5039 51095
rect 7277 51049 7329 51095
rect 7401 51049 7453 51095
rect 7525 51049 7577 51095
rect 7649 51049 7701 51095
rect 9939 51049 9991 51095
rect 10063 51049 10115 51095
rect 4863 51046 4915 51049
rect 4987 51046 5039 51049
rect 7277 51046 7329 51049
rect 7401 51046 7453 51049
rect 7525 51046 7577 51049
rect 7649 51046 7701 51049
rect 9939 51046 9991 51049
rect 10063 51046 10115 51049
rect 4863 50941 4915 50974
rect 4987 50941 5039 50974
rect 7277 50941 7329 50974
rect 7401 50941 7453 50974
rect 7525 50941 7577 50974
rect 7649 50941 7701 50974
rect 9939 50941 9991 50974
rect 10063 50941 10115 50974
rect 4863 50922 4915 50941
rect 4987 50922 5039 50941
rect 7277 50922 7329 50941
rect 7401 50922 7453 50941
rect 7525 50922 7577 50941
rect 7649 50922 7701 50941
rect 9939 50922 9991 50941
rect 10063 50922 10115 50941
rect 3559 50692 3611 50693
rect 3683 50692 3735 50693
rect 3807 50692 3859 50693
rect 3931 50692 3983 50693
rect 4055 50692 4107 50693
rect 4179 50692 4231 50693
rect 4303 50692 4355 50693
rect 4427 50692 4479 50693
rect 4551 50692 4603 50693
rect 4675 50692 4727 50693
rect 5180 50692 5232 50693
rect 5304 50692 5356 50693
rect 5428 50692 5480 50693
rect 5552 50692 5604 50693
rect 5676 50692 5728 50693
rect 5800 50692 5852 50693
rect 5924 50692 5976 50693
rect 6048 50692 6100 50693
rect 6172 50692 6224 50693
rect 6296 50692 6348 50693
rect 6420 50692 6472 50693
rect 6544 50692 6596 50693
rect 6668 50692 6720 50693
rect 6792 50692 6844 50693
rect 6916 50692 6968 50693
rect 7040 50692 7092 50693
rect 7886 50692 7938 50693
rect 8010 50692 8062 50693
rect 8134 50692 8186 50693
rect 8258 50692 8310 50693
rect 8382 50692 8434 50693
rect 8506 50692 8558 50693
rect 8630 50692 8682 50693
rect 8754 50692 8806 50693
rect 8878 50692 8930 50693
rect 9002 50692 9054 50693
rect 9126 50692 9178 50693
rect 9250 50692 9302 50693
rect 9374 50692 9426 50693
rect 9498 50692 9550 50693
rect 9622 50692 9674 50693
rect 9746 50692 9798 50693
rect 10251 50692 10303 50693
rect 10375 50692 10427 50693
rect 10499 50692 10551 50693
rect 10623 50692 10675 50693
rect 10747 50692 10799 50693
rect 10871 50692 10923 50693
rect 10995 50692 11047 50693
rect 11119 50692 11171 50693
rect 11243 50692 11295 50693
rect 11367 50692 11419 50693
rect 3559 50646 3611 50692
rect 3683 50646 3735 50692
rect 3807 50646 3859 50692
rect 3931 50646 3983 50692
rect 4055 50646 4107 50692
rect 4179 50646 4231 50692
rect 4303 50646 4355 50692
rect 4427 50646 4479 50692
rect 4551 50646 4603 50692
rect 4675 50646 4727 50692
rect 5180 50646 5232 50692
rect 5304 50646 5356 50692
rect 5428 50646 5480 50692
rect 5552 50646 5604 50692
rect 5676 50646 5728 50692
rect 5800 50646 5852 50692
rect 5924 50646 5976 50692
rect 6048 50646 6100 50692
rect 6172 50646 6224 50692
rect 6296 50646 6348 50692
rect 6420 50646 6472 50692
rect 6544 50646 6596 50692
rect 6668 50646 6720 50692
rect 6792 50646 6844 50692
rect 6916 50646 6968 50692
rect 7040 50646 7092 50692
rect 7886 50646 7938 50692
rect 8010 50646 8062 50692
rect 8134 50646 8186 50692
rect 8258 50646 8310 50692
rect 8382 50646 8434 50692
rect 8506 50646 8558 50692
rect 8630 50646 8682 50692
rect 8754 50646 8806 50692
rect 8878 50646 8930 50692
rect 9002 50646 9054 50692
rect 9126 50646 9178 50692
rect 9250 50646 9302 50692
rect 9374 50646 9426 50692
rect 9498 50646 9550 50692
rect 9622 50646 9674 50692
rect 9746 50646 9798 50692
rect 10251 50646 10303 50692
rect 10375 50646 10427 50692
rect 10499 50646 10551 50692
rect 10623 50646 10675 50692
rect 10747 50646 10799 50692
rect 10871 50646 10923 50692
rect 10995 50646 11047 50692
rect 11119 50646 11171 50692
rect 11243 50646 11295 50692
rect 11367 50646 11419 50692
rect 3559 50641 3611 50646
rect 3683 50641 3735 50646
rect 3807 50641 3859 50646
rect 3931 50641 3983 50646
rect 4055 50641 4107 50646
rect 4179 50641 4231 50646
rect 4303 50641 4355 50646
rect 4427 50641 4479 50646
rect 4551 50641 4603 50646
rect 4675 50641 4727 50646
rect 5180 50641 5232 50646
rect 5304 50641 5356 50646
rect 5428 50641 5480 50646
rect 5552 50641 5604 50646
rect 5676 50641 5728 50646
rect 5800 50641 5852 50646
rect 5924 50641 5976 50646
rect 6048 50641 6100 50646
rect 6172 50641 6224 50646
rect 6296 50641 6348 50646
rect 6420 50641 6472 50646
rect 6544 50641 6596 50646
rect 6668 50641 6720 50646
rect 6792 50641 6844 50646
rect 6916 50641 6968 50646
rect 7040 50641 7092 50646
rect 7886 50641 7938 50646
rect 8010 50641 8062 50646
rect 8134 50641 8186 50646
rect 8258 50641 8310 50646
rect 8382 50641 8434 50646
rect 8506 50641 8558 50646
rect 8630 50641 8682 50646
rect 8754 50641 8806 50646
rect 8878 50641 8930 50646
rect 9002 50641 9054 50646
rect 9126 50641 9178 50646
rect 9250 50641 9302 50646
rect 9374 50641 9426 50646
rect 9498 50641 9550 50646
rect 9622 50641 9674 50646
rect 9746 50641 9798 50646
rect 10251 50641 10303 50646
rect 10375 50641 10427 50646
rect 10499 50641 10551 50646
rect 10623 50641 10675 50646
rect 10747 50641 10799 50646
rect 10871 50641 10923 50646
rect 10995 50641 11047 50646
rect 11119 50641 11171 50646
rect 11243 50641 11295 50646
rect 11367 50641 11419 50646
rect 3559 50564 3611 50569
rect 3683 50564 3735 50569
rect 3807 50564 3859 50569
rect 3931 50564 3983 50569
rect 4055 50564 4107 50569
rect 4179 50564 4231 50569
rect 4303 50564 4355 50569
rect 4427 50564 4479 50569
rect 4551 50564 4603 50569
rect 4675 50564 4727 50569
rect 5180 50564 5232 50569
rect 5304 50564 5356 50569
rect 5428 50564 5480 50569
rect 5552 50564 5604 50569
rect 5676 50564 5728 50569
rect 5800 50564 5852 50569
rect 5924 50564 5976 50569
rect 6048 50564 6100 50569
rect 6172 50564 6224 50569
rect 6296 50564 6348 50569
rect 6420 50564 6472 50569
rect 6544 50564 6596 50569
rect 6668 50564 6720 50569
rect 6792 50564 6844 50569
rect 6916 50564 6968 50569
rect 7040 50564 7092 50569
rect 7886 50564 7938 50569
rect 8010 50564 8062 50569
rect 8134 50564 8186 50569
rect 8258 50564 8310 50569
rect 8382 50564 8434 50569
rect 8506 50564 8558 50569
rect 8630 50564 8682 50569
rect 8754 50564 8806 50569
rect 8878 50564 8930 50569
rect 9002 50564 9054 50569
rect 9126 50564 9178 50569
rect 9250 50564 9302 50569
rect 9374 50564 9426 50569
rect 9498 50564 9550 50569
rect 9622 50564 9674 50569
rect 9746 50564 9798 50569
rect 10251 50564 10303 50569
rect 10375 50564 10427 50569
rect 10499 50564 10551 50569
rect 10623 50564 10675 50569
rect 10747 50564 10799 50569
rect 10871 50564 10923 50569
rect 10995 50564 11047 50569
rect 11119 50564 11171 50569
rect 11243 50564 11295 50569
rect 11367 50564 11419 50569
rect 3559 50518 3611 50564
rect 3683 50518 3735 50564
rect 3807 50518 3859 50564
rect 3931 50518 3983 50564
rect 4055 50518 4107 50564
rect 4179 50518 4231 50564
rect 4303 50518 4355 50564
rect 4427 50518 4479 50564
rect 4551 50518 4603 50564
rect 4675 50518 4727 50564
rect 5180 50518 5232 50564
rect 5304 50518 5356 50564
rect 5428 50518 5480 50564
rect 5552 50518 5604 50564
rect 5676 50518 5728 50564
rect 5800 50518 5852 50564
rect 5924 50518 5976 50564
rect 6048 50518 6100 50564
rect 6172 50518 6224 50564
rect 6296 50518 6348 50564
rect 6420 50518 6472 50564
rect 6544 50518 6596 50564
rect 6668 50518 6720 50564
rect 6792 50518 6844 50564
rect 6916 50518 6968 50564
rect 7040 50518 7092 50564
rect 7886 50518 7938 50564
rect 8010 50518 8062 50564
rect 8134 50518 8186 50564
rect 8258 50518 8310 50564
rect 8382 50518 8434 50564
rect 8506 50518 8558 50564
rect 8630 50518 8682 50564
rect 8754 50518 8806 50564
rect 8878 50518 8930 50564
rect 9002 50518 9054 50564
rect 9126 50518 9178 50564
rect 9250 50518 9302 50564
rect 9374 50518 9426 50564
rect 9498 50518 9550 50564
rect 9622 50518 9674 50564
rect 9746 50518 9798 50564
rect 10251 50518 10303 50564
rect 10375 50518 10427 50564
rect 10499 50518 10551 50564
rect 10623 50518 10675 50564
rect 10747 50518 10799 50564
rect 10871 50518 10923 50564
rect 10995 50518 11047 50564
rect 11119 50518 11171 50564
rect 11243 50518 11295 50564
rect 11367 50518 11419 50564
rect 3559 50517 3611 50518
rect 3683 50517 3735 50518
rect 3807 50517 3859 50518
rect 3931 50517 3983 50518
rect 4055 50517 4107 50518
rect 4179 50517 4231 50518
rect 4303 50517 4355 50518
rect 4427 50517 4479 50518
rect 4551 50517 4603 50518
rect 4675 50517 4727 50518
rect 5180 50517 5232 50518
rect 5304 50517 5356 50518
rect 5428 50517 5480 50518
rect 5552 50517 5604 50518
rect 5676 50517 5728 50518
rect 5800 50517 5852 50518
rect 5924 50517 5976 50518
rect 6048 50517 6100 50518
rect 6172 50517 6224 50518
rect 6296 50517 6348 50518
rect 6420 50517 6472 50518
rect 6544 50517 6596 50518
rect 6668 50517 6720 50518
rect 6792 50517 6844 50518
rect 6916 50517 6968 50518
rect 7040 50517 7092 50518
rect 7886 50517 7938 50518
rect 8010 50517 8062 50518
rect 8134 50517 8186 50518
rect 8258 50517 8310 50518
rect 8382 50517 8434 50518
rect 8506 50517 8558 50518
rect 8630 50517 8682 50518
rect 8754 50517 8806 50518
rect 8878 50517 8930 50518
rect 9002 50517 9054 50518
rect 9126 50517 9178 50518
rect 9250 50517 9302 50518
rect 9374 50517 9426 50518
rect 9498 50517 9550 50518
rect 9622 50517 9674 50518
rect 9746 50517 9798 50518
rect 10251 50517 10303 50518
rect 10375 50517 10427 50518
rect 10499 50517 10551 50518
rect 10623 50517 10675 50518
rect 10747 50517 10799 50518
rect 10871 50517 10923 50518
rect 10995 50517 11047 50518
rect 11119 50517 11171 50518
rect 11243 50517 11295 50518
rect 11367 50517 11419 50518
rect 4863 50269 4915 50288
rect 4987 50269 5039 50288
rect 7277 50269 7329 50288
rect 7401 50269 7453 50288
rect 7525 50269 7577 50288
rect 7649 50269 7701 50288
rect 9939 50269 9991 50288
rect 10063 50269 10115 50288
rect 4863 50236 4915 50269
rect 4987 50236 5039 50269
rect 7277 50236 7329 50269
rect 7401 50236 7453 50269
rect 7525 50236 7577 50269
rect 7649 50236 7701 50269
rect 9939 50236 9991 50269
rect 10063 50236 10115 50269
rect 4863 50161 4915 50164
rect 4987 50161 5039 50164
rect 7277 50161 7329 50164
rect 7401 50161 7453 50164
rect 7525 50161 7577 50164
rect 7649 50161 7701 50164
rect 9939 50161 9991 50164
rect 10063 50161 10115 50164
rect 4863 50115 4915 50161
rect 4987 50115 5039 50161
rect 7277 50115 7329 50161
rect 7401 50115 7453 50161
rect 7525 50115 7577 50161
rect 7649 50115 7701 50161
rect 9939 50115 9991 50161
rect 10063 50115 10115 50161
rect 4863 50112 4915 50115
rect 4987 50112 5039 50115
rect 7277 50112 7329 50115
rect 7401 50112 7453 50115
rect 7525 50112 7577 50115
rect 7649 50112 7701 50115
rect 9939 50112 9991 50115
rect 10063 50112 10115 50115
rect 4863 50007 4915 50040
rect 4987 50007 5039 50040
rect 7277 50007 7329 50040
rect 7401 50007 7453 50040
rect 7525 50007 7577 50040
rect 7649 50007 7701 50040
rect 9939 50007 9991 50040
rect 10063 50007 10115 50040
rect 4863 49988 4915 50007
rect 4987 49988 5039 50007
rect 7277 49988 7329 50007
rect 7401 49988 7453 50007
rect 7525 49988 7577 50007
rect 7649 49988 7701 50007
rect 9939 49988 9991 50007
rect 10063 49988 10115 50007
rect 3559 49758 3611 49759
rect 3683 49758 3735 49759
rect 3807 49758 3859 49759
rect 3931 49758 3983 49759
rect 4055 49758 4107 49759
rect 4179 49758 4231 49759
rect 4303 49758 4355 49759
rect 4427 49758 4479 49759
rect 4551 49758 4603 49759
rect 4675 49758 4727 49759
rect 5180 49758 5232 49759
rect 5304 49758 5356 49759
rect 5428 49758 5480 49759
rect 5552 49758 5604 49759
rect 5676 49758 5728 49759
rect 5800 49758 5852 49759
rect 5924 49758 5976 49759
rect 6048 49758 6100 49759
rect 6172 49758 6224 49759
rect 6296 49758 6348 49759
rect 6420 49758 6472 49759
rect 6544 49758 6596 49759
rect 6668 49758 6720 49759
rect 6792 49758 6844 49759
rect 6916 49758 6968 49759
rect 7040 49758 7092 49759
rect 7886 49758 7938 49759
rect 8010 49758 8062 49759
rect 8134 49758 8186 49759
rect 8258 49758 8310 49759
rect 8382 49758 8434 49759
rect 8506 49758 8558 49759
rect 8630 49758 8682 49759
rect 8754 49758 8806 49759
rect 8878 49758 8930 49759
rect 9002 49758 9054 49759
rect 9126 49758 9178 49759
rect 9250 49758 9302 49759
rect 9374 49758 9426 49759
rect 9498 49758 9550 49759
rect 9622 49758 9674 49759
rect 9746 49758 9798 49759
rect 10251 49758 10303 49759
rect 10375 49758 10427 49759
rect 10499 49758 10551 49759
rect 10623 49758 10675 49759
rect 10747 49758 10799 49759
rect 10871 49758 10923 49759
rect 10995 49758 11047 49759
rect 11119 49758 11171 49759
rect 11243 49758 11295 49759
rect 11367 49758 11419 49759
rect 3559 49712 3611 49758
rect 3683 49712 3735 49758
rect 3807 49712 3859 49758
rect 3931 49712 3983 49758
rect 4055 49712 4107 49758
rect 4179 49712 4231 49758
rect 4303 49712 4355 49758
rect 4427 49712 4479 49758
rect 4551 49712 4603 49758
rect 4675 49712 4727 49758
rect 5180 49712 5232 49758
rect 5304 49712 5356 49758
rect 5428 49712 5480 49758
rect 5552 49712 5604 49758
rect 5676 49712 5728 49758
rect 5800 49712 5852 49758
rect 5924 49712 5976 49758
rect 6048 49712 6100 49758
rect 6172 49712 6224 49758
rect 6296 49712 6348 49758
rect 6420 49712 6472 49758
rect 6544 49712 6596 49758
rect 6668 49712 6720 49758
rect 6792 49712 6844 49758
rect 6916 49712 6968 49758
rect 7040 49712 7092 49758
rect 7886 49712 7938 49758
rect 8010 49712 8062 49758
rect 8134 49712 8186 49758
rect 8258 49712 8310 49758
rect 8382 49712 8434 49758
rect 8506 49712 8558 49758
rect 8630 49712 8682 49758
rect 8754 49712 8806 49758
rect 8878 49712 8930 49758
rect 9002 49712 9054 49758
rect 9126 49712 9178 49758
rect 9250 49712 9302 49758
rect 9374 49712 9426 49758
rect 9498 49712 9550 49758
rect 9622 49712 9674 49758
rect 9746 49712 9798 49758
rect 10251 49712 10303 49758
rect 10375 49712 10427 49758
rect 10499 49712 10551 49758
rect 10623 49712 10675 49758
rect 10747 49712 10799 49758
rect 10871 49712 10923 49758
rect 10995 49712 11047 49758
rect 11119 49712 11171 49758
rect 11243 49712 11295 49758
rect 11367 49712 11419 49758
rect 3559 49707 3611 49712
rect 3683 49707 3735 49712
rect 3807 49707 3859 49712
rect 3931 49707 3983 49712
rect 4055 49707 4107 49712
rect 4179 49707 4231 49712
rect 4303 49707 4355 49712
rect 4427 49707 4479 49712
rect 4551 49707 4603 49712
rect 4675 49707 4727 49712
rect 5180 49707 5232 49712
rect 5304 49707 5356 49712
rect 5428 49707 5480 49712
rect 5552 49707 5604 49712
rect 5676 49707 5728 49712
rect 5800 49707 5852 49712
rect 5924 49707 5976 49712
rect 6048 49707 6100 49712
rect 6172 49707 6224 49712
rect 6296 49707 6348 49712
rect 6420 49707 6472 49712
rect 6544 49707 6596 49712
rect 6668 49707 6720 49712
rect 6792 49707 6844 49712
rect 6916 49707 6968 49712
rect 7040 49707 7092 49712
rect 7886 49707 7938 49712
rect 8010 49707 8062 49712
rect 8134 49707 8186 49712
rect 8258 49707 8310 49712
rect 8382 49707 8434 49712
rect 8506 49707 8558 49712
rect 8630 49707 8682 49712
rect 8754 49707 8806 49712
rect 8878 49707 8930 49712
rect 9002 49707 9054 49712
rect 9126 49707 9178 49712
rect 9250 49707 9302 49712
rect 9374 49707 9426 49712
rect 9498 49707 9550 49712
rect 9622 49707 9674 49712
rect 9746 49707 9798 49712
rect 10251 49707 10303 49712
rect 10375 49707 10427 49712
rect 10499 49707 10551 49712
rect 10623 49707 10675 49712
rect 10747 49707 10799 49712
rect 10871 49707 10923 49712
rect 10995 49707 11047 49712
rect 11119 49707 11171 49712
rect 11243 49707 11295 49712
rect 11367 49707 11419 49712
rect 3559 49630 3611 49635
rect 3683 49630 3735 49635
rect 3807 49630 3859 49635
rect 3931 49630 3983 49635
rect 4055 49630 4107 49635
rect 4179 49630 4231 49635
rect 4303 49630 4355 49635
rect 4427 49630 4479 49635
rect 4551 49630 4603 49635
rect 4675 49630 4727 49635
rect 5180 49630 5232 49635
rect 5304 49630 5356 49635
rect 5428 49630 5480 49635
rect 5552 49630 5604 49635
rect 5676 49630 5728 49635
rect 5800 49630 5852 49635
rect 5924 49630 5976 49635
rect 6048 49630 6100 49635
rect 6172 49630 6224 49635
rect 6296 49630 6348 49635
rect 6420 49630 6472 49635
rect 6544 49630 6596 49635
rect 6668 49630 6720 49635
rect 6792 49630 6844 49635
rect 6916 49630 6968 49635
rect 7040 49630 7092 49635
rect 7886 49630 7938 49635
rect 8010 49630 8062 49635
rect 8134 49630 8186 49635
rect 8258 49630 8310 49635
rect 8382 49630 8434 49635
rect 8506 49630 8558 49635
rect 8630 49630 8682 49635
rect 8754 49630 8806 49635
rect 8878 49630 8930 49635
rect 9002 49630 9054 49635
rect 9126 49630 9178 49635
rect 9250 49630 9302 49635
rect 9374 49630 9426 49635
rect 9498 49630 9550 49635
rect 9622 49630 9674 49635
rect 9746 49630 9798 49635
rect 10251 49630 10303 49635
rect 10375 49630 10427 49635
rect 10499 49630 10551 49635
rect 10623 49630 10675 49635
rect 10747 49630 10799 49635
rect 10871 49630 10923 49635
rect 10995 49630 11047 49635
rect 11119 49630 11171 49635
rect 11243 49630 11295 49635
rect 11367 49630 11419 49635
rect 3559 49584 3611 49630
rect 3683 49584 3735 49630
rect 3807 49584 3859 49630
rect 3931 49584 3983 49630
rect 4055 49584 4107 49630
rect 4179 49584 4231 49630
rect 4303 49584 4355 49630
rect 4427 49584 4479 49630
rect 4551 49584 4603 49630
rect 4675 49584 4727 49630
rect 5180 49584 5232 49630
rect 5304 49584 5356 49630
rect 5428 49584 5480 49630
rect 5552 49584 5604 49630
rect 5676 49584 5728 49630
rect 5800 49584 5852 49630
rect 5924 49584 5976 49630
rect 6048 49584 6100 49630
rect 6172 49584 6224 49630
rect 6296 49584 6348 49630
rect 6420 49584 6472 49630
rect 6544 49584 6596 49630
rect 6668 49584 6720 49630
rect 6792 49584 6844 49630
rect 6916 49584 6968 49630
rect 7040 49584 7092 49630
rect 7886 49584 7938 49630
rect 8010 49584 8062 49630
rect 8134 49584 8186 49630
rect 8258 49584 8310 49630
rect 8382 49584 8434 49630
rect 8506 49584 8558 49630
rect 8630 49584 8682 49630
rect 8754 49584 8806 49630
rect 8878 49584 8930 49630
rect 9002 49584 9054 49630
rect 9126 49584 9178 49630
rect 9250 49584 9302 49630
rect 9374 49584 9426 49630
rect 9498 49584 9550 49630
rect 9622 49584 9674 49630
rect 9746 49584 9798 49630
rect 10251 49584 10303 49630
rect 10375 49584 10427 49630
rect 10499 49584 10551 49630
rect 10623 49584 10675 49630
rect 10747 49584 10799 49630
rect 10871 49584 10923 49630
rect 10995 49584 11047 49630
rect 11119 49584 11171 49630
rect 11243 49584 11295 49630
rect 11367 49584 11419 49630
rect 3559 49583 3611 49584
rect 3683 49583 3735 49584
rect 3807 49583 3859 49584
rect 3931 49583 3983 49584
rect 4055 49583 4107 49584
rect 4179 49583 4231 49584
rect 4303 49583 4355 49584
rect 4427 49583 4479 49584
rect 4551 49583 4603 49584
rect 4675 49583 4727 49584
rect 5180 49583 5232 49584
rect 5304 49583 5356 49584
rect 5428 49583 5480 49584
rect 5552 49583 5604 49584
rect 5676 49583 5728 49584
rect 5800 49583 5852 49584
rect 5924 49583 5976 49584
rect 6048 49583 6100 49584
rect 6172 49583 6224 49584
rect 6296 49583 6348 49584
rect 6420 49583 6472 49584
rect 6544 49583 6596 49584
rect 6668 49583 6720 49584
rect 6792 49583 6844 49584
rect 6916 49583 6968 49584
rect 7040 49583 7092 49584
rect 7886 49583 7938 49584
rect 8010 49583 8062 49584
rect 8134 49583 8186 49584
rect 8258 49583 8310 49584
rect 8382 49583 8434 49584
rect 8506 49583 8558 49584
rect 8630 49583 8682 49584
rect 8754 49583 8806 49584
rect 8878 49583 8930 49584
rect 9002 49583 9054 49584
rect 9126 49583 9178 49584
rect 9250 49583 9302 49584
rect 9374 49583 9426 49584
rect 9498 49583 9550 49584
rect 9622 49583 9674 49584
rect 9746 49583 9798 49584
rect 10251 49583 10303 49584
rect 10375 49583 10427 49584
rect 10499 49583 10551 49584
rect 10623 49583 10675 49584
rect 10747 49583 10799 49584
rect 10871 49583 10923 49584
rect 10995 49583 11047 49584
rect 11119 49583 11171 49584
rect 11243 49583 11295 49584
rect 11367 49583 11419 49584
rect 4863 49335 4915 49354
rect 4987 49335 5039 49354
rect 7277 49335 7329 49354
rect 7401 49335 7453 49354
rect 7525 49335 7577 49354
rect 7649 49335 7701 49354
rect 9939 49335 9991 49354
rect 10063 49335 10115 49354
rect 4863 49302 4915 49335
rect 4987 49302 5039 49335
rect 7277 49302 7329 49335
rect 7401 49302 7453 49335
rect 7525 49302 7577 49335
rect 7649 49302 7701 49335
rect 9939 49302 9991 49335
rect 10063 49302 10115 49335
rect 4863 49227 4915 49230
rect 4987 49227 5039 49230
rect 7277 49227 7329 49230
rect 7401 49227 7453 49230
rect 7525 49227 7577 49230
rect 7649 49227 7701 49230
rect 9939 49227 9991 49230
rect 10063 49227 10115 49230
rect 4863 49181 4915 49227
rect 4987 49181 5039 49227
rect 7277 49181 7329 49227
rect 7401 49181 7453 49227
rect 7525 49181 7577 49227
rect 7649 49181 7701 49227
rect 9939 49181 9991 49227
rect 10063 49181 10115 49227
rect 4863 49178 4915 49181
rect 4987 49178 5039 49181
rect 7277 49178 7329 49181
rect 7401 49178 7453 49181
rect 7525 49178 7577 49181
rect 7649 49178 7701 49181
rect 9939 49178 9991 49181
rect 10063 49178 10115 49181
rect 4863 49073 4915 49106
rect 4987 49073 5039 49106
rect 7277 49073 7329 49106
rect 7401 49073 7453 49106
rect 7525 49073 7577 49106
rect 7649 49073 7701 49106
rect 9939 49073 9991 49106
rect 10063 49073 10115 49106
rect 4863 49054 4915 49073
rect 4987 49054 5039 49073
rect 7277 49054 7329 49073
rect 7401 49054 7453 49073
rect 7525 49054 7577 49073
rect 7649 49054 7701 49073
rect 9939 49054 9991 49073
rect 10063 49054 10115 49073
rect 3559 48824 3611 48825
rect 3683 48824 3735 48825
rect 3807 48824 3859 48825
rect 3931 48824 3983 48825
rect 4055 48824 4107 48825
rect 4179 48824 4231 48825
rect 4303 48824 4355 48825
rect 4427 48824 4479 48825
rect 4551 48824 4603 48825
rect 4675 48824 4727 48825
rect 5180 48824 5232 48825
rect 5304 48824 5356 48825
rect 5428 48824 5480 48825
rect 5552 48824 5604 48825
rect 5676 48824 5728 48825
rect 5800 48824 5852 48825
rect 5924 48824 5976 48825
rect 6048 48824 6100 48825
rect 6172 48824 6224 48825
rect 6296 48824 6348 48825
rect 6420 48824 6472 48825
rect 6544 48824 6596 48825
rect 6668 48824 6720 48825
rect 6792 48824 6844 48825
rect 6916 48824 6968 48825
rect 7040 48824 7092 48825
rect 7886 48824 7938 48825
rect 8010 48824 8062 48825
rect 8134 48824 8186 48825
rect 8258 48824 8310 48825
rect 8382 48824 8434 48825
rect 8506 48824 8558 48825
rect 8630 48824 8682 48825
rect 8754 48824 8806 48825
rect 8878 48824 8930 48825
rect 9002 48824 9054 48825
rect 9126 48824 9178 48825
rect 9250 48824 9302 48825
rect 9374 48824 9426 48825
rect 9498 48824 9550 48825
rect 9622 48824 9674 48825
rect 9746 48824 9798 48825
rect 10251 48824 10303 48825
rect 10375 48824 10427 48825
rect 10499 48824 10551 48825
rect 10623 48824 10675 48825
rect 10747 48824 10799 48825
rect 10871 48824 10923 48825
rect 10995 48824 11047 48825
rect 11119 48824 11171 48825
rect 11243 48824 11295 48825
rect 11367 48824 11419 48825
rect 3559 48778 3611 48824
rect 3683 48778 3735 48824
rect 3807 48778 3859 48824
rect 3931 48778 3983 48824
rect 4055 48778 4107 48824
rect 4179 48778 4231 48824
rect 4303 48778 4355 48824
rect 4427 48778 4479 48824
rect 4551 48778 4603 48824
rect 4675 48778 4727 48824
rect 5180 48778 5232 48824
rect 5304 48778 5356 48824
rect 5428 48778 5480 48824
rect 5552 48778 5604 48824
rect 5676 48778 5728 48824
rect 5800 48778 5852 48824
rect 5924 48778 5976 48824
rect 6048 48778 6100 48824
rect 6172 48778 6224 48824
rect 6296 48778 6348 48824
rect 6420 48778 6472 48824
rect 6544 48778 6596 48824
rect 6668 48778 6720 48824
rect 6792 48778 6844 48824
rect 6916 48778 6968 48824
rect 7040 48778 7092 48824
rect 7886 48778 7938 48824
rect 8010 48778 8062 48824
rect 8134 48778 8186 48824
rect 8258 48778 8310 48824
rect 8382 48778 8434 48824
rect 8506 48778 8558 48824
rect 8630 48778 8682 48824
rect 8754 48778 8806 48824
rect 8878 48778 8930 48824
rect 9002 48778 9054 48824
rect 9126 48778 9178 48824
rect 9250 48778 9302 48824
rect 9374 48778 9426 48824
rect 9498 48778 9550 48824
rect 9622 48778 9674 48824
rect 9746 48778 9798 48824
rect 10251 48778 10303 48824
rect 10375 48778 10427 48824
rect 10499 48778 10551 48824
rect 10623 48778 10675 48824
rect 10747 48778 10799 48824
rect 10871 48778 10923 48824
rect 10995 48778 11047 48824
rect 11119 48778 11171 48824
rect 11243 48778 11295 48824
rect 11367 48778 11419 48824
rect 3559 48773 3611 48778
rect 3683 48773 3735 48778
rect 3807 48773 3859 48778
rect 3931 48773 3983 48778
rect 4055 48773 4107 48778
rect 4179 48773 4231 48778
rect 4303 48773 4355 48778
rect 4427 48773 4479 48778
rect 4551 48773 4603 48778
rect 4675 48773 4727 48778
rect 5180 48773 5232 48778
rect 5304 48773 5356 48778
rect 5428 48773 5480 48778
rect 5552 48773 5604 48778
rect 5676 48773 5728 48778
rect 5800 48773 5852 48778
rect 5924 48773 5976 48778
rect 6048 48773 6100 48778
rect 6172 48773 6224 48778
rect 6296 48773 6348 48778
rect 6420 48773 6472 48778
rect 6544 48773 6596 48778
rect 6668 48773 6720 48778
rect 6792 48773 6844 48778
rect 6916 48773 6968 48778
rect 7040 48773 7092 48778
rect 7886 48773 7938 48778
rect 8010 48773 8062 48778
rect 8134 48773 8186 48778
rect 8258 48773 8310 48778
rect 8382 48773 8434 48778
rect 8506 48773 8558 48778
rect 8630 48773 8682 48778
rect 8754 48773 8806 48778
rect 8878 48773 8930 48778
rect 9002 48773 9054 48778
rect 9126 48773 9178 48778
rect 9250 48773 9302 48778
rect 9374 48773 9426 48778
rect 9498 48773 9550 48778
rect 9622 48773 9674 48778
rect 9746 48773 9798 48778
rect 10251 48773 10303 48778
rect 10375 48773 10427 48778
rect 10499 48773 10551 48778
rect 10623 48773 10675 48778
rect 10747 48773 10799 48778
rect 10871 48773 10923 48778
rect 10995 48773 11047 48778
rect 11119 48773 11171 48778
rect 11243 48773 11295 48778
rect 11367 48773 11419 48778
rect 3559 48696 3611 48701
rect 3683 48696 3735 48701
rect 3807 48696 3859 48701
rect 3931 48696 3983 48701
rect 4055 48696 4107 48701
rect 4179 48696 4231 48701
rect 4303 48696 4355 48701
rect 4427 48696 4479 48701
rect 4551 48696 4603 48701
rect 4675 48696 4727 48701
rect 5180 48696 5232 48701
rect 5304 48696 5356 48701
rect 5428 48696 5480 48701
rect 5552 48696 5604 48701
rect 5676 48696 5728 48701
rect 5800 48696 5852 48701
rect 5924 48696 5976 48701
rect 6048 48696 6100 48701
rect 6172 48696 6224 48701
rect 6296 48696 6348 48701
rect 6420 48696 6472 48701
rect 6544 48696 6596 48701
rect 6668 48696 6720 48701
rect 6792 48696 6844 48701
rect 6916 48696 6968 48701
rect 7040 48696 7092 48701
rect 7886 48696 7938 48701
rect 8010 48696 8062 48701
rect 8134 48696 8186 48701
rect 8258 48696 8310 48701
rect 8382 48696 8434 48701
rect 8506 48696 8558 48701
rect 8630 48696 8682 48701
rect 8754 48696 8806 48701
rect 8878 48696 8930 48701
rect 9002 48696 9054 48701
rect 9126 48696 9178 48701
rect 9250 48696 9302 48701
rect 9374 48696 9426 48701
rect 9498 48696 9550 48701
rect 9622 48696 9674 48701
rect 9746 48696 9798 48701
rect 10251 48696 10303 48701
rect 10375 48696 10427 48701
rect 10499 48696 10551 48701
rect 10623 48696 10675 48701
rect 10747 48696 10799 48701
rect 10871 48696 10923 48701
rect 10995 48696 11047 48701
rect 11119 48696 11171 48701
rect 11243 48696 11295 48701
rect 11367 48696 11419 48701
rect 3559 48650 3611 48696
rect 3683 48650 3735 48696
rect 3807 48650 3859 48696
rect 3931 48650 3983 48696
rect 4055 48650 4107 48696
rect 4179 48650 4231 48696
rect 4303 48650 4355 48696
rect 4427 48650 4479 48696
rect 4551 48650 4603 48696
rect 4675 48650 4727 48696
rect 5180 48650 5232 48696
rect 5304 48650 5356 48696
rect 5428 48650 5480 48696
rect 5552 48650 5604 48696
rect 5676 48650 5728 48696
rect 5800 48650 5852 48696
rect 5924 48650 5976 48696
rect 6048 48650 6100 48696
rect 6172 48650 6224 48696
rect 6296 48650 6348 48696
rect 6420 48650 6472 48696
rect 6544 48650 6596 48696
rect 6668 48650 6720 48696
rect 6792 48650 6844 48696
rect 6916 48650 6968 48696
rect 7040 48650 7092 48696
rect 7886 48650 7938 48696
rect 8010 48650 8062 48696
rect 8134 48650 8186 48696
rect 8258 48650 8310 48696
rect 8382 48650 8434 48696
rect 8506 48650 8558 48696
rect 8630 48650 8682 48696
rect 8754 48650 8806 48696
rect 8878 48650 8930 48696
rect 9002 48650 9054 48696
rect 9126 48650 9178 48696
rect 9250 48650 9302 48696
rect 9374 48650 9426 48696
rect 9498 48650 9550 48696
rect 9622 48650 9674 48696
rect 9746 48650 9798 48696
rect 10251 48650 10303 48696
rect 10375 48650 10427 48696
rect 10499 48650 10551 48696
rect 10623 48650 10675 48696
rect 10747 48650 10799 48696
rect 10871 48650 10923 48696
rect 10995 48650 11047 48696
rect 11119 48650 11171 48696
rect 11243 48650 11295 48696
rect 11367 48650 11419 48696
rect 3559 48649 3611 48650
rect 3683 48649 3735 48650
rect 3807 48649 3859 48650
rect 3931 48649 3983 48650
rect 4055 48649 4107 48650
rect 4179 48649 4231 48650
rect 4303 48649 4355 48650
rect 4427 48649 4479 48650
rect 4551 48649 4603 48650
rect 4675 48649 4727 48650
rect 5180 48649 5232 48650
rect 5304 48649 5356 48650
rect 5428 48649 5480 48650
rect 5552 48649 5604 48650
rect 5676 48649 5728 48650
rect 5800 48649 5852 48650
rect 5924 48649 5976 48650
rect 6048 48649 6100 48650
rect 6172 48649 6224 48650
rect 6296 48649 6348 48650
rect 6420 48649 6472 48650
rect 6544 48649 6596 48650
rect 6668 48649 6720 48650
rect 6792 48649 6844 48650
rect 6916 48649 6968 48650
rect 7040 48649 7092 48650
rect 7886 48649 7938 48650
rect 8010 48649 8062 48650
rect 8134 48649 8186 48650
rect 8258 48649 8310 48650
rect 8382 48649 8434 48650
rect 8506 48649 8558 48650
rect 8630 48649 8682 48650
rect 8754 48649 8806 48650
rect 8878 48649 8930 48650
rect 9002 48649 9054 48650
rect 9126 48649 9178 48650
rect 9250 48649 9302 48650
rect 9374 48649 9426 48650
rect 9498 48649 9550 48650
rect 9622 48649 9674 48650
rect 9746 48649 9798 48650
rect 10251 48649 10303 48650
rect 10375 48649 10427 48650
rect 10499 48649 10551 48650
rect 10623 48649 10675 48650
rect 10747 48649 10799 48650
rect 10871 48649 10923 48650
rect 10995 48649 11047 48650
rect 11119 48649 11171 48650
rect 11243 48649 11295 48650
rect 11367 48649 11419 48650
rect 4863 48401 4915 48435
rect 4987 48401 5039 48435
rect 7277 48401 7329 48435
rect 7401 48401 7453 48435
rect 7525 48401 7577 48435
rect 7649 48401 7701 48435
rect 9939 48401 9991 48435
rect 10063 48401 10115 48435
rect 4863 48383 4915 48401
rect 4987 48383 5039 48401
rect 7277 48383 7329 48401
rect 7401 48383 7453 48401
rect 7525 48383 7577 48401
rect 7649 48383 7701 48401
rect 9939 48383 9991 48401
rect 10063 48383 10115 48401
rect 4863 48293 4915 48311
rect 4987 48293 5039 48311
rect 7277 48293 7329 48311
rect 7401 48293 7453 48311
rect 7525 48293 7577 48311
rect 7649 48293 7701 48311
rect 9939 48293 9991 48311
rect 10063 48293 10115 48311
rect 4863 48259 4915 48293
rect 4987 48259 5039 48293
rect 7277 48259 7329 48293
rect 7401 48259 7453 48293
rect 7525 48259 7577 48293
rect 7649 48259 7701 48293
rect 9939 48259 9991 48293
rect 10063 48259 10115 48293
rect 2810 47936 2862 47988
rect 2934 47936 2986 47988
rect 3058 47936 3110 47988
rect 3182 47936 3234 47988
rect 3306 47936 3358 47988
rect 3430 47936 3482 47988
rect 3554 47936 3606 47988
rect 3678 47936 3730 47988
rect 3802 47936 3854 47988
rect 3926 47936 3978 47988
rect 4050 47936 4102 47988
rect 4174 47936 4226 47988
rect 4298 47936 4350 47988
rect 4422 47936 4474 47988
rect 4546 47936 4598 47988
rect 4670 47936 4722 47988
rect 5180 47936 5232 47988
rect 5304 47936 5356 47988
rect 5428 47936 5480 47988
rect 5552 47936 5604 47988
rect 5676 47936 5728 47988
rect 5800 47936 5852 47988
rect 5924 47936 5976 47988
rect 6048 47936 6100 47988
rect 6172 47936 6224 47988
rect 6296 47936 6348 47988
rect 6420 47936 6472 47988
rect 6544 47936 6596 47988
rect 6668 47936 6720 47988
rect 6792 47936 6844 47988
rect 6916 47936 6968 47988
rect 7040 47936 7092 47988
rect 7886 47936 7938 47988
rect 8010 47936 8062 47988
rect 8134 47936 8186 47988
rect 8258 47936 8310 47988
rect 8382 47936 8434 47988
rect 8506 47936 8558 47988
rect 8630 47936 8682 47988
rect 8754 47936 8806 47988
rect 8878 47936 8930 47988
rect 9002 47936 9054 47988
rect 9126 47936 9178 47988
rect 9250 47936 9302 47988
rect 9374 47936 9426 47988
rect 9498 47936 9550 47988
rect 9622 47936 9674 47988
rect 9746 47936 9798 47988
rect 10256 47936 10308 47988
rect 10380 47936 10432 47988
rect 10504 47936 10556 47988
rect 10628 47936 10680 47988
rect 10752 47936 10804 47988
rect 10876 47936 10928 47988
rect 11000 47936 11052 47988
rect 11124 47936 11176 47988
rect 11248 47936 11300 47988
rect 11372 47936 11424 47988
rect 11496 47936 11548 47988
rect 11620 47936 11672 47988
rect 11744 47936 11796 47988
rect 11868 47936 11920 47988
rect 11992 47936 12044 47988
rect 12116 47936 12168 47988
rect 2810 47812 2862 47864
rect 2934 47812 2986 47864
rect 3058 47812 3110 47864
rect 3182 47812 3234 47864
rect 3306 47812 3358 47864
rect 3430 47812 3482 47864
rect 3554 47812 3606 47864
rect 3678 47812 3730 47864
rect 3802 47812 3854 47864
rect 3926 47812 3978 47864
rect 4050 47812 4102 47864
rect 4174 47812 4226 47864
rect 4298 47812 4350 47864
rect 4422 47812 4474 47864
rect 4546 47812 4598 47864
rect 4670 47812 4722 47864
rect 5180 47812 5232 47864
rect 5304 47812 5356 47864
rect 5428 47812 5480 47864
rect 5552 47812 5604 47864
rect 5676 47812 5728 47864
rect 5800 47812 5852 47864
rect 5924 47812 5976 47864
rect 6048 47812 6100 47864
rect 6172 47812 6224 47864
rect 6296 47812 6348 47864
rect 6420 47812 6472 47864
rect 6544 47812 6596 47864
rect 6668 47812 6720 47864
rect 6792 47812 6844 47864
rect 6916 47812 6968 47864
rect 7040 47812 7092 47864
rect 7886 47812 7938 47864
rect 8010 47812 8062 47864
rect 8134 47812 8186 47864
rect 8258 47812 8310 47864
rect 8382 47812 8434 47864
rect 8506 47812 8558 47864
rect 8630 47812 8682 47864
rect 8754 47812 8806 47864
rect 8878 47812 8930 47864
rect 9002 47812 9054 47864
rect 9126 47812 9178 47864
rect 9250 47812 9302 47864
rect 9374 47812 9426 47864
rect 9498 47812 9550 47864
rect 9622 47812 9674 47864
rect 9746 47812 9798 47864
rect 10256 47812 10308 47864
rect 10380 47812 10432 47864
rect 10504 47812 10556 47864
rect 10628 47812 10680 47864
rect 10752 47812 10804 47864
rect 10876 47812 10928 47864
rect 11000 47812 11052 47864
rect 11124 47812 11176 47864
rect 11248 47812 11300 47864
rect 11372 47812 11424 47864
rect 11496 47812 11548 47864
rect 11620 47812 11672 47864
rect 11744 47812 11796 47864
rect 11868 47812 11920 47864
rect 11992 47812 12044 47864
rect 12116 47812 12168 47864
rect 2810 47688 2862 47740
rect 2934 47688 2986 47740
rect 3058 47688 3110 47740
rect 3182 47688 3234 47740
rect 3306 47688 3358 47740
rect 3430 47688 3482 47740
rect 3554 47688 3606 47740
rect 3678 47688 3730 47740
rect 3802 47688 3854 47740
rect 3926 47688 3978 47740
rect 4050 47688 4102 47740
rect 4174 47688 4226 47740
rect 4298 47688 4350 47740
rect 4422 47688 4474 47740
rect 4546 47688 4598 47740
rect 4670 47688 4722 47740
rect 5180 47688 5232 47740
rect 5304 47688 5356 47740
rect 5428 47688 5480 47740
rect 5552 47688 5604 47740
rect 5676 47688 5728 47740
rect 5800 47688 5852 47740
rect 5924 47688 5976 47740
rect 6048 47688 6100 47740
rect 6172 47688 6224 47740
rect 6296 47688 6348 47740
rect 6420 47688 6472 47740
rect 6544 47688 6596 47740
rect 6668 47688 6720 47740
rect 6792 47688 6844 47740
rect 6916 47688 6968 47740
rect 7040 47688 7092 47740
rect 7886 47688 7938 47740
rect 8010 47688 8062 47740
rect 8134 47688 8186 47740
rect 8258 47688 8310 47740
rect 8382 47688 8434 47740
rect 8506 47688 8558 47740
rect 8630 47688 8682 47740
rect 8754 47688 8806 47740
rect 8878 47688 8930 47740
rect 9002 47688 9054 47740
rect 9126 47688 9178 47740
rect 9250 47688 9302 47740
rect 9374 47688 9426 47740
rect 9498 47688 9550 47740
rect 9622 47688 9674 47740
rect 9746 47688 9798 47740
rect 10256 47688 10308 47740
rect 10380 47688 10432 47740
rect 10504 47688 10556 47740
rect 10628 47688 10680 47740
rect 10752 47688 10804 47740
rect 10876 47688 10928 47740
rect 11000 47688 11052 47740
rect 11124 47688 11176 47740
rect 11248 47688 11300 47740
rect 11372 47688 11424 47740
rect 11496 47688 11548 47740
rect 11620 47688 11672 47740
rect 11744 47688 11796 47740
rect 11868 47688 11920 47740
rect 11992 47688 12044 47740
rect 12116 47688 12168 47740
rect 14904 52522 14956 52574
rect 14904 52414 14956 52466
rect 14904 52306 14956 52358
rect 14904 52198 14956 52250
rect 14904 52090 14956 52142
rect 14904 51982 14956 52034
rect 14904 51874 14956 51926
rect 14904 51766 14956 51818
rect 14904 51658 14956 51710
rect 14904 51550 14956 51602
rect 14904 51442 14956 51494
rect 14904 51334 14956 51386
rect 14904 51226 14956 51278
rect 22 38122 74 38174
rect 22 38014 74 38066
rect 22 37906 74 37958
rect 22 37798 74 37850
rect 22 37690 74 37742
rect 22 37582 74 37634
rect 22 37474 74 37526
rect 22 37366 74 37418
rect 22 37258 74 37310
rect 22 37150 74 37202
rect 22 37042 74 37094
rect 22 36934 74 36986
rect 22 36826 74 36878
rect 14904 38122 14956 38174
rect 14904 38014 14956 38066
rect 14904 37906 14956 37958
rect 14904 37798 14956 37850
rect 14904 37690 14956 37742
rect 14904 37582 14956 37634
rect 14904 37474 14956 37526
rect 14904 37366 14956 37418
rect 14904 37258 14956 37310
rect 14904 37150 14956 37202
rect 14904 37042 14956 37094
rect 14904 36934 14956 36986
rect 14904 36826 14956 36878
<< metal2 >>
rect 261 56669 2161 57600
rect 261 56617 917 56669
rect 969 56617 1041 56669
rect 1093 56617 1165 56669
rect 1217 56617 1289 56669
rect 1341 56617 1413 56669
rect 1465 56617 1537 56669
rect 1589 56617 1661 56669
rect 1713 56617 1785 56669
rect 1837 56617 2161 56669
rect 261 56545 2161 56617
rect 261 56493 917 56545
rect 969 56493 1041 56545
rect 1093 56493 1165 56545
rect 1217 56493 1289 56545
rect 1341 56493 1413 56545
rect 1465 56493 1537 56545
rect 1589 56493 1661 56545
rect 1713 56493 1785 56545
rect 1837 56493 2161 56545
rect 261 56421 2161 56493
rect 261 56369 917 56421
rect 969 56369 1041 56421
rect 1093 56369 1165 56421
rect 1217 56369 1289 56421
rect 1341 56369 1413 56421
rect 1465 56369 1537 56421
rect 1589 56369 1661 56421
rect 1713 56369 1785 56421
rect 1837 56369 2161 56421
rect 261 56297 2161 56369
rect 261 56245 917 56297
rect 969 56245 1041 56297
rect 1093 56245 1165 56297
rect 1217 56245 1289 56297
rect 1341 56245 1413 56297
rect 1465 56245 1537 56297
rect 1589 56245 1661 56297
rect 1713 56245 1785 56297
rect 1837 56245 2161 56297
rect 261 56173 2161 56245
rect 261 56121 917 56173
rect 969 56121 1041 56173
rect 1093 56121 1165 56173
rect 1217 56121 1289 56173
rect 1341 56121 1413 56173
rect 1465 56121 1537 56173
rect 1589 56121 1661 56173
rect 1713 56121 1785 56173
rect 1837 56121 2161 56173
rect 261 56049 2161 56121
rect 261 55997 917 56049
rect 969 55997 1041 56049
rect 1093 55997 1165 56049
rect 1217 55997 1289 56049
rect 1341 55997 1413 56049
rect 1465 55997 1537 56049
rect 1589 55997 1661 56049
rect 1713 55997 1785 56049
rect 1837 55997 2161 56049
rect 261 55925 2161 55997
rect 261 55873 917 55925
rect 969 55873 1041 55925
rect 1093 55873 1165 55925
rect 1217 55873 1289 55925
rect 1341 55873 1413 55925
rect 1465 55873 1537 55925
rect 1589 55873 1661 55925
rect 1713 55873 1785 55925
rect 1837 55873 2161 55925
rect 261 55801 2161 55873
rect 261 55749 917 55801
rect 969 55749 1041 55801
rect 1093 55749 1165 55801
rect 1217 55749 1289 55801
rect 1341 55749 1413 55801
rect 1465 55749 1537 55801
rect 1589 55749 1661 55801
rect 1713 55749 1785 55801
rect 1837 55749 2161 55801
rect 261 55748 2161 55749
rect 261 55692 315 55748
rect 371 55692 439 55748
rect 495 55692 563 55748
rect 619 55692 687 55748
rect 743 55692 811 55748
rect 867 55692 935 55748
rect 991 55692 1059 55748
rect 1115 55692 1183 55748
rect 1239 55692 1307 55748
rect 1363 55692 1431 55748
rect 1487 55692 1555 55748
rect 1611 55692 1679 55748
rect 1735 55692 1803 55748
rect 1859 55692 1927 55748
rect 1983 55692 2051 55748
rect 2107 55692 2161 55748
rect 261 55677 2161 55692
rect 261 55625 917 55677
rect 969 55625 1041 55677
rect 1093 55625 1165 55677
rect 1217 55625 1289 55677
rect 1341 55625 1413 55677
rect 1465 55625 1537 55677
rect 1589 55625 1661 55677
rect 1713 55625 1785 55677
rect 1837 55625 2161 55677
rect 261 55624 2161 55625
rect 261 55568 315 55624
rect 371 55568 439 55624
rect 495 55568 563 55624
rect 619 55568 687 55624
rect 743 55568 811 55624
rect 867 55568 935 55624
rect 991 55568 1059 55624
rect 1115 55568 1183 55624
rect 1239 55568 1307 55624
rect 1363 55568 1431 55624
rect 1487 55568 1555 55624
rect 1611 55568 1679 55624
rect 1735 55568 1803 55624
rect 1859 55568 1927 55624
rect 1983 55568 2051 55624
rect 2107 55568 2161 55624
rect 261 55553 2161 55568
rect 261 55501 917 55553
rect 969 55501 1041 55553
rect 1093 55501 1165 55553
rect 1217 55501 1289 55553
rect 1341 55501 1413 55553
rect 1465 55501 1537 55553
rect 1589 55501 1661 55553
rect 1713 55501 1785 55553
rect 1837 55501 2161 55553
rect 261 55500 2161 55501
rect 261 55444 315 55500
rect 371 55444 439 55500
rect 495 55444 563 55500
rect 619 55444 687 55500
rect 743 55444 811 55500
rect 867 55444 935 55500
rect 991 55444 1059 55500
rect 1115 55444 1183 55500
rect 1239 55444 1307 55500
rect 1363 55444 1431 55500
rect 1487 55444 1555 55500
rect 1611 55444 1679 55500
rect 1735 55444 1803 55500
rect 1859 55444 1927 55500
rect 1983 55444 2051 55500
rect 2107 55444 2161 55500
rect 261 55429 2161 55444
rect 261 55377 917 55429
rect 969 55377 1041 55429
rect 1093 55377 1165 55429
rect 1217 55377 1289 55429
rect 1341 55377 1413 55429
rect 1465 55377 1537 55429
rect 1589 55377 1661 55429
rect 1713 55377 1785 55429
rect 1837 55377 2161 55429
rect 261 55376 2161 55377
rect 261 55320 315 55376
rect 371 55320 439 55376
rect 495 55320 563 55376
rect 619 55320 687 55376
rect 743 55320 811 55376
rect 867 55320 935 55376
rect 991 55320 1059 55376
rect 1115 55320 1183 55376
rect 1239 55320 1307 55376
rect 1363 55320 1431 55376
rect 1487 55320 1555 55376
rect 1611 55320 1679 55376
rect 1735 55320 1803 55376
rect 1859 55320 1927 55376
rect 1983 55320 2051 55376
rect 2107 55320 2161 55376
rect 261 55305 2161 55320
rect 261 55253 917 55305
rect 969 55253 1041 55305
rect 1093 55253 1165 55305
rect 1217 55253 1289 55305
rect 1341 55253 1413 55305
rect 1465 55253 1537 55305
rect 1589 55253 1661 55305
rect 1713 55253 1785 55305
rect 1837 55253 2161 55305
rect 261 55252 2161 55253
rect 261 55196 315 55252
rect 371 55196 439 55252
rect 495 55196 563 55252
rect 619 55196 687 55252
rect 743 55196 811 55252
rect 867 55196 935 55252
rect 991 55196 1059 55252
rect 1115 55196 1183 55252
rect 1239 55196 1307 55252
rect 1363 55196 1431 55252
rect 1487 55196 1555 55252
rect 1611 55196 1679 55252
rect 1735 55196 1803 55252
rect 1859 55196 1927 55252
rect 1983 55196 2051 55252
rect 2107 55196 2161 55252
rect 261 55181 2161 55196
rect 261 55129 917 55181
rect 969 55129 1041 55181
rect 1093 55129 1165 55181
rect 1217 55129 1289 55181
rect 1341 55129 1413 55181
rect 1465 55129 1537 55181
rect 1589 55129 1661 55181
rect 1713 55129 1785 55181
rect 1837 55129 2161 55181
rect 261 55128 2161 55129
rect 261 55072 315 55128
rect 371 55072 439 55128
rect 495 55072 563 55128
rect 619 55072 687 55128
rect 743 55072 811 55128
rect 867 55072 935 55128
rect 991 55072 1059 55128
rect 1115 55072 1183 55128
rect 1239 55072 1307 55128
rect 1363 55072 1431 55128
rect 1487 55072 1555 55128
rect 1611 55072 1679 55128
rect 1735 55072 1803 55128
rect 1859 55072 1927 55128
rect 1983 55072 2051 55128
rect 2107 55072 2161 55128
rect 261 55057 2161 55072
rect 261 55005 917 55057
rect 969 55005 1041 55057
rect 1093 55005 1165 55057
rect 1217 55005 1289 55057
rect 1341 55005 1413 55057
rect 1465 55005 1537 55057
rect 1589 55005 1661 55057
rect 1713 55005 1785 55057
rect 1837 55005 2161 55057
rect 261 55004 2161 55005
rect 261 54948 315 55004
rect 371 54948 439 55004
rect 495 54948 563 55004
rect 619 54948 687 55004
rect 743 54948 811 55004
rect 867 54948 935 55004
rect 991 54948 1059 55004
rect 1115 54948 1183 55004
rect 1239 54948 1307 55004
rect 1363 54948 1431 55004
rect 1487 54948 1555 55004
rect 1611 54948 1679 55004
rect 1735 54948 1803 55004
rect 1859 54948 1927 55004
rect 1983 54948 2051 55004
rect 2107 54948 2161 55004
rect 261 54933 2161 54948
rect 261 54881 917 54933
rect 969 54881 1041 54933
rect 1093 54881 1165 54933
rect 1217 54881 1289 54933
rect 1341 54881 1413 54933
rect 1465 54881 1537 54933
rect 1589 54881 1661 54933
rect 1713 54881 1785 54933
rect 1837 54881 2161 54933
rect 261 54880 2161 54881
rect 261 54824 315 54880
rect 371 54824 439 54880
rect 495 54824 563 54880
rect 619 54824 687 54880
rect 743 54824 811 54880
rect 867 54824 935 54880
rect 991 54824 1059 54880
rect 1115 54824 1183 54880
rect 1239 54824 1307 54880
rect 1363 54824 1431 54880
rect 1487 54824 1555 54880
rect 1611 54824 1679 54880
rect 1735 54824 1803 54880
rect 1859 54824 1927 54880
rect 1983 54824 2051 54880
rect 2107 54824 2161 54880
rect 261 54809 2161 54824
rect 261 54757 917 54809
rect 969 54757 1041 54809
rect 1093 54757 1165 54809
rect 1217 54757 1289 54809
rect 1341 54757 1413 54809
rect 1465 54757 1537 54809
rect 1589 54757 1661 54809
rect 1713 54757 1785 54809
rect 1837 54757 2161 54809
rect 261 54756 2161 54757
rect 261 54700 315 54756
rect 371 54700 439 54756
rect 495 54700 563 54756
rect 619 54700 687 54756
rect 743 54700 811 54756
rect 867 54700 935 54756
rect 991 54700 1059 54756
rect 1115 54700 1183 54756
rect 1239 54700 1307 54756
rect 1363 54700 1431 54756
rect 1487 54700 1555 54756
rect 1611 54700 1679 54756
rect 1735 54700 1803 54756
rect 1859 54700 1927 54756
rect 1983 54700 2051 54756
rect 2107 54700 2161 54756
rect 261 54685 2161 54700
rect 261 54633 917 54685
rect 969 54633 1041 54685
rect 1093 54633 1165 54685
rect 1217 54633 1289 54685
rect 1341 54633 1413 54685
rect 1465 54633 1537 54685
rect 1589 54633 1661 54685
rect 1713 54633 1785 54685
rect 1837 54633 2161 54685
rect 261 54632 2161 54633
rect 261 54576 315 54632
rect 371 54576 439 54632
rect 495 54576 563 54632
rect 619 54576 687 54632
rect 743 54576 811 54632
rect 867 54576 935 54632
rect 991 54576 1059 54632
rect 1115 54576 1183 54632
rect 1239 54576 1307 54632
rect 1363 54576 1431 54632
rect 1487 54576 1555 54632
rect 1611 54576 1679 54632
rect 1735 54576 1803 54632
rect 1859 54576 1927 54632
rect 1983 54576 2051 54632
rect 2107 54576 2161 54632
rect 261 54561 2161 54576
rect 261 54509 917 54561
rect 969 54509 1041 54561
rect 1093 54509 1165 54561
rect 1217 54509 1289 54561
rect 1341 54509 1413 54561
rect 1465 54509 1537 54561
rect 1589 54509 1661 54561
rect 1713 54509 1785 54561
rect 1837 54509 2161 54561
rect 261 54508 2161 54509
rect 261 54452 315 54508
rect 371 54452 439 54508
rect 495 54452 563 54508
rect 619 54452 687 54508
rect 743 54452 811 54508
rect 867 54452 935 54508
rect 991 54452 1059 54508
rect 1115 54452 1183 54508
rect 1239 54452 1307 54508
rect 1363 54452 1431 54508
rect 1487 54452 1555 54508
rect 1611 54452 1679 54508
rect 1735 54452 1803 54508
rect 1859 54452 1927 54508
rect 1983 54452 2051 54508
rect 2107 54452 2161 54508
rect 261 54437 2161 54452
rect 261 54385 917 54437
rect 969 54385 1041 54437
rect 1093 54385 1165 54437
rect 1217 54385 1289 54437
rect 1341 54385 1413 54437
rect 1465 54385 1537 54437
rect 1589 54385 1661 54437
rect 1713 54385 1785 54437
rect 1837 54385 2161 54437
rect 261 54313 2161 54385
rect 261 54261 917 54313
rect 969 54261 1041 54313
rect 1093 54261 1165 54313
rect 1217 54261 1289 54313
rect 1341 54261 1413 54313
rect 1465 54261 1537 54313
rect 1589 54261 1661 54313
rect 1713 54261 1785 54313
rect 1837 54261 2161 54313
rect 261 54189 2161 54261
rect 261 54137 917 54189
rect 969 54137 1041 54189
rect 1093 54137 1165 54189
rect 1217 54137 1289 54189
rect 1341 54137 1413 54189
rect 1465 54137 1537 54189
rect 1589 54137 1661 54189
rect 1713 54137 1785 54189
rect 1837 54137 2161 54189
rect 261 54065 2161 54137
rect 261 54013 917 54065
rect 969 54013 1041 54065
rect 1093 54013 1165 54065
rect 1217 54013 1289 54065
rect 1341 54013 1413 54065
rect 1465 54013 1537 54065
rect 1589 54013 1661 54065
rect 1713 54013 1785 54065
rect 1837 54013 2161 54065
rect 261 53941 2161 54013
rect 261 53889 917 53941
rect 969 53889 1041 53941
rect 1093 53889 1165 53941
rect 1217 53889 1289 53941
rect 1341 53889 1413 53941
rect 1465 53889 1537 53941
rect 1589 53889 1661 53941
rect 1713 53889 1785 53941
rect 1837 53889 2161 53941
rect 261 53817 2161 53889
rect 261 53765 917 53817
rect 969 53765 1041 53817
rect 1093 53765 1165 53817
rect 1217 53765 1289 53817
rect 1341 53765 1413 53817
rect 1465 53765 1537 53817
rect 1589 53765 1661 53817
rect 1713 53765 1785 53817
rect 1837 53765 2161 53817
rect 261 53693 2161 53765
rect 261 53641 917 53693
rect 969 53641 1041 53693
rect 1093 53641 1165 53693
rect 1217 53641 1289 53693
rect 1341 53641 1413 53693
rect 1465 53641 1537 53693
rect 1589 53641 1661 53693
rect 1713 53641 1785 53693
rect 1837 53641 2161 53693
rect -11 52576 86 52600
rect -11 51224 20 52576
rect 76 51224 86 52576
rect -11 51200 86 51224
rect 261 50948 2161 53641
rect 2481 57225 2681 57278
rect 2481 57169 2491 57225
rect 2547 57169 2615 57225
rect 2671 57169 2681 57225
rect 2481 57108 2681 57169
rect 2481 57101 2501 57108
rect 2481 57045 2491 57101
rect 2553 57056 2609 57108
rect 2661 57101 2681 57108
rect 2547 57045 2615 57056
rect 2671 57045 2681 57101
rect 2481 56977 2681 57045
rect 2481 56921 2491 56977
rect 2547 56921 2615 56977
rect 2671 56921 2681 56977
rect 2481 56853 2681 56921
rect 2481 56797 2491 56853
rect 2547 56797 2615 56853
rect 2671 56797 2681 56853
rect 2481 56729 2681 56797
rect 2481 56673 2491 56729
rect 2547 56673 2615 56729
rect 2671 56673 2681 56729
rect 2481 56605 2681 56673
rect 2481 56549 2491 56605
rect 2547 56549 2615 56605
rect 2671 56549 2681 56605
rect 2481 56481 2681 56549
rect 2481 56425 2491 56481
rect 2547 56425 2615 56481
rect 2671 56425 2681 56481
rect 2481 56357 2681 56425
rect 2481 56301 2491 56357
rect 2547 56301 2615 56357
rect 2671 56301 2681 56357
rect 2481 56233 2681 56301
rect 2481 56177 2491 56233
rect 2547 56177 2615 56233
rect 2671 56177 2681 56233
rect 2481 56109 2681 56177
rect 2481 56053 2491 56109
rect 2547 56053 2615 56109
rect 2671 56053 2681 56109
rect 2481 54148 2681 56053
rect 2481 54092 2491 54148
rect 2547 54092 2615 54148
rect 2671 54092 2681 54148
rect 2481 54024 2681 54092
rect 2481 53968 2491 54024
rect 2547 53968 2615 54024
rect 2671 53968 2681 54024
rect 2481 53900 2681 53968
rect 2481 53844 2491 53900
rect 2547 53844 2615 53900
rect 2671 53844 2681 53900
rect 2481 53776 2681 53844
rect 2481 53720 2491 53776
rect 2547 53720 2615 53776
rect 2671 53720 2681 53776
rect 2481 53652 2681 53720
rect 2481 53596 2491 53652
rect 2547 53596 2615 53652
rect 2671 53596 2681 53652
rect 2481 53528 2681 53596
rect 2481 53472 2491 53528
rect 2547 53484 2615 53528
rect 2481 53432 2501 53472
rect 2553 53432 2609 53484
rect 2671 53472 2681 53528
rect 2661 53432 2681 53472
rect 2481 53404 2681 53432
rect 2481 53348 2491 53404
rect 2547 53376 2615 53404
rect 2481 53324 2501 53348
rect 2553 53324 2609 53376
rect 2671 53348 2681 53404
rect 2661 53324 2681 53348
rect 2481 53280 2681 53324
rect 2481 53224 2491 53280
rect 2547 53268 2615 53280
rect 2481 53216 2501 53224
rect 2553 53216 2609 53268
rect 2671 53224 2681 53280
rect 2661 53216 2681 53224
rect 2481 53156 2681 53216
rect 2481 53100 2491 53156
rect 2547 53100 2615 53156
rect 2671 53100 2681 53156
rect 2481 53032 2681 53100
rect 2481 52976 2491 53032
rect 2547 52976 2615 53032
rect 2671 52976 2681 53032
rect 2481 52908 2681 52976
rect 2481 52852 2491 52908
rect 2547 52852 2615 52908
rect 2671 52852 2681 52908
rect 261 50892 315 50948
rect 371 50892 439 50948
rect 495 50892 563 50948
rect 619 50892 687 50948
rect 743 50892 811 50948
rect 867 50892 935 50948
rect 991 50892 1059 50948
rect 1115 50892 1183 50948
rect 1239 50892 1307 50948
rect 1363 50892 1431 50948
rect 1487 50892 1555 50948
rect 1611 50892 1679 50948
rect 1735 50892 1803 50948
rect 1859 50892 1927 50948
rect 1983 50892 2051 50948
rect 2107 50892 2161 50948
rect 261 50824 2161 50892
rect 261 50768 315 50824
rect 371 50768 439 50824
rect 495 50768 563 50824
rect 619 50768 687 50824
rect 743 50768 811 50824
rect 867 50768 935 50824
rect 991 50768 1059 50824
rect 1115 50768 1183 50824
rect 1239 50768 1307 50824
rect 1363 50768 1431 50824
rect 1487 50768 1555 50824
rect 1611 50768 1679 50824
rect 1735 50768 1803 50824
rect 1859 50768 1927 50824
rect 1983 50768 2051 50824
rect 2107 50768 2161 50824
rect 261 50700 2161 50768
rect 261 50644 315 50700
rect 371 50644 439 50700
rect 495 50644 563 50700
rect 619 50644 687 50700
rect 743 50644 811 50700
rect 867 50644 935 50700
rect 991 50644 1059 50700
rect 1115 50644 1183 50700
rect 1239 50644 1307 50700
rect 1363 50644 1431 50700
rect 1487 50644 1555 50700
rect 1611 50644 1679 50700
rect 1735 50644 1803 50700
rect 1859 50644 1927 50700
rect 1983 50644 2051 50700
rect 2107 50644 2161 50700
rect 261 50576 2161 50644
rect 261 50520 315 50576
rect 371 50520 439 50576
rect 495 50520 563 50576
rect 619 50520 687 50576
rect 743 50520 811 50576
rect 867 50520 935 50576
rect 991 50520 1059 50576
rect 1115 50520 1183 50576
rect 1239 50520 1307 50576
rect 1363 50520 1431 50576
rect 1487 50520 1555 50576
rect 1611 50520 1679 50576
rect 1735 50520 1803 50576
rect 1859 50520 1927 50576
rect 1983 50520 2051 50576
rect 2107 50520 2161 50576
rect 261 50452 2161 50520
rect 261 50396 315 50452
rect 371 50396 439 50452
rect 495 50396 563 50452
rect 619 50396 687 50452
rect 743 50396 811 50452
rect 867 50396 935 50452
rect 991 50396 1059 50452
rect 1115 50396 1183 50452
rect 1239 50396 1307 50452
rect 1363 50396 1431 50452
rect 1487 50396 1555 50452
rect 1611 50396 1679 50452
rect 1735 50396 1803 50452
rect 1859 50396 1927 50452
rect 1983 50396 2051 50452
rect 2107 50396 2161 50452
rect 261 50328 2161 50396
rect 261 50272 315 50328
rect 371 50272 439 50328
rect 495 50272 563 50328
rect 619 50272 687 50328
rect 743 50272 811 50328
rect 867 50272 935 50328
rect 991 50272 1059 50328
rect 1115 50272 1183 50328
rect 1239 50272 1307 50328
rect 1363 50272 1431 50328
rect 1487 50272 1555 50328
rect 1611 50272 1679 50328
rect 1735 50272 1803 50328
rect 1859 50272 1927 50328
rect 1983 50272 2051 50328
rect 2107 50272 2161 50328
rect 261 50204 2161 50272
rect 261 50148 315 50204
rect 371 50148 439 50204
rect 495 50148 563 50204
rect 619 50148 687 50204
rect 743 50148 811 50204
rect 867 50148 935 50204
rect 991 50148 1059 50204
rect 1115 50148 1183 50204
rect 1239 50148 1307 50204
rect 1363 50148 1431 50204
rect 1487 50148 1555 50204
rect 1611 50148 1679 50204
rect 1735 50148 1803 50204
rect 1859 50148 1927 50204
rect 1983 50148 2051 50204
rect 2107 50148 2161 50204
rect 261 50080 2161 50148
rect 261 50024 315 50080
rect 371 50024 439 50080
rect 495 50024 563 50080
rect 619 50024 687 50080
rect 743 50024 811 50080
rect 867 50024 935 50080
rect 991 50024 1059 50080
rect 1115 50024 1183 50080
rect 1239 50024 1307 50080
rect 1363 50024 1431 50080
rect 1487 50024 1555 50080
rect 1611 50024 1679 50080
rect 1735 50024 1803 50080
rect 1859 50024 1927 50080
rect 1983 50024 2051 50080
rect 2107 50024 2161 50080
rect 261 49956 2161 50024
rect 261 49900 315 49956
rect 371 49900 439 49956
rect 495 49900 563 49956
rect 619 49900 687 49956
rect 743 49900 811 49956
rect 867 49900 935 49956
rect 991 49900 1059 49956
rect 1115 49900 1183 49956
rect 1239 49900 1307 49956
rect 1363 49900 1431 49956
rect 1487 49900 1555 49956
rect 1611 49900 1679 49956
rect 1735 49900 1803 49956
rect 1859 49900 1927 49956
rect 1983 49900 2051 49956
rect 2107 49900 2161 49956
rect 261 49832 2161 49900
rect 261 49776 315 49832
rect 371 49776 439 49832
rect 495 49776 563 49832
rect 619 49776 687 49832
rect 743 49776 811 49832
rect 867 49776 935 49832
rect 991 49776 1059 49832
rect 1115 49776 1183 49832
rect 1239 49776 1307 49832
rect 1363 49776 1431 49832
rect 1487 49776 1555 49832
rect 1611 49776 1679 49832
rect 1735 49776 1803 49832
rect 1859 49776 1927 49832
rect 1983 49776 2051 49832
rect 2107 49776 2161 49832
rect 261 49708 2161 49776
rect 261 49652 315 49708
rect 371 49652 439 49708
rect 495 49652 563 49708
rect 619 49652 687 49708
rect 743 49652 811 49708
rect 867 49652 935 49708
rect 991 49652 1059 49708
rect 1115 49652 1183 49708
rect 1239 49652 1307 49708
rect 1363 49652 1431 49708
rect 1487 49652 1555 49708
rect 1611 49652 1679 49708
rect 1735 49652 1803 49708
rect 1859 49652 1927 49708
rect 1983 49652 2051 49708
rect 2107 49652 2161 49708
rect 261 47748 2161 49652
rect 261 47692 315 47748
rect 371 47692 439 47748
rect 495 47692 563 47748
rect 619 47692 687 47748
rect 743 47692 811 47748
rect 867 47692 935 47748
rect 991 47692 1059 47748
rect 1115 47692 1183 47748
rect 1239 47692 1307 47748
rect 1363 47692 1431 47748
rect 1487 47692 1555 47748
rect 1611 47692 1679 47748
rect 1735 47692 1803 47748
rect 1859 47692 1927 47748
rect 1983 47692 2051 47748
rect 2107 47692 2161 47748
rect 261 47624 2161 47692
rect 261 47568 315 47624
rect 371 47568 439 47624
rect 495 47568 563 47624
rect 619 47568 687 47624
rect 743 47568 811 47624
rect 867 47568 935 47624
rect 991 47568 1059 47624
rect 1115 47568 1183 47624
rect 1239 47568 1307 47624
rect 1363 47568 1431 47624
rect 1487 47568 1555 47624
rect 1611 47568 1679 47624
rect 1735 47568 1803 47624
rect 1859 47568 1927 47624
rect 1983 47568 2051 47624
rect 2107 47568 2161 47624
rect 261 47500 2161 47568
rect 261 47444 315 47500
rect 371 47444 439 47500
rect 495 47444 563 47500
rect 619 47444 687 47500
rect 743 47444 811 47500
rect 867 47444 935 47500
rect 991 47444 1059 47500
rect 1115 47444 1183 47500
rect 1239 47444 1307 47500
rect 1363 47444 1431 47500
rect 1487 47444 1555 47500
rect 1611 47444 1679 47500
rect 1735 47444 1803 47500
rect 1859 47444 1927 47500
rect 1983 47444 2051 47500
rect 2107 47444 2161 47500
rect 261 47376 2161 47444
rect 261 47320 315 47376
rect 371 47320 439 47376
rect 495 47320 563 47376
rect 619 47320 687 47376
rect 743 47320 811 47376
rect 867 47320 935 47376
rect 991 47320 1059 47376
rect 1115 47320 1183 47376
rect 1239 47320 1307 47376
rect 1363 47320 1431 47376
rect 1487 47320 1555 47376
rect 1611 47320 1679 47376
rect 1735 47320 1803 47376
rect 1859 47320 1927 47376
rect 1983 47320 2051 47376
rect 2107 47320 2161 47376
rect 261 47281 2161 47320
rect 2279 52521 2355 52600
rect 2279 52465 2289 52521
rect 2345 52465 2355 52521
rect 2279 52389 2355 52465
rect 2279 52333 2289 52389
rect 2345 52333 2355 52389
rect 2279 52257 2355 52333
rect 2279 52201 2289 52257
rect 2345 52201 2355 52257
rect 2279 52125 2355 52201
rect 2279 52069 2289 52125
rect 2345 52069 2355 52125
rect 2279 51993 2355 52069
rect 2279 51937 2289 51993
rect 2345 51937 2355 51993
rect 2279 51861 2355 51937
rect 2279 51805 2289 51861
rect 2345 51805 2355 51861
rect 2279 51729 2355 51805
rect 2279 51673 2289 51729
rect 2345 51673 2355 51729
rect 2279 51597 2355 51673
rect 2279 51541 2289 51597
rect 2345 51541 2355 51597
rect 2279 51465 2355 51541
rect 2279 51409 2289 51465
rect 2345 51409 2355 51465
rect 2279 51333 2355 51409
rect 2279 51277 2289 51333
rect 2345 51277 2355 51333
rect 305 47252 2117 47281
rect 305 47196 315 47252
rect 371 47196 439 47252
rect 495 47196 563 47252
rect 619 47196 687 47252
rect 743 47196 811 47252
rect 867 47196 935 47252
rect 991 47196 1059 47252
rect 1115 47196 1183 47252
rect 1239 47196 1307 47252
rect 1363 47196 1431 47252
rect 1487 47196 1555 47252
rect 1611 47196 1679 47252
rect 1735 47196 1803 47252
rect 1859 47196 1927 47252
rect 1983 47196 2051 47252
rect 2107 47196 2117 47252
rect 305 47128 2117 47196
rect 305 47072 315 47128
rect 371 47072 439 47128
rect 495 47072 563 47128
rect 619 47072 687 47128
rect 743 47072 811 47128
rect 867 47072 935 47128
rect 991 47072 1059 47128
rect 1115 47072 1183 47128
rect 1239 47072 1307 47128
rect 1363 47072 1431 47128
rect 1487 47072 1555 47128
rect 1611 47072 1679 47128
rect 1735 47072 1803 47128
rect 1859 47072 1927 47128
rect 1983 47072 2051 47128
rect 2107 47072 2117 47128
rect 305 47004 2117 47072
rect 305 46948 315 47004
rect 371 46948 439 47004
rect 495 46948 563 47004
rect 619 46948 687 47004
rect 743 46948 811 47004
rect 867 46948 935 47004
rect 991 46948 1059 47004
rect 1115 46948 1183 47004
rect 1239 46948 1307 47004
rect 1363 46948 1431 47004
rect 1487 46948 1555 47004
rect 1611 46948 1679 47004
rect 1735 46948 1803 47004
rect 1859 46948 1927 47004
rect 1983 46948 2051 47004
rect 2107 46948 2117 47004
rect 305 46880 2117 46948
rect 305 46824 315 46880
rect 371 46824 439 46880
rect 495 46824 563 46880
rect 619 46824 687 46880
rect 743 46824 811 46880
rect 867 46824 935 46880
rect 991 46824 1059 46880
rect 1115 46824 1183 46880
rect 1239 46824 1307 46880
rect 1363 46824 1431 46880
rect 1487 46824 1555 46880
rect 1611 46824 1679 46880
rect 1735 46824 1803 46880
rect 1859 46824 1927 46880
rect 1983 46824 2051 46880
rect 2107 46824 2117 46880
rect 305 46756 2117 46824
rect 305 46700 315 46756
rect 371 46700 439 46756
rect 495 46700 563 46756
rect 619 46700 687 46756
rect 743 46700 811 46756
rect 867 46700 935 46756
rect 991 46700 1059 46756
rect 1115 46700 1183 46756
rect 1239 46700 1307 46756
rect 1363 46700 1431 46756
rect 1487 46700 1555 46756
rect 1611 46700 1679 46756
rect 1735 46700 1803 46756
rect 1859 46700 1927 46756
rect 1983 46700 2051 46756
rect 2107 46700 2117 46756
rect 305 46632 2117 46700
rect 305 46576 315 46632
rect 371 46576 439 46632
rect 495 46576 563 46632
rect 619 46576 687 46632
rect 743 46576 811 46632
rect 867 46576 935 46632
rect 991 46576 1059 46632
rect 1115 46576 1183 46632
rect 1239 46576 1307 46632
rect 1363 46576 1431 46632
rect 1487 46576 1555 46632
rect 1611 46576 1679 46632
rect 1735 46576 1803 46632
rect 1859 46576 1927 46632
rect 1983 46576 2051 46632
rect 2107 46576 2117 46632
rect 305 46508 2117 46576
rect 305 46452 315 46508
rect 371 46452 439 46508
rect 495 46452 563 46508
rect 619 46452 687 46508
rect 743 46452 811 46508
rect 867 46452 935 46508
rect 991 46452 1059 46508
rect 1115 46452 1183 46508
rect 1239 46452 1307 46508
rect 1363 46452 1431 46508
rect 1487 46452 1555 46508
rect 1611 46452 1679 46508
rect 1735 46452 1803 46508
rect 1859 46452 1927 46508
rect 1983 46452 2051 46508
rect 2107 46452 2117 46508
rect 305 46442 2117 46452
rect 305 44548 2117 44558
rect 305 44492 315 44548
rect 371 44492 439 44548
rect 495 44492 563 44548
rect 619 44492 687 44548
rect 743 44492 811 44548
rect 867 44492 935 44548
rect 991 44492 1059 44548
rect 1115 44492 1183 44548
rect 1239 44492 1307 44548
rect 1363 44492 1431 44548
rect 1487 44492 1555 44548
rect 1611 44492 1679 44548
rect 1735 44492 1803 44548
rect 1859 44492 1927 44548
rect 1983 44492 2051 44548
rect 2107 44492 2117 44548
rect 305 44424 2117 44492
rect 305 44368 315 44424
rect 371 44368 439 44424
rect 495 44368 563 44424
rect 619 44368 687 44424
rect 743 44368 811 44424
rect 867 44368 935 44424
rect 991 44368 1059 44424
rect 1115 44368 1183 44424
rect 1239 44368 1307 44424
rect 1363 44368 1431 44424
rect 1487 44368 1555 44424
rect 1611 44368 1679 44424
rect 1735 44368 1803 44424
rect 1859 44368 1927 44424
rect 1983 44368 2051 44424
rect 2107 44368 2117 44424
rect 305 44300 2117 44368
rect 305 44244 315 44300
rect 371 44244 439 44300
rect 495 44244 563 44300
rect 619 44244 687 44300
rect 743 44244 811 44300
rect 867 44244 935 44300
rect 991 44244 1059 44300
rect 1115 44244 1183 44300
rect 1239 44244 1307 44300
rect 1363 44244 1431 44300
rect 1487 44244 1555 44300
rect 1611 44244 1679 44300
rect 1735 44244 1803 44300
rect 1859 44244 1927 44300
rect 1983 44244 2051 44300
rect 2107 44244 2117 44300
rect 305 44176 2117 44244
rect 305 44120 315 44176
rect 371 44120 439 44176
rect 495 44120 563 44176
rect 619 44120 687 44176
rect 743 44120 811 44176
rect 867 44120 935 44176
rect 991 44120 1059 44176
rect 1115 44120 1183 44176
rect 1239 44120 1307 44176
rect 1363 44120 1431 44176
rect 1487 44120 1555 44176
rect 1611 44120 1679 44176
rect 1735 44120 1803 44176
rect 1859 44120 1927 44176
rect 1983 44120 2051 44176
rect 2107 44120 2117 44176
rect 305 44052 2117 44120
rect 305 43996 315 44052
rect 371 43996 439 44052
rect 495 43996 563 44052
rect 619 43996 687 44052
rect 743 43996 811 44052
rect 867 43996 935 44052
rect 991 43996 1059 44052
rect 1115 43996 1183 44052
rect 1239 43996 1307 44052
rect 1363 43996 1431 44052
rect 1487 43996 1555 44052
rect 1611 43996 1679 44052
rect 1735 43996 1803 44052
rect 1859 43996 1927 44052
rect 1983 43996 2051 44052
rect 2107 43996 2117 44052
rect 305 43928 2117 43996
rect 305 43872 315 43928
rect 371 43872 439 43928
rect 495 43872 563 43928
rect 619 43872 687 43928
rect 743 43872 811 43928
rect 867 43872 935 43928
rect 991 43872 1059 43928
rect 1115 43872 1183 43928
rect 1239 43872 1307 43928
rect 1363 43872 1431 43928
rect 1487 43872 1555 43928
rect 1611 43872 1679 43928
rect 1735 43872 1803 43928
rect 1859 43872 1927 43928
rect 1983 43872 2051 43928
rect 2107 43872 2117 43928
rect 305 43804 2117 43872
rect 305 43748 315 43804
rect 371 43748 439 43804
rect 495 43748 563 43804
rect 619 43748 687 43804
rect 743 43748 811 43804
rect 867 43748 935 43804
rect 991 43748 1059 43804
rect 1115 43748 1183 43804
rect 1239 43748 1307 43804
rect 1363 43748 1431 43804
rect 1487 43748 1555 43804
rect 1611 43748 1679 43804
rect 1735 43748 1803 43804
rect 1859 43748 1927 43804
rect 1983 43748 2051 43804
rect 2107 43748 2117 43804
rect 305 43680 2117 43748
rect 305 43624 315 43680
rect 371 43624 439 43680
rect 495 43624 563 43680
rect 619 43624 687 43680
rect 743 43624 811 43680
rect 867 43624 935 43680
rect 991 43624 1059 43680
rect 1115 43624 1183 43680
rect 1239 43624 1307 43680
rect 1363 43624 1431 43680
rect 1487 43624 1555 43680
rect 1611 43624 1679 43680
rect 1735 43624 1803 43680
rect 1859 43624 1927 43680
rect 1983 43624 2051 43680
rect 2107 43624 2117 43680
rect 305 43556 2117 43624
rect 305 43500 315 43556
rect 371 43500 439 43556
rect 495 43500 563 43556
rect 619 43500 687 43556
rect 743 43500 811 43556
rect 867 43500 935 43556
rect 991 43500 1059 43556
rect 1115 43500 1183 43556
rect 1239 43500 1307 43556
rect 1363 43500 1431 43556
rect 1487 43500 1555 43556
rect 1611 43500 1679 43556
rect 1735 43500 1803 43556
rect 1859 43500 1927 43556
rect 1983 43500 2051 43556
rect 2107 43500 2117 43556
rect 305 43432 2117 43500
rect 305 43376 315 43432
rect 371 43376 439 43432
rect 495 43376 563 43432
rect 619 43376 687 43432
rect 743 43376 811 43432
rect 867 43376 935 43432
rect 991 43376 1059 43432
rect 1115 43376 1183 43432
rect 1239 43376 1307 43432
rect 1363 43376 1431 43432
rect 1487 43376 1555 43432
rect 1611 43376 1679 43432
rect 1735 43376 1803 43432
rect 1859 43376 1927 43432
rect 1983 43376 2051 43432
rect 2107 43376 2117 43432
rect 305 43308 2117 43376
rect 305 43252 315 43308
rect 371 43252 439 43308
rect 495 43252 563 43308
rect 619 43252 687 43308
rect 743 43252 811 43308
rect 867 43252 935 43308
rect 991 43252 1059 43308
rect 1115 43252 1183 43308
rect 1239 43252 1307 43308
rect 1363 43252 1431 43308
rect 1487 43252 1555 43308
rect 1611 43252 1679 43308
rect 1735 43252 1803 43308
rect 1859 43252 1927 43308
rect 1983 43252 2051 43308
rect 2107 43252 2117 43308
rect 305 43242 2117 43252
rect 305 42948 2117 42958
rect 305 42892 315 42948
rect 371 42892 439 42948
rect 495 42892 563 42948
rect 619 42892 687 42948
rect 743 42892 811 42948
rect 867 42892 935 42948
rect 991 42892 1059 42948
rect 1115 42892 1183 42948
rect 1239 42892 1307 42948
rect 1363 42892 1431 42948
rect 1487 42892 1555 42948
rect 1611 42892 1679 42948
rect 1735 42892 1803 42948
rect 1859 42892 1927 42948
rect 1983 42892 2051 42948
rect 2107 42892 2117 42948
rect 305 42824 2117 42892
rect 305 42768 315 42824
rect 371 42768 439 42824
rect 495 42768 563 42824
rect 619 42768 687 42824
rect 743 42768 811 42824
rect 867 42768 935 42824
rect 991 42768 1059 42824
rect 1115 42768 1183 42824
rect 1239 42768 1307 42824
rect 1363 42768 1431 42824
rect 1487 42768 1555 42824
rect 1611 42768 1679 42824
rect 1735 42768 1803 42824
rect 1859 42768 1927 42824
rect 1983 42768 2051 42824
rect 2107 42768 2117 42824
rect 305 42700 2117 42768
rect 305 42644 315 42700
rect 371 42644 439 42700
rect 495 42644 563 42700
rect 619 42644 687 42700
rect 743 42644 811 42700
rect 867 42644 935 42700
rect 991 42644 1059 42700
rect 1115 42644 1183 42700
rect 1239 42644 1307 42700
rect 1363 42644 1431 42700
rect 1487 42644 1555 42700
rect 1611 42644 1679 42700
rect 1735 42644 1803 42700
rect 1859 42644 1927 42700
rect 1983 42644 2051 42700
rect 2107 42644 2117 42700
rect 305 42576 2117 42644
rect 305 42520 315 42576
rect 371 42520 439 42576
rect 495 42520 563 42576
rect 619 42520 687 42576
rect 743 42520 811 42576
rect 867 42520 935 42576
rect 991 42520 1059 42576
rect 1115 42520 1183 42576
rect 1239 42520 1307 42576
rect 1363 42520 1431 42576
rect 1487 42520 1555 42576
rect 1611 42520 1679 42576
rect 1735 42520 1803 42576
rect 1859 42520 1927 42576
rect 1983 42520 2051 42576
rect 2107 42520 2117 42576
rect 305 42452 2117 42520
rect 305 42396 315 42452
rect 371 42396 439 42452
rect 495 42396 563 42452
rect 619 42396 687 42452
rect 743 42396 811 42452
rect 867 42396 935 42452
rect 991 42396 1059 42452
rect 1115 42396 1183 42452
rect 1239 42396 1307 42452
rect 1363 42396 1431 42452
rect 1487 42396 1555 42452
rect 1611 42396 1679 42452
rect 1735 42396 1803 42452
rect 1859 42396 1927 42452
rect 1983 42396 2051 42452
rect 2107 42396 2117 42452
rect 305 42328 2117 42396
rect 305 42272 315 42328
rect 371 42272 439 42328
rect 495 42272 563 42328
rect 619 42272 687 42328
rect 743 42272 811 42328
rect 867 42272 935 42328
rect 991 42272 1059 42328
rect 1115 42272 1183 42328
rect 1239 42272 1307 42328
rect 1363 42272 1431 42328
rect 1487 42272 1555 42328
rect 1611 42272 1679 42328
rect 1735 42272 1803 42328
rect 1859 42272 1927 42328
rect 1983 42272 2051 42328
rect 2107 42272 2117 42328
rect 305 42204 2117 42272
rect 305 42148 315 42204
rect 371 42148 439 42204
rect 495 42148 563 42204
rect 619 42148 687 42204
rect 743 42148 811 42204
rect 867 42148 935 42204
rect 991 42148 1059 42204
rect 1115 42148 1183 42204
rect 1239 42148 1307 42204
rect 1363 42148 1431 42204
rect 1487 42148 1555 42204
rect 1611 42148 1679 42204
rect 1735 42148 1803 42204
rect 1859 42148 1927 42204
rect 1983 42148 2051 42204
rect 2107 42148 2117 42204
rect 305 42080 2117 42148
rect 305 42024 315 42080
rect 371 42024 439 42080
rect 495 42024 563 42080
rect 619 42024 687 42080
rect 743 42024 811 42080
rect 867 42024 935 42080
rect 991 42024 1059 42080
rect 1115 42024 1183 42080
rect 1239 42024 1307 42080
rect 1363 42024 1431 42080
rect 1487 42024 1555 42080
rect 1611 42024 1679 42080
rect 1735 42024 1803 42080
rect 1859 42024 1927 42080
rect 1983 42024 2051 42080
rect 2107 42024 2117 42080
rect 305 41956 2117 42024
rect 305 41900 315 41956
rect 371 41900 439 41956
rect 495 41900 563 41956
rect 619 41900 687 41956
rect 743 41900 811 41956
rect 867 41900 935 41956
rect 991 41900 1059 41956
rect 1115 41900 1183 41956
rect 1239 41900 1307 41956
rect 1363 41900 1431 41956
rect 1487 41900 1555 41956
rect 1611 41900 1679 41956
rect 1735 41900 1803 41956
rect 1859 41900 1927 41956
rect 1983 41900 2051 41956
rect 2107 41900 2117 41956
rect 305 41832 2117 41900
rect 305 41776 315 41832
rect 371 41776 439 41832
rect 495 41776 563 41832
rect 619 41776 687 41832
rect 743 41776 811 41832
rect 867 41776 935 41832
rect 991 41776 1059 41832
rect 1115 41776 1183 41832
rect 1239 41776 1307 41832
rect 1363 41776 1431 41832
rect 1487 41776 1555 41832
rect 1611 41776 1679 41832
rect 1735 41776 1803 41832
rect 1859 41776 1927 41832
rect 1983 41776 2051 41832
rect 2107 41776 2117 41832
rect 305 41708 2117 41776
rect 305 41652 315 41708
rect 371 41652 439 41708
rect 495 41652 563 41708
rect 619 41652 687 41708
rect 743 41652 811 41708
rect 867 41652 935 41708
rect 991 41652 1059 41708
rect 1115 41652 1183 41708
rect 1239 41652 1307 41708
rect 1363 41652 1431 41708
rect 1487 41652 1555 41708
rect 1611 41652 1679 41708
rect 1735 41652 1803 41708
rect 1859 41652 1927 41708
rect 1983 41652 2051 41708
rect 2107 41652 2117 41708
rect 305 41642 2117 41652
rect 305 41348 2117 41358
rect 305 41292 315 41348
rect 371 41292 439 41348
rect 495 41292 563 41348
rect 619 41292 687 41348
rect 743 41292 811 41348
rect 867 41292 935 41348
rect 991 41292 1059 41348
rect 1115 41292 1183 41348
rect 1239 41292 1307 41348
rect 1363 41292 1431 41348
rect 1487 41292 1555 41348
rect 1611 41292 1679 41348
rect 1735 41292 1803 41348
rect 1859 41292 1927 41348
rect 1983 41292 2051 41348
rect 2107 41292 2117 41348
rect 305 41224 2117 41292
rect 305 41168 315 41224
rect 371 41168 439 41224
rect 495 41168 563 41224
rect 619 41168 687 41224
rect 743 41168 811 41224
rect 867 41168 935 41224
rect 991 41168 1059 41224
rect 1115 41168 1183 41224
rect 1239 41168 1307 41224
rect 1363 41168 1431 41224
rect 1487 41168 1555 41224
rect 1611 41168 1679 41224
rect 1735 41168 1803 41224
rect 1859 41168 1927 41224
rect 1983 41168 2051 41224
rect 2107 41168 2117 41224
rect 305 41100 2117 41168
rect 305 41044 315 41100
rect 371 41044 439 41100
rect 495 41044 563 41100
rect 619 41044 687 41100
rect 743 41044 811 41100
rect 867 41044 935 41100
rect 991 41044 1059 41100
rect 1115 41044 1183 41100
rect 1239 41044 1307 41100
rect 1363 41044 1431 41100
rect 1487 41044 1555 41100
rect 1611 41044 1679 41100
rect 1735 41044 1803 41100
rect 1859 41044 1927 41100
rect 1983 41044 2051 41100
rect 2107 41044 2117 41100
rect 305 40976 2117 41044
rect 305 40920 315 40976
rect 371 40920 439 40976
rect 495 40920 563 40976
rect 619 40920 687 40976
rect 743 40920 811 40976
rect 867 40920 935 40976
rect 991 40920 1059 40976
rect 1115 40920 1183 40976
rect 1239 40920 1307 40976
rect 1363 40920 1431 40976
rect 1487 40920 1555 40976
rect 1611 40920 1679 40976
rect 1735 40920 1803 40976
rect 1859 40920 1927 40976
rect 1983 40920 2051 40976
rect 2107 40920 2117 40976
rect 305 40852 2117 40920
rect 305 40796 315 40852
rect 371 40796 439 40852
rect 495 40796 563 40852
rect 619 40796 687 40852
rect 743 40796 811 40852
rect 867 40796 935 40852
rect 991 40796 1059 40852
rect 1115 40796 1183 40852
rect 1239 40796 1307 40852
rect 1363 40796 1431 40852
rect 1487 40796 1555 40852
rect 1611 40796 1679 40852
rect 1735 40796 1803 40852
rect 1859 40796 1927 40852
rect 1983 40796 2051 40852
rect 2107 40796 2117 40852
rect 305 40728 2117 40796
rect 305 40672 315 40728
rect 371 40672 439 40728
rect 495 40672 563 40728
rect 619 40672 687 40728
rect 743 40672 811 40728
rect 867 40672 935 40728
rect 991 40672 1059 40728
rect 1115 40672 1183 40728
rect 1239 40672 1307 40728
rect 1363 40672 1431 40728
rect 1487 40672 1555 40728
rect 1611 40672 1679 40728
rect 1735 40672 1803 40728
rect 1859 40672 1927 40728
rect 1983 40672 2051 40728
rect 2107 40672 2117 40728
rect 305 40604 2117 40672
rect 305 40548 315 40604
rect 371 40548 439 40604
rect 495 40548 563 40604
rect 619 40548 687 40604
rect 743 40548 811 40604
rect 867 40548 935 40604
rect 991 40548 1059 40604
rect 1115 40548 1183 40604
rect 1239 40548 1307 40604
rect 1363 40548 1431 40604
rect 1487 40548 1555 40604
rect 1611 40548 1679 40604
rect 1735 40548 1803 40604
rect 1859 40548 1927 40604
rect 1983 40548 2051 40604
rect 2107 40548 2117 40604
rect 305 40480 2117 40548
rect 305 40424 315 40480
rect 371 40424 439 40480
rect 495 40424 563 40480
rect 619 40424 687 40480
rect 743 40424 811 40480
rect 867 40424 935 40480
rect 991 40424 1059 40480
rect 1115 40424 1183 40480
rect 1239 40424 1307 40480
rect 1363 40424 1431 40480
rect 1487 40424 1555 40480
rect 1611 40424 1679 40480
rect 1735 40424 1803 40480
rect 1859 40424 1927 40480
rect 1983 40424 2051 40480
rect 2107 40424 2117 40480
rect 305 40356 2117 40424
rect 305 40300 315 40356
rect 371 40300 439 40356
rect 495 40300 563 40356
rect 619 40300 687 40356
rect 743 40300 811 40356
rect 867 40300 935 40356
rect 991 40300 1059 40356
rect 1115 40300 1183 40356
rect 1239 40300 1307 40356
rect 1363 40300 1431 40356
rect 1487 40300 1555 40356
rect 1611 40300 1679 40356
rect 1735 40300 1803 40356
rect 1859 40300 1927 40356
rect 1983 40300 2051 40356
rect 2107 40300 2117 40356
rect 305 40232 2117 40300
rect 305 40176 315 40232
rect 371 40176 439 40232
rect 495 40176 563 40232
rect 619 40176 687 40232
rect 743 40176 811 40232
rect 867 40176 935 40232
rect 991 40176 1059 40232
rect 1115 40176 1183 40232
rect 1239 40176 1307 40232
rect 1363 40176 1431 40232
rect 1487 40176 1555 40232
rect 1611 40176 1679 40232
rect 1735 40176 1803 40232
rect 1859 40176 1927 40232
rect 1983 40176 2051 40232
rect 2107 40176 2117 40232
rect 305 40108 2117 40176
rect 305 40052 315 40108
rect 371 40052 439 40108
rect 495 40052 563 40108
rect 619 40052 687 40108
rect 743 40052 811 40108
rect 867 40052 935 40108
rect 991 40052 1059 40108
rect 1115 40052 1183 40108
rect 1239 40052 1307 40108
rect 1363 40052 1431 40108
rect 1487 40052 1555 40108
rect 1611 40052 1679 40108
rect 1735 40052 1803 40108
rect 1859 40052 1927 40108
rect 1983 40052 2051 40108
rect 2107 40052 2117 40108
rect 305 40042 2117 40052
rect 305 39748 2117 39758
rect 305 39692 315 39748
rect 371 39692 439 39748
rect 495 39692 563 39748
rect 619 39692 687 39748
rect 743 39692 811 39748
rect 867 39692 935 39748
rect 991 39692 1059 39748
rect 1115 39692 1183 39748
rect 1239 39692 1307 39748
rect 1363 39692 1431 39748
rect 1487 39692 1555 39748
rect 1611 39692 1679 39748
rect 1735 39692 1803 39748
rect 1859 39692 1927 39748
rect 1983 39692 2051 39748
rect 2107 39692 2117 39748
rect 305 39624 2117 39692
rect 305 39568 315 39624
rect 371 39568 439 39624
rect 495 39568 563 39624
rect 619 39568 687 39624
rect 743 39568 811 39624
rect 867 39568 935 39624
rect 991 39568 1059 39624
rect 1115 39568 1183 39624
rect 1239 39568 1307 39624
rect 1363 39568 1431 39624
rect 1487 39568 1555 39624
rect 1611 39568 1679 39624
rect 1735 39568 1803 39624
rect 1859 39568 1927 39624
rect 1983 39568 2051 39624
rect 2107 39568 2117 39624
rect 305 39500 2117 39568
rect 305 39444 315 39500
rect 371 39444 439 39500
rect 495 39444 563 39500
rect 619 39444 687 39500
rect 743 39444 811 39500
rect 867 39444 935 39500
rect 991 39444 1059 39500
rect 1115 39444 1183 39500
rect 1239 39444 1307 39500
rect 1363 39444 1431 39500
rect 1487 39444 1555 39500
rect 1611 39444 1679 39500
rect 1735 39444 1803 39500
rect 1859 39444 1927 39500
rect 1983 39444 2051 39500
rect 2107 39444 2117 39500
rect 305 39376 2117 39444
rect 305 39320 315 39376
rect 371 39320 439 39376
rect 495 39320 563 39376
rect 619 39320 687 39376
rect 743 39320 811 39376
rect 867 39320 935 39376
rect 991 39320 1059 39376
rect 1115 39320 1183 39376
rect 1239 39320 1307 39376
rect 1363 39320 1431 39376
rect 1487 39320 1555 39376
rect 1611 39320 1679 39376
rect 1735 39320 1803 39376
rect 1859 39320 1927 39376
rect 1983 39320 2051 39376
rect 2107 39320 2117 39376
rect 305 39252 2117 39320
rect 305 39196 315 39252
rect 371 39196 439 39252
rect 495 39196 563 39252
rect 619 39196 687 39252
rect 743 39196 811 39252
rect 867 39196 935 39252
rect 991 39196 1059 39252
rect 1115 39196 1183 39252
rect 1239 39196 1307 39252
rect 1363 39196 1431 39252
rect 1487 39196 1555 39252
rect 1611 39196 1679 39252
rect 1735 39196 1803 39252
rect 1859 39196 1927 39252
rect 1983 39196 2051 39252
rect 2107 39196 2117 39252
rect 305 39128 2117 39196
rect 305 39072 315 39128
rect 371 39072 439 39128
rect 495 39072 563 39128
rect 619 39072 687 39128
rect 743 39072 811 39128
rect 867 39072 935 39128
rect 991 39072 1059 39128
rect 1115 39072 1183 39128
rect 1239 39072 1307 39128
rect 1363 39072 1431 39128
rect 1487 39072 1555 39128
rect 1611 39072 1679 39128
rect 1735 39072 1803 39128
rect 1859 39072 1927 39128
rect 1983 39072 2051 39128
rect 2107 39072 2117 39128
rect 305 39004 2117 39072
rect 305 38948 315 39004
rect 371 38948 439 39004
rect 495 38948 563 39004
rect 619 38948 687 39004
rect 743 38948 811 39004
rect 867 38948 935 39004
rect 991 38948 1059 39004
rect 1115 38948 1183 39004
rect 1239 38948 1307 39004
rect 1363 38948 1431 39004
rect 1487 38948 1555 39004
rect 1611 38948 1679 39004
rect 1735 38948 1803 39004
rect 1859 38948 1927 39004
rect 1983 38948 2051 39004
rect 2107 38948 2117 39004
rect 305 38880 2117 38948
rect 305 38824 315 38880
rect 371 38824 439 38880
rect 495 38824 563 38880
rect 619 38824 687 38880
rect 743 38824 811 38880
rect 867 38824 935 38880
rect 991 38824 1059 38880
rect 1115 38824 1183 38880
rect 1239 38824 1307 38880
rect 1363 38824 1431 38880
rect 1487 38824 1555 38880
rect 1611 38824 1679 38880
rect 1735 38824 1803 38880
rect 1859 38824 1927 38880
rect 1983 38824 2051 38880
rect 2107 38824 2117 38880
rect 305 38756 2117 38824
rect 305 38700 315 38756
rect 371 38700 439 38756
rect 495 38700 563 38756
rect 619 38700 687 38756
rect 743 38700 811 38756
rect 867 38700 935 38756
rect 991 38700 1059 38756
rect 1115 38700 1183 38756
rect 1239 38700 1307 38756
rect 1363 38700 1431 38756
rect 1487 38700 1555 38756
rect 1611 38700 1679 38756
rect 1735 38700 1803 38756
rect 1859 38700 1927 38756
rect 1983 38700 2051 38756
rect 2107 38700 2117 38756
rect 305 38632 2117 38700
rect 305 38576 315 38632
rect 371 38576 439 38632
rect 495 38576 563 38632
rect 619 38576 687 38632
rect 743 38576 811 38632
rect 867 38576 935 38632
rect 991 38576 1059 38632
rect 1115 38576 1183 38632
rect 1239 38576 1307 38632
rect 1363 38576 1431 38632
rect 1487 38576 1555 38632
rect 1611 38576 1679 38632
rect 1735 38576 1803 38632
rect 1859 38576 1927 38632
rect 1983 38576 2051 38632
rect 2107 38576 2117 38632
rect 305 38508 2117 38576
rect 305 38452 315 38508
rect 371 38452 439 38508
rect 495 38452 563 38508
rect 619 38452 687 38508
rect 743 38452 811 38508
rect 867 38452 935 38508
rect 991 38452 1059 38508
rect 1115 38452 1183 38508
rect 1239 38452 1307 38508
rect 1363 38452 1431 38508
rect 1487 38452 1555 38508
rect 1611 38452 1679 38508
rect 1735 38452 1803 38508
rect 1859 38452 1927 38508
rect 1983 38452 2051 38508
rect 2107 38452 2117 38508
rect 305 38442 2117 38452
rect -11 38176 86 38200
rect -11 36824 20 38176
rect 76 36824 86 38176
rect -11 36800 86 36824
rect 2279 38135 2355 51277
rect 2481 49348 2681 52852
rect 2481 49292 2491 49348
rect 2547 49292 2615 49348
rect 2671 49292 2681 49348
rect 2481 49224 2681 49292
rect 2481 49168 2491 49224
rect 2547 49168 2615 49224
rect 2671 49168 2681 49224
rect 2481 49100 2681 49168
rect 2481 49044 2491 49100
rect 2547 49044 2615 49100
rect 2671 49044 2681 49100
rect 2481 48976 2681 49044
rect 2481 48920 2491 48976
rect 2547 48920 2615 48976
rect 2671 48920 2681 48976
rect 2481 48852 2681 48920
rect 2481 48796 2491 48852
rect 2547 48796 2615 48852
rect 2671 48796 2681 48852
rect 2481 48728 2681 48796
rect 2481 48672 2491 48728
rect 2547 48672 2615 48728
rect 2671 48672 2681 48728
rect 2481 48604 2681 48672
rect 2481 48548 2491 48604
rect 2547 48548 2615 48604
rect 2671 48548 2681 48604
rect 2481 48480 2681 48548
rect 2481 48424 2491 48480
rect 2547 48424 2615 48480
rect 2671 48424 2681 48480
rect 2481 48356 2681 48424
rect 2481 48300 2491 48356
rect 2547 48300 2615 48356
rect 2671 48300 2681 48356
rect 2481 48232 2681 48300
rect 2481 48176 2491 48232
rect 2547 48176 2615 48232
rect 2671 48176 2681 48232
rect 2481 48108 2681 48176
rect 2481 48052 2491 48108
rect 2547 48052 2615 48108
rect 2671 48052 2681 48108
rect 2481 47281 2681 48052
rect 2741 56669 4791 57600
rect 2741 56617 2833 56669
rect 2885 56617 2957 56669
rect 3009 56617 3081 56669
rect 3133 56617 3205 56669
rect 3257 56617 3329 56669
rect 3381 56617 3453 56669
rect 3505 56617 3577 56669
rect 3629 56617 3701 56669
rect 3753 56617 4340 56669
rect 4392 56617 4464 56669
rect 4516 56617 4588 56669
rect 4640 56617 4712 56669
rect 4764 56617 4791 56669
rect 2741 56545 4791 56617
rect 2741 56493 2833 56545
rect 2885 56493 2957 56545
rect 3009 56493 3081 56545
rect 3133 56493 3205 56545
rect 3257 56493 3329 56545
rect 3381 56493 3453 56545
rect 3505 56493 3577 56545
rect 3629 56493 3701 56545
rect 3753 56493 4340 56545
rect 4392 56493 4464 56545
rect 4516 56493 4588 56545
rect 4640 56493 4712 56545
rect 4764 56493 4791 56545
rect 2741 56421 4791 56493
rect 2741 56369 2833 56421
rect 2885 56369 2957 56421
rect 3009 56369 3081 56421
rect 3133 56369 3205 56421
rect 3257 56369 3329 56421
rect 3381 56369 3453 56421
rect 3505 56369 3577 56421
rect 3629 56369 3701 56421
rect 3753 56369 4340 56421
rect 4392 56369 4464 56421
rect 4516 56369 4588 56421
rect 4640 56369 4712 56421
rect 4764 56369 4791 56421
rect 2741 56297 4791 56369
rect 2741 56245 2833 56297
rect 2885 56245 2957 56297
rect 3009 56245 3081 56297
rect 3133 56245 3205 56297
rect 3257 56245 3329 56297
rect 3381 56245 3453 56297
rect 3505 56245 3577 56297
rect 3629 56245 3701 56297
rect 3753 56245 4340 56297
rect 4392 56245 4464 56297
rect 4516 56245 4588 56297
rect 4640 56245 4712 56297
rect 4764 56245 4791 56297
rect 2741 56173 4791 56245
rect 2741 56121 2833 56173
rect 2885 56121 2957 56173
rect 3009 56121 3081 56173
rect 3133 56121 3205 56173
rect 3257 56121 3329 56173
rect 3381 56121 3453 56173
rect 3505 56121 3577 56173
rect 3629 56121 3701 56173
rect 3753 56121 4340 56173
rect 4392 56121 4464 56173
rect 4516 56121 4588 56173
rect 4640 56121 4712 56173
rect 4764 56121 4791 56173
rect 2741 56049 4791 56121
rect 2741 55997 2833 56049
rect 2885 55997 2957 56049
rect 3009 55997 3081 56049
rect 3133 55997 3205 56049
rect 3257 55997 3329 56049
rect 3381 55997 3453 56049
rect 3505 55997 3577 56049
rect 3629 55997 3701 56049
rect 3753 55997 4340 56049
rect 4392 55997 4464 56049
rect 4516 55997 4588 56049
rect 4640 55997 4712 56049
rect 4764 55997 4791 56049
rect 2741 55925 4791 55997
rect 2741 55873 2833 55925
rect 2885 55873 2957 55925
rect 3009 55873 3081 55925
rect 3133 55873 3205 55925
rect 3257 55873 3329 55925
rect 3381 55873 3453 55925
rect 3505 55873 3577 55925
rect 3629 55873 3701 55925
rect 3753 55873 4340 55925
rect 4392 55873 4464 55925
rect 4516 55873 4588 55925
rect 4640 55873 4712 55925
rect 4764 55873 4791 55925
rect 2741 55801 4791 55873
rect 2741 55749 2833 55801
rect 2885 55749 2957 55801
rect 3009 55749 3081 55801
rect 3133 55749 3205 55801
rect 3257 55749 3329 55801
rect 3381 55749 3453 55801
rect 3505 55749 3577 55801
rect 3629 55749 3701 55801
rect 3753 55749 4340 55801
rect 4392 55749 4464 55801
rect 4516 55749 4588 55801
rect 4640 55749 4712 55801
rect 4764 55749 4791 55801
rect 2741 55748 4791 55749
rect 2741 55692 2808 55748
rect 2864 55692 2932 55748
rect 2988 55692 3056 55748
rect 3112 55692 3180 55748
rect 3236 55692 3304 55748
rect 3360 55692 3428 55748
rect 3484 55692 3552 55748
rect 3608 55692 3676 55748
rect 3732 55692 3800 55748
rect 3856 55692 3924 55748
rect 3980 55692 4048 55748
rect 4104 55692 4172 55748
rect 4228 55692 4296 55748
rect 4352 55692 4420 55748
rect 4476 55692 4544 55748
rect 4600 55692 4668 55748
rect 4724 55692 4791 55748
rect 2741 55677 4791 55692
rect 2741 55625 2833 55677
rect 2885 55625 2957 55677
rect 3009 55625 3081 55677
rect 3133 55625 3205 55677
rect 3257 55625 3329 55677
rect 3381 55625 3453 55677
rect 3505 55625 3577 55677
rect 3629 55625 3701 55677
rect 3753 55625 4340 55677
rect 4392 55625 4464 55677
rect 4516 55625 4588 55677
rect 4640 55625 4712 55677
rect 4764 55625 4791 55677
rect 2741 55624 4791 55625
rect 2741 55568 2808 55624
rect 2864 55568 2932 55624
rect 2988 55568 3056 55624
rect 3112 55568 3180 55624
rect 3236 55568 3304 55624
rect 3360 55568 3428 55624
rect 3484 55568 3552 55624
rect 3608 55568 3676 55624
rect 3732 55568 3800 55624
rect 3856 55568 3924 55624
rect 3980 55568 4048 55624
rect 4104 55568 4172 55624
rect 4228 55568 4296 55624
rect 4352 55568 4420 55624
rect 4476 55568 4544 55624
rect 4600 55568 4668 55624
rect 4724 55568 4791 55624
rect 2741 55553 4791 55568
rect 2741 55501 2833 55553
rect 2885 55501 2957 55553
rect 3009 55501 3081 55553
rect 3133 55501 3205 55553
rect 3257 55501 3329 55553
rect 3381 55501 3453 55553
rect 3505 55501 3577 55553
rect 3629 55501 3701 55553
rect 3753 55501 4340 55553
rect 4392 55501 4464 55553
rect 4516 55501 4588 55553
rect 4640 55501 4712 55553
rect 4764 55501 4791 55553
rect 2741 55500 4791 55501
rect 2741 55444 2808 55500
rect 2864 55444 2932 55500
rect 2988 55444 3056 55500
rect 3112 55444 3180 55500
rect 3236 55444 3304 55500
rect 3360 55444 3428 55500
rect 3484 55444 3552 55500
rect 3608 55444 3676 55500
rect 3732 55444 3800 55500
rect 3856 55444 3924 55500
rect 3980 55444 4048 55500
rect 4104 55444 4172 55500
rect 4228 55444 4296 55500
rect 4352 55444 4420 55500
rect 4476 55444 4544 55500
rect 4600 55444 4668 55500
rect 4724 55444 4791 55500
rect 2741 55429 4791 55444
rect 2741 55377 2833 55429
rect 2885 55377 2957 55429
rect 3009 55377 3081 55429
rect 3133 55377 3205 55429
rect 3257 55377 3329 55429
rect 3381 55377 3453 55429
rect 3505 55377 3577 55429
rect 3629 55377 3701 55429
rect 3753 55377 4340 55429
rect 4392 55377 4464 55429
rect 4516 55377 4588 55429
rect 4640 55377 4712 55429
rect 4764 55377 4791 55429
rect 2741 55376 4791 55377
rect 2741 55320 2808 55376
rect 2864 55320 2932 55376
rect 2988 55320 3056 55376
rect 3112 55320 3180 55376
rect 3236 55320 3304 55376
rect 3360 55320 3428 55376
rect 3484 55320 3552 55376
rect 3608 55320 3676 55376
rect 3732 55320 3800 55376
rect 3856 55320 3924 55376
rect 3980 55320 4048 55376
rect 4104 55320 4172 55376
rect 4228 55320 4296 55376
rect 4352 55320 4420 55376
rect 4476 55320 4544 55376
rect 4600 55320 4668 55376
rect 4724 55320 4791 55376
rect 2741 55305 4791 55320
rect 2741 55253 2833 55305
rect 2885 55253 2957 55305
rect 3009 55253 3081 55305
rect 3133 55253 3205 55305
rect 3257 55253 3329 55305
rect 3381 55253 3453 55305
rect 3505 55253 3577 55305
rect 3629 55253 3701 55305
rect 3753 55253 4340 55305
rect 4392 55253 4464 55305
rect 4516 55253 4588 55305
rect 4640 55253 4712 55305
rect 4764 55253 4791 55305
rect 2741 55252 4791 55253
rect 2741 55196 2808 55252
rect 2864 55196 2932 55252
rect 2988 55196 3056 55252
rect 3112 55196 3180 55252
rect 3236 55196 3304 55252
rect 3360 55196 3428 55252
rect 3484 55196 3552 55252
rect 3608 55196 3676 55252
rect 3732 55196 3800 55252
rect 3856 55196 3924 55252
rect 3980 55196 4048 55252
rect 4104 55196 4172 55252
rect 4228 55196 4296 55252
rect 4352 55196 4420 55252
rect 4476 55196 4544 55252
rect 4600 55196 4668 55252
rect 4724 55196 4791 55252
rect 2741 55181 4791 55196
rect 2741 55129 2833 55181
rect 2885 55129 2957 55181
rect 3009 55129 3081 55181
rect 3133 55129 3205 55181
rect 3257 55129 3329 55181
rect 3381 55129 3453 55181
rect 3505 55129 3577 55181
rect 3629 55129 3701 55181
rect 3753 55129 4340 55181
rect 4392 55129 4464 55181
rect 4516 55129 4588 55181
rect 4640 55129 4712 55181
rect 4764 55129 4791 55181
rect 2741 55128 4791 55129
rect 2741 55072 2808 55128
rect 2864 55072 2932 55128
rect 2988 55072 3056 55128
rect 3112 55072 3180 55128
rect 3236 55072 3304 55128
rect 3360 55072 3428 55128
rect 3484 55072 3552 55128
rect 3608 55072 3676 55128
rect 3732 55072 3800 55128
rect 3856 55072 3924 55128
rect 3980 55072 4048 55128
rect 4104 55072 4172 55128
rect 4228 55072 4296 55128
rect 4352 55072 4420 55128
rect 4476 55072 4544 55128
rect 4600 55072 4668 55128
rect 4724 55072 4791 55128
rect 2741 55057 4791 55072
rect 2741 55005 2833 55057
rect 2885 55005 2957 55057
rect 3009 55005 3081 55057
rect 3133 55005 3205 55057
rect 3257 55005 3329 55057
rect 3381 55005 3453 55057
rect 3505 55005 3577 55057
rect 3629 55005 3701 55057
rect 3753 55005 4340 55057
rect 4392 55005 4464 55057
rect 4516 55005 4588 55057
rect 4640 55005 4712 55057
rect 4764 55005 4791 55057
rect 2741 55004 4791 55005
rect 2741 54948 2808 55004
rect 2864 54948 2932 55004
rect 2988 54948 3056 55004
rect 3112 54948 3180 55004
rect 3236 54948 3304 55004
rect 3360 54948 3428 55004
rect 3484 54948 3552 55004
rect 3608 54948 3676 55004
rect 3732 54948 3800 55004
rect 3856 54948 3924 55004
rect 3980 54948 4048 55004
rect 4104 54948 4172 55004
rect 4228 54948 4296 55004
rect 4352 54948 4420 55004
rect 4476 54948 4544 55004
rect 4600 54948 4668 55004
rect 4724 54948 4791 55004
rect 2741 54933 4791 54948
rect 2741 54881 2833 54933
rect 2885 54881 2957 54933
rect 3009 54881 3081 54933
rect 3133 54881 3205 54933
rect 3257 54881 3329 54933
rect 3381 54881 3453 54933
rect 3505 54881 3577 54933
rect 3629 54881 3701 54933
rect 3753 54881 4340 54933
rect 4392 54881 4464 54933
rect 4516 54881 4588 54933
rect 4640 54881 4712 54933
rect 4764 54881 4791 54933
rect 2741 54880 4791 54881
rect 2741 54824 2808 54880
rect 2864 54824 2932 54880
rect 2988 54824 3056 54880
rect 3112 54824 3180 54880
rect 3236 54824 3304 54880
rect 3360 54824 3428 54880
rect 3484 54824 3552 54880
rect 3608 54824 3676 54880
rect 3732 54824 3800 54880
rect 3856 54824 3924 54880
rect 3980 54824 4048 54880
rect 4104 54824 4172 54880
rect 4228 54824 4296 54880
rect 4352 54824 4420 54880
rect 4476 54824 4544 54880
rect 4600 54824 4668 54880
rect 4724 54824 4791 54880
rect 2741 54809 4791 54824
rect 2741 54757 2833 54809
rect 2885 54757 2957 54809
rect 3009 54757 3081 54809
rect 3133 54757 3205 54809
rect 3257 54757 3329 54809
rect 3381 54757 3453 54809
rect 3505 54757 3577 54809
rect 3629 54757 3701 54809
rect 3753 54757 4340 54809
rect 4392 54757 4464 54809
rect 4516 54757 4588 54809
rect 4640 54757 4712 54809
rect 4764 54757 4791 54809
rect 2741 54756 4791 54757
rect 2741 54700 2808 54756
rect 2864 54700 2932 54756
rect 2988 54700 3056 54756
rect 3112 54700 3180 54756
rect 3236 54700 3304 54756
rect 3360 54700 3428 54756
rect 3484 54700 3552 54756
rect 3608 54700 3676 54756
rect 3732 54700 3800 54756
rect 3856 54700 3924 54756
rect 3980 54700 4048 54756
rect 4104 54700 4172 54756
rect 4228 54700 4296 54756
rect 4352 54700 4420 54756
rect 4476 54700 4544 54756
rect 4600 54700 4668 54756
rect 4724 54700 4791 54756
rect 2741 54685 4791 54700
rect 2741 54633 2833 54685
rect 2885 54633 2957 54685
rect 3009 54633 3081 54685
rect 3133 54633 3205 54685
rect 3257 54633 3329 54685
rect 3381 54633 3453 54685
rect 3505 54633 3577 54685
rect 3629 54633 3701 54685
rect 3753 54633 4340 54685
rect 4392 54633 4464 54685
rect 4516 54633 4588 54685
rect 4640 54633 4712 54685
rect 4764 54633 4791 54685
rect 2741 54632 4791 54633
rect 2741 54576 2808 54632
rect 2864 54576 2932 54632
rect 2988 54576 3056 54632
rect 3112 54576 3180 54632
rect 3236 54576 3304 54632
rect 3360 54576 3428 54632
rect 3484 54576 3552 54632
rect 3608 54576 3676 54632
rect 3732 54576 3800 54632
rect 3856 54576 3924 54632
rect 3980 54576 4048 54632
rect 4104 54576 4172 54632
rect 4228 54576 4296 54632
rect 4352 54576 4420 54632
rect 4476 54576 4544 54632
rect 4600 54576 4668 54632
rect 4724 54576 4791 54632
rect 2741 54561 4791 54576
rect 2741 54509 2833 54561
rect 2885 54509 2957 54561
rect 3009 54509 3081 54561
rect 3133 54509 3205 54561
rect 3257 54509 3329 54561
rect 3381 54509 3453 54561
rect 3505 54509 3577 54561
rect 3629 54509 3701 54561
rect 3753 54509 4340 54561
rect 4392 54509 4464 54561
rect 4516 54509 4588 54561
rect 4640 54509 4712 54561
rect 4764 54509 4791 54561
rect 2741 54508 4791 54509
rect 2741 54452 2808 54508
rect 2864 54452 2932 54508
rect 2988 54452 3056 54508
rect 3112 54452 3180 54508
rect 3236 54452 3304 54508
rect 3360 54452 3428 54508
rect 3484 54452 3552 54508
rect 3608 54452 3676 54508
rect 3732 54452 3800 54508
rect 3856 54452 3924 54508
rect 3980 54452 4048 54508
rect 4104 54452 4172 54508
rect 4228 54452 4296 54508
rect 4352 54452 4420 54508
rect 4476 54452 4544 54508
rect 4600 54452 4668 54508
rect 4724 54452 4791 54508
rect 2741 54437 4791 54452
rect 2741 54385 2833 54437
rect 2885 54385 2957 54437
rect 3009 54385 3081 54437
rect 3133 54385 3205 54437
rect 3257 54385 3329 54437
rect 3381 54385 3453 54437
rect 3505 54385 3577 54437
rect 3629 54385 3701 54437
rect 3753 54385 4340 54437
rect 4392 54385 4464 54437
rect 4516 54385 4588 54437
rect 4640 54385 4712 54437
rect 4764 54385 4791 54437
rect 2741 54313 4791 54385
rect 2741 54261 2833 54313
rect 2885 54261 2957 54313
rect 3009 54261 3081 54313
rect 3133 54261 3205 54313
rect 3257 54261 3329 54313
rect 3381 54261 3453 54313
rect 3505 54261 3577 54313
rect 3629 54261 3701 54313
rect 3753 54261 4340 54313
rect 4392 54261 4464 54313
rect 4516 54261 4588 54313
rect 4640 54261 4712 54313
rect 4764 54261 4791 54313
rect 2741 54189 4791 54261
rect 2741 54137 2833 54189
rect 2885 54137 2957 54189
rect 3009 54137 3081 54189
rect 3133 54137 3205 54189
rect 3257 54137 3329 54189
rect 3381 54137 3453 54189
rect 3505 54137 3577 54189
rect 3629 54137 3701 54189
rect 3753 54137 4340 54189
rect 4392 54137 4464 54189
rect 4516 54137 4588 54189
rect 4640 54137 4712 54189
rect 4764 54137 4791 54189
rect 2741 54065 4791 54137
rect 2741 54013 2833 54065
rect 2885 54013 2957 54065
rect 3009 54013 3081 54065
rect 3133 54013 3205 54065
rect 3257 54013 3329 54065
rect 3381 54013 3453 54065
rect 3505 54013 3577 54065
rect 3629 54013 3701 54065
rect 3753 54013 4340 54065
rect 4392 54013 4464 54065
rect 4516 54013 4588 54065
rect 4640 54013 4712 54065
rect 4764 54013 4791 54065
rect 2741 53941 4791 54013
rect 2741 53889 2833 53941
rect 2885 53889 2957 53941
rect 3009 53889 3081 53941
rect 3133 53889 3205 53941
rect 3257 53889 3329 53941
rect 3381 53889 3453 53941
rect 3505 53889 3577 53941
rect 3629 53889 3701 53941
rect 3753 53889 4340 53941
rect 4392 53889 4464 53941
rect 4516 53889 4588 53941
rect 4640 53889 4712 53941
rect 4764 53889 4791 53941
rect 2741 53817 4791 53889
rect 2741 53765 2833 53817
rect 2885 53765 2957 53817
rect 3009 53765 3081 53817
rect 3133 53765 3205 53817
rect 3257 53765 3329 53817
rect 3381 53765 3453 53817
rect 3505 53765 3577 53817
rect 3629 53765 3701 53817
rect 3753 53765 4340 53817
rect 4392 53765 4464 53817
rect 4516 53765 4588 53817
rect 4640 53765 4712 53817
rect 4764 53765 4791 53817
rect 2741 53693 4791 53765
rect 2741 53641 2833 53693
rect 2885 53641 2957 53693
rect 3009 53641 3081 53693
rect 3133 53641 3205 53693
rect 3257 53641 3329 53693
rect 3381 53641 3453 53693
rect 3505 53641 3577 53693
rect 3629 53641 3701 53693
rect 3753 53641 4340 53693
rect 4392 53641 4464 53693
rect 4516 53641 4588 53693
rect 4640 53641 4712 53693
rect 4764 53641 4791 53693
rect 2741 52588 4791 53641
rect 2741 52536 2810 52588
rect 2862 52536 2934 52588
rect 2986 52536 3058 52588
rect 3110 52536 3182 52588
rect 3234 52536 3306 52588
rect 3358 52536 3430 52588
rect 3482 52536 3554 52588
rect 3606 52536 3678 52588
rect 3730 52536 3802 52588
rect 3854 52536 3926 52588
rect 3978 52536 4050 52588
rect 4102 52536 4174 52588
rect 4226 52536 4298 52588
rect 4350 52536 4422 52588
rect 4474 52536 4546 52588
rect 4598 52536 4670 52588
rect 4722 52536 4791 52588
rect 2741 52464 4791 52536
rect 2741 52412 2810 52464
rect 2862 52412 2934 52464
rect 2986 52412 3058 52464
rect 3110 52412 3182 52464
rect 3234 52412 3306 52464
rect 3358 52412 3430 52464
rect 3482 52412 3554 52464
rect 3606 52412 3678 52464
rect 3730 52412 3802 52464
rect 3854 52412 3926 52464
rect 3978 52412 4050 52464
rect 4102 52412 4174 52464
rect 4226 52412 4298 52464
rect 4350 52412 4422 52464
rect 4474 52412 4546 52464
rect 4598 52412 4670 52464
rect 4722 52412 4791 52464
rect 2741 52340 4791 52412
rect 2741 52288 2810 52340
rect 2862 52288 2934 52340
rect 2986 52288 3058 52340
rect 3110 52288 3182 52340
rect 3234 52288 3306 52340
rect 3358 52288 3430 52340
rect 3482 52288 3554 52340
rect 3606 52288 3678 52340
rect 3730 52288 3802 52340
rect 3854 52288 3926 52340
rect 3978 52288 4050 52340
rect 4102 52288 4174 52340
rect 4226 52288 4298 52340
rect 4350 52288 4422 52340
rect 4474 52288 4546 52340
rect 4598 52288 4670 52340
rect 4722 52288 4791 52340
rect 2741 51627 4791 52288
rect 2741 51575 3559 51627
rect 3611 51575 3683 51627
rect 3735 51575 3807 51627
rect 3859 51575 3931 51627
rect 3983 51575 4055 51627
rect 4107 51575 4179 51627
rect 4231 51575 4303 51627
rect 4355 51575 4427 51627
rect 4479 51575 4551 51627
rect 4603 51575 4675 51627
rect 4727 51575 4791 51627
rect 2741 51503 4791 51575
rect 2741 51451 3559 51503
rect 3611 51451 3683 51503
rect 3735 51451 3807 51503
rect 3859 51451 3931 51503
rect 3983 51451 4055 51503
rect 4107 51451 4179 51503
rect 4231 51451 4303 51503
rect 4355 51451 4427 51503
rect 4479 51451 4551 51503
rect 4603 51451 4675 51503
rect 4727 51451 4791 51503
rect 2741 50948 4791 51451
rect 2741 50892 2808 50948
rect 2864 50892 2932 50948
rect 2988 50892 3056 50948
rect 3112 50892 3180 50948
rect 3236 50892 3304 50948
rect 3360 50892 3428 50948
rect 3484 50892 3552 50948
rect 3608 50892 3676 50948
rect 3732 50892 3800 50948
rect 3856 50892 3924 50948
rect 3980 50892 4048 50948
rect 4104 50892 4172 50948
rect 4228 50892 4296 50948
rect 4352 50892 4420 50948
rect 4476 50892 4544 50948
rect 4600 50892 4668 50948
rect 4724 50892 4791 50948
rect 2741 50824 4791 50892
rect 2741 50768 2808 50824
rect 2864 50768 2932 50824
rect 2988 50768 3056 50824
rect 3112 50768 3180 50824
rect 3236 50768 3304 50824
rect 3360 50768 3428 50824
rect 3484 50768 3552 50824
rect 3608 50768 3676 50824
rect 3732 50768 3800 50824
rect 3856 50768 3924 50824
rect 3980 50768 4048 50824
rect 4104 50768 4172 50824
rect 4228 50768 4296 50824
rect 4352 50768 4420 50824
rect 4476 50768 4544 50824
rect 4600 50768 4668 50824
rect 4724 50768 4791 50824
rect 2741 50700 4791 50768
rect 2741 50644 2808 50700
rect 2864 50644 2932 50700
rect 2988 50644 3056 50700
rect 3112 50644 3180 50700
rect 3236 50644 3304 50700
rect 3360 50644 3428 50700
rect 3484 50644 3552 50700
rect 3608 50693 3676 50700
rect 3732 50693 3800 50700
rect 3856 50693 3924 50700
rect 3980 50693 4048 50700
rect 4104 50693 4172 50700
rect 4228 50693 4296 50700
rect 4352 50693 4420 50700
rect 4476 50693 4544 50700
rect 4600 50693 4668 50700
rect 4724 50693 4791 50700
rect 3611 50644 3676 50693
rect 3735 50644 3800 50693
rect 3859 50644 3924 50693
rect 3983 50644 4048 50693
rect 4107 50644 4172 50693
rect 4231 50644 4296 50693
rect 4355 50644 4420 50693
rect 4479 50644 4544 50693
rect 4603 50644 4668 50693
rect 2741 50641 3559 50644
rect 3611 50641 3683 50644
rect 3735 50641 3807 50644
rect 3859 50641 3931 50644
rect 3983 50641 4055 50644
rect 4107 50641 4179 50644
rect 4231 50641 4303 50644
rect 4355 50641 4427 50644
rect 4479 50641 4551 50644
rect 4603 50641 4675 50644
rect 4727 50641 4791 50693
rect 2741 50576 4791 50641
rect 2741 50520 2808 50576
rect 2864 50520 2932 50576
rect 2988 50520 3056 50576
rect 3112 50520 3180 50576
rect 3236 50520 3304 50576
rect 3360 50520 3428 50576
rect 3484 50520 3552 50576
rect 3608 50569 3676 50576
rect 3732 50569 3800 50576
rect 3856 50569 3924 50576
rect 3980 50569 4048 50576
rect 4104 50569 4172 50576
rect 4228 50569 4296 50576
rect 4352 50569 4420 50576
rect 4476 50569 4544 50576
rect 4600 50569 4668 50576
rect 4724 50569 4791 50576
rect 3611 50520 3676 50569
rect 3735 50520 3800 50569
rect 3859 50520 3924 50569
rect 3983 50520 4048 50569
rect 4107 50520 4172 50569
rect 4231 50520 4296 50569
rect 4355 50520 4420 50569
rect 4479 50520 4544 50569
rect 4603 50520 4668 50569
rect 2741 50517 3559 50520
rect 3611 50517 3683 50520
rect 3735 50517 3807 50520
rect 3859 50517 3931 50520
rect 3983 50517 4055 50520
rect 4107 50517 4179 50520
rect 4231 50517 4303 50520
rect 4355 50517 4427 50520
rect 4479 50517 4551 50520
rect 4603 50517 4675 50520
rect 4727 50517 4791 50569
rect 2741 50452 4791 50517
rect 2741 50396 2808 50452
rect 2864 50396 2932 50452
rect 2988 50396 3056 50452
rect 3112 50396 3180 50452
rect 3236 50396 3304 50452
rect 3360 50396 3428 50452
rect 3484 50396 3552 50452
rect 3608 50396 3676 50452
rect 3732 50396 3800 50452
rect 3856 50396 3924 50452
rect 3980 50396 4048 50452
rect 4104 50396 4172 50452
rect 4228 50396 4296 50452
rect 4352 50396 4420 50452
rect 4476 50396 4544 50452
rect 4600 50396 4668 50452
rect 4724 50396 4791 50452
rect 2741 50328 4791 50396
rect 2741 50272 2808 50328
rect 2864 50272 2932 50328
rect 2988 50272 3056 50328
rect 3112 50272 3180 50328
rect 3236 50272 3304 50328
rect 3360 50272 3428 50328
rect 3484 50272 3552 50328
rect 3608 50272 3676 50328
rect 3732 50272 3800 50328
rect 3856 50272 3924 50328
rect 3980 50272 4048 50328
rect 4104 50272 4172 50328
rect 4228 50272 4296 50328
rect 4352 50272 4420 50328
rect 4476 50272 4544 50328
rect 4600 50272 4668 50328
rect 4724 50272 4791 50328
rect 2741 50204 4791 50272
rect 2741 50148 2808 50204
rect 2864 50148 2932 50204
rect 2988 50148 3056 50204
rect 3112 50148 3180 50204
rect 3236 50148 3304 50204
rect 3360 50148 3428 50204
rect 3484 50148 3552 50204
rect 3608 50148 3676 50204
rect 3732 50148 3800 50204
rect 3856 50148 3924 50204
rect 3980 50148 4048 50204
rect 4104 50148 4172 50204
rect 4228 50148 4296 50204
rect 4352 50148 4420 50204
rect 4476 50148 4544 50204
rect 4600 50148 4668 50204
rect 4724 50148 4791 50204
rect 2741 50080 4791 50148
rect 2741 50024 2808 50080
rect 2864 50024 2932 50080
rect 2988 50024 3056 50080
rect 3112 50024 3180 50080
rect 3236 50024 3304 50080
rect 3360 50024 3428 50080
rect 3484 50024 3552 50080
rect 3608 50024 3676 50080
rect 3732 50024 3800 50080
rect 3856 50024 3924 50080
rect 3980 50024 4048 50080
rect 4104 50024 4172 50080
rect 4228 50024 4296 50080
rect 4352 50024 4420 50080
rect 4476 50024 4544 50080
rect 4600 50024 4668 50080
rect 4724 50024 4791 50080
rect 2741 49956 4791 50024
rect 2741 49900 2808 49956
rect 2864 49900 2932 49956
rect 2988 49900 3056 49956
rect 3112 49900 3180 49956
rect 3236 49900 3304 49956
rect 3360 49900 3428 49956
rect 3484 49900 3552 49956
rect 3608 49900 3676 49956
rect 3732 49900 3800 49956
rect 3856 49900 3924 49956
rect 3980 49900 4048 49956
rect 4104 49900 4172 49956
rect 4228 49900 4296 49956
rect 4352 49900 4420 49956
rect 4476 49900 4544 49956
rect 4600 49900 4668 49956
rect 4724 49900 4791 49956
rect 2741 49832 4791 49900
rect 2741 49776 2808 49832
rect 2864 49776 2932 49832
rect 2988 49776 3056 49832
rect 3112 49776 3180 49832
rect 3236 49776 3304 49832
rect 3360 49776 3428 49832
rect 3484 49776 3552 49832
rect 3608 49776 3676 49832
rect 3732 49776 3800 49832
rect 3856 49776 3924 49832
rect 3980 49776 4048 49832
rect 4104 49776 4172 49832
rect 4228 49776 4296 49832
rect 4352 49776 4420 49832
rect 4476 49776 4544 49832
rect 4600 49776 4668 49832
rect 4724 49776 4791 49832
rect 2741 49759 4791 49776
rect 2741 49708 3559 49759
rect 3611 49708 3683 49759
rect 3735 49708 3807 49759
rect 3859 49708 3931 49759
rect 3983 49708 4055 49759
rect 4107 49708 4179 49759
rect 4231 49708 4303 49759
rect 4355 49708 4427 49759
rect 4479 49708 4551 49759
rect 4603 49708 4675 49759
rect 2741 49652 2808 49708
rect 2864 49652 2932 49708
rect 2988 49652 3056 49708
rect 3112 49652 3180 49708
rect 3236 49652 3304 49708
rect 3360 49652 3428 49708
rect 3484 49652 3552 49708
rect 3611 49707 3676 49708
rect 3735 49707 3800 49708
rect 3859 49707 3924 49708
rect 3983 49707 4048 49708
rect 4107 49707 4172 49708
rect 4231 49707 4296 49708
rect 4355 49707 4420 49708
rect 4479 49707 4544 49708
rect 4603 49707 4668 49708
rect 4727 49707 4791 49759
rect 3608 49652 3676 49707
rect 3732 49652 3800 49707
rect 3856 49652 3924 49707
rect 3980 49652 4048 49707
rect 4104 49652 4172 49707
rect 4228 49652 4296 49707
rect 4352 49652 4420 49707
rect 4476 49652 4544 49707
rect 4600 49652 4668 49707
rect 4724 49652 4791 49707
rect 2741 49635 4791 49652
rect 2741 49583 3559 49635
rect 3611 49583 3683 49635
rect 3735 49583 3807 49635
rect 3859 49583 3931 49635
rect 3983 49583 4055 49635
rect 4107 49583 4179 49635
rect 4231 49583 4303 49635
rect 4355 49583 4427 49635
rect 4479 49583 4551 49635
rect 4603 49583 4675 49635
rect 4727 49583 4791 49635
rect 2741 48825 4791 49583
rect 2741 48773 3559 48825
rect 3611 48773 3683 48825
rect 3735 48773 3807 48825
rect 3859 48773 3931 48825
rect 3983 48773 4055 48825
rect 4107 48773 4179 48825
rect 4231 48773 4303 48825
rect 4355 48773 4427 48825
rect 4479 48773 4551 48825
rect 4603 48773 4675 48825
rect 4727 48773 4791 48825
rect 2741 48701 4791 48773
rect 2741 48649 3559 48701
rect 3611 48649 3683 48701
rect 3735 48649 3807 48701
rect 3859 48649 3931 48701
rect 3983 48649 4055 48701
rect 4107 48649 4179 48701
rect 4231 48649 4303 48701
rect 4355 48649 4427 48701
rect 4479 48649 4551 48701
rect 4603 48649 4675 48701
rect 4727 48649 4791 48701
rect 2741 47988 4791 48649
rect 2741 47936 2810 47988
rect 2862 47936 2934 47988
rect 2986 47936 3058 47988
rect 3110 47936 3182 47988
rect 3234 47936 3306 47988
rect 3358 47936 3430 47988
rect 3482 47936 3554 47988
rect 3606 47936 3678 47988
rect 3730 47936 3802 47988
rect 3854 47936 3926 47988
rect 3978 47936 4050 47988
rect 4102 47936 4174 47988
rect 4226 47936 4298 47988
rect 4350 47936 4422 47988
rect 4474 47936 4546 47988
rect 4598 47936 4670 47988
rect 4722 47936 4791 47988
rect 2741 47864 4791 47936
rect 2741 47812 2810 47864
rect 2862 47812 2934 47864
rect 2986 47812 3058 47864
rect 3110 47812 3182 47864
rect 3234 47812 3306 47864
rect 3358 47812 3430 47864
rect 3482 47812 3554 47864
rect 3606 47812 3678 47864
rect 3730 47812 3802 47864
rect 3854 47812 3926 47864
rect 3978 47812 4050 47864
rect 4102 47812 4174 47864
rect 4226 47812 4298 47864
rect 4350 47812 4422 47864
rect 4474 47812 4546 47864
rect 4598 47812 4670 47864
rect 4722 47812 4791 47864
rect 2741 47748 4791 47812
rect 2741 47692 2808 47748
rect 2864 47692 2932 47748
rect 2988 47692 3056 47748
rect 3112 47692 3180 47748
rect 3236 47692 3304 47748
rect 3360 47692 3428 47748
rect 3484 47692 3552 47748
rect 3608 47692 3676 47748
rect 3732 47692 3800 47748
rect 3856 47692 3924 47748
rect 3980 47692 4048 47748
rect 4104 47692 4172 47748
rect 4228 47692 4296 47748
rect 4352 47692 4420 47748
rect 4476 47692 4544 47748
rect 4600 47692 4668 47748
rect 4724 47692 4791 47748
rect 2741 47688 2810 47692
rect 2862 47688 2934 47692
rect 2986 47688 3058 47692
rect 3110 47688 3182 47692
rect 3234 47688 3306 47692
rect 3358 47688 3430 47692
rect 3482 47688 3554 47692
rect 3606 47688 3678 47692
rect 3730 47688 3802 47692
rect 3854 47688 3926 47692
rect 3978 47688 4050 47692
rect 4102 47688 4174 47692
rect 4226 47688 4298 47692
rect 4350 47688 4422 47692
rect 4474 47688 4546 47692
rect 4598 47688 4670 47692
rect 4722 47688 4791 47692
rect 2741 47624 4791 47688
rect 2741 47568 2808 47624
rect 2864 47568 2932 47624
rect 2988 47568 3056 47624
rect 3112 47568 3180 47624
rect 3236 47568 3304 47624
rect 3360 47568 3428 47624
rect 3484 47568 3552 47624
rect 3608 47568 3676 47624
rect 3732 47568 3800 47624
rect 3856 47568 3924 47624
rect 3980 47568 4048 47624
rect 4104 47568 4172 47624
rect 4228 47568 4296 47624
rect 4352 47568 4420 47624
rect 4476 47568 4544 47624
rect 4600 47568 4668 47624
rect 4724 47568 4791 47624
rect 2741 47500 4791 47568
rect 2741 47444 2808 47500
rect 2864 47444 2932 47500
rect 2988 47444 3056 47500
rect 3112 47444 3180 47500
rect 3236 47444 3304 47500
rect 3360 47444 3428 47500
rect 3484 47444 3552 47500
rect 3608 47444 3676 47500
rect 3732 47444 3800 47500
rect 3856 47444 3924 47500
rect 3980 47444 4048 47500
rect 4104 47444 4172 47500
rect 4228 47444 4296 47500
rect 4352 47444 4420 47500
rect 4476 47444 4544 47500
rect 4600 47444 4668 47500
rect 4724 47444 4791 47500
rect 2741 47376 4791 47444
rect 2741 47320 2808 47376
rect 2864 47320 2932 47376
rect 2988 47320 3056 47376
rect 3112 47320 3180 47376
rect 3236 47320 3304 47376
rect 3360 47320 3428 47376
rect 3484 47320 3552 47376
rect 3608 47320 3676 47376
rect 3732 47320 3800 47376
rect 3856 47320 3924 47376
rect 3980 47320 4048 47376
rect 4104 47320 4172 47376
rect 4228 47320 4296 47376
rect 4352 47320 4420 47376
rect 4476 47320 4544 47376
rect 4600 47320 4668 47376
rect 4724 47320 4791 47376
rect 2741 47281 4791 47320
rect 4851 57225 5051 57278
rect 4851 57169 4861 57225
rect 4917 57169 4985 57225
rect 5041 57169 5051 57225
rect 4851 57108 5051 57169
rect 4851 57101 4871 57108
rect 4851 57045 4861 57101
rect 4923 57056 4979 57108
rect 5031 57101 5051 57108
rect 4917 57045 4985 57056
rect 5041 57045 5051 57101
rect 4851 56977 5051 57045
rect 4851 56921 4861 56977
rect 4917 56921 4985 56977
rect 5041 56921 5051 56977
rect 4851 56853 5051 56921
rect 4851 56797 4861 56853
rect 4917 56797 4985 56853
rect 5041 56797 5051 56853
rect 4851 56729 5051 56797
rect 4851 56673 4861 56729
rect 4917 56673 4985 56729
rect 5041 56673 5051 56729
rect 4851 56605 5051 56673
rect 4851 56549 4861 56605
rect 4917 56549 4985 56605
rect 5041 56549 5051 56605
rect 4851 56481 5051 56549
rect 4851 56425 4861 56481
rect 4917 56425 4985 56481
rect 5041 56425 5051 56481
rect 4851 56357 5051 56425
rect 4851 56301 4861 56357
rect 4917 56301 4985 56357
rect 5041 56301 5051 56357
rect 4851 56233 5051 56301
rect 4851 56177 4861 56233
rect 4917 56177 4985 56233
rect 5041 56177 5051 56233
rect 4851 56109 5051 56177
rect 4851 56053 4861 56109
rect 4917 56053 4985 56109
rect 5041 56053 5051 56109
rect 4851 54148 5051 56053
rect 4851 54092 4861 54148
rect 4917 54092 4985 54148
rect 5041 54092 5051 54148
rect 4851 54024 5051 54092
rect 4851 53968 4861 54024
rect 4917 53968 4985 54024
rect 5041 53968 5051 54024
rect 4851 53900 5051 53968
rect 4851 53844 4861 53900
rect 4917 53844 4985 53900
rect 5041 53844 5051 53900
rect 4851 53776 5051 53844
rect 4851 53720 4861 53776
rect 4917 53720 4985 53776
rect 5041 53720 5051 53776
rect 4851 53652 5051 53720
rect 4851 53596 4861 53652
rect 4917 53596 4985 53652
rect 5041 53596 5051 53652
rect 4851 53528 5051 53596
rect 4851 53472 4861 53528
rect 4917 53484 4985 53528
rect 4851 53432 4871 53472
rect 4923 53432 4979 53484
rect 5041 53472 5051 53528
rect 5031 53432 5051 53472
rect 4851 53404 5051 53432
rect 4851 53348 4861 53404
rect 4917 53376 4985 53404
rect 4851 53324 4871 53348
rect 4923 53324 4979 53376
rect 5041 53348 5051 53404
rect 5031 53324 5051 53348
rect 4851 53280 5051 53324
rect 4851 53224 4861 53280
rect 4917 53268 4985 53280
rect 4851 53216 4871 53224
rect 4923 53216 4979 53268
rect 5041 53224 5051 53280
rect 5031 53216 5051 53224
rect 4851 53156 5051 53216
rect 4851 53100 4861 53156
rect 4917 53100 4985 53156
rect 5041 53100 5051 53156
rect 4851 53032 5051 53100
rect 4851 52976 4861 53032
rect 4917 52976 4985 53032
rect 5041 52976 5051 53032
rect 4851 52908 5051 52976
rect 4851 52852 4861 52908
rect 4917 52852 4985 52908
rect 5041 52852 5051 52908
rect 4851 52017 5051 52852
rect 4851 51965 4863 52017
rect 4915 51965 4987 52017
rect 5039 51965 5051 52017
rect 4851 51893 5051 51965
rect 4851 51841 4863 51893
rect 4915 51841 4987 51893
rect 5039 51841 5051 51893
rect 4851 51222 5051 51841
rect 4851 51170 4863 51222
rect 4915 51170 4987 51222
rect 5039 51170 5051 51222
rect 4851 51098 5051 51170
rect 4851 51046 4863 51098
rect 4915 51046 4987 51098
rect 5039 51046 5051 51098
rect 4851 50974 5051 51046
rect 4851 50922 4863 50974
rect 4915 50922 4987 50974
rect 5039 50922 5051 50974
rect 4851 50288 5051 50922
rect 4851 50236 4863 50288
rect 4915 50236 4987 50288
rect 5039 50236 5051 50288
rect 4851 50164 5051 50236
rect 4851 50112 4863 50164
rect 4915 50112 4987 50164
rect 5039 50112 5051 50164
rect 4851 50040 5051 50112
rect 4851 49988 4863 50040
rect 4915 49988 4987 50040
rect 5039 49988 5051 50040
rect 4851 49354 5051 49988
rect 4851 49348 4863 49354
rect 4915 49348 4987 49354
rect 5039 49348 5051 49354
rect 4851 49292 4861 49348
rect 4917 49292 4985 49348
rect 5041 49292 5051 49348
rect 4851 49230 5051 49292
rect 4851 49224 4863 49230
rect 4915 49224 4987 49230
rect 5039 49224 5051 49230
rect 4851 49168 4861 49224
rect 4917 49168 4985 49224
rect 5041 49168 5051 49224
rect 4851 49106 5051 49168
rect 4851 49100 4863 49106
rect 4915 49100 4987 49106
rect 5039 49100 5051 49106
rect 4851 49044 4861 49100
rect 4917 49044 4985 49100
rect 5041 49044 5051 49100
rect 4851 48976 5051 49044
rect 4851 48920 4861 48976
rect 4917 48920 4985 48976
rect 5041 48920 5051 48976
rect 4851 48852 5051 48920
rect 4851 48796 4861 48852
rect 4917 48796 4985 48852
rect 5041 48796 5051 48852
rect 4851 48728 5051 48796
rect 4851 48672 4861 48728
rect 4917 48672 4985 48728
rect 5041 48672 5051 48728
rect 4851 48604 5051 48672
rect 4851 48548 4861 48604
rect 4917 48548 4985 48604
rect 5041 48548 5051 48604
rect 4851 48480 5051 48548
rect 4851 48424 4861 48480
rect 4917 48424 4985 48480
rect 5041 48424 5051 48480
rect 4851 48383 4863 48424
rect 4915 48383 4987 48424
rect 5039 48383 5051 48424
rect 4851 48356 5051 48383
rect 4851 48300 4861 48356
rect 4917 48300 4985 48356
rect 5041 48300 5051 48356
rect 4851 48259 4863 48300
rect 4915 48259 4987 48300
rect 5039 48259 5051 48300
rect 4851 48232 5051 48259
rect 4851 48176 4861 48232
rect 4917 48176 4985 48232
rect 5041 48176 5051 48232
rect 4851 48108 5051 48176
rect 4851 48052 4861 48108
rect 4917 48052 4985 48108
rect 5041 48052 5051 48108
rect 4851 47281 5051 48052
rect 5111 56669 7161 57600
rect 5111 56617 6297 56669
rect 6349 56617 6421 56669
rect 6473 56617 6545 56669
rect 6597 56617 6669 56669
rect 6721 56617 6793 56669
rect 6845 56617 6917 56669
rect 6969 56617 7041 56669
rect 7093 56617 7161 56669
rect 5111 56545 7161 56617
rect 5111 56493 6297 56545
rect 6349 56493 6421 56545
rect 6473 56493 6545 56545
rect 6597 56493 6669 56545
rect 6721 56493 6793 56545
rect 6845 56493 6917 56545
rect 6969 56493 7041 56545
rect 7093 56493 7161 56545
rect 5111 56421 7161 56493
rect 5111 56369 6297 56421
rect 6349 56369 6421 56421
rect 6473 56369 6545 56421
rect 6597 56369 6669 56421
rect 6721 56369 6793 56421
rect 6845 56369 6917 56421
rect 6969 56369 7041 56421
rect 7093 56369 7161 56421
rect 5111 56297 7161 56369
rect 5111 56245 6297 56297
rect 6349 56245 6421 56297
rect 6473 56245 6545 56297
rect 6597 56245 6669 56297
rect 6721 56245 6793 56297
rect 6845 56245 6917 56297
rect 6969 56245 7041 56297
rect 7093 56245 7161 56297
rect 5111 56173 7161 56245
rect 5111 56121 6297 56173
rect 6349 56121 6421 56173
rect 6473 56121 6545 56173
rect 6597 56121 6669 56173
rect 6721 56121 6793 56173
rect 6845 56121 6917 56173
rect 6969 56121 7041 56173
rect 7093 56121 7161 56173
rect 5111 56049 7161 56121
rect 5111 55997 6297 56049
rect 6349 55997 6421 56049
rect 6473 55997 6545 56049
rect 6597 55997 6669 56049
rect 6721 55997 6793 56049
rect 6845 55997 6917 56049
rect 6969 55997 7041 56049
rect 7093 55997 7161 56049
rect 5111 55925 7161 55997
rect 5111 55873 6297 55925
rect 6349 55873 6421 55925
rect 6473 55873 6545 55925
rect 6597 55873 6669 55925
rect 6721 55873 6793 55925
rect 6845 55873 6917 55925
rect 6969 55873 7041 55925
rect 7093 55873 7161 55925
rect 5111 55801 7161 55873
rect 5111 55749 6297 55801
rect 6349 55749 6421 55801
rect 6473 55749 6545 55801
rect 6597 55749 6669 55801
rect 6721 55749 6793 55801
rect 6845 55749 6917 55801
rect 6969 55749 7041 55801
rect 7093 55749 7161 55801
rect 5111 55748 7161 55749
rect 5111 55692 5178 55748
rect 5234 55692 5302 55748
rect 5358 55692 5426 55748
rect 5482 55692 5550 55748
rect 5606 55692 5674 55748
rect 5730 55692 5798 55748
rect 5854 55692 5922 55748
rect 5978 55692 6046 55748
rect 6102 55692 6170 55748
rect 6226 55692 6294 55748
rect 6350 55692 6418 55748
rect 6474 55692 6542 55748
rect 6598 55692 6666 55748
rect 6722 55692 6790 55748
rect 6846 55692 6914 55748
rect 6970 55692 7038 55748
rect 7094 55692 7161 55748
rect 5111 55677 7161 55692
rect 5111 55625 6297 55677
rect 6349 55625 6421 55677
rect 6473 55625 6545 55677
rect 6597 55625 6669 55677
rect 6721 55625 6793 55677
rect 6845 55625 6917 55677
rect 6969 55625 7041 55677
rect 7093 55625 7161 55677
rect 5111 55624 7161 55625
rect 5111 55568 5178 55624
rect 5234 55568 5302 55624
rect 5358 55568 5426 55624
rect 5482 55568 5550 55624
rect 5606 55568 5674 55624
rect 5730 55568 5798 55624
rect 5854 55568 5922 55624
rect 5978 55568 6046 55624
rect 6102 55568 6170 55624
rect 6226 55568 6294 55624
rect 6350 55568 6418 55624
rect 6474 55568 6542 55624
rect 6598 55568 6666 55624
rect 6722 55568 6790 55624
rect 6846 55568 6914 55624
rect 6970 55568 7038 55624
rect 7094 55568 7161 55624
rect 5111 55553 7161 55568
rect 5111 55501 6297 55553
rect 6349 55501 6421 55553
rect 6473 55501 6545 55553
rect 6597 55501 6669 55553
rect 6721 55501 6793 55553
rect 6845 55501 6917 55553
rect 6969 55501 7041 55553
rect 7093 55501 7161 55553
rect 5111 55500 7161 55501
rect 5111 55444 5178 55500
rect 5234 55444 5302 55500
rect 5358 55444 5426 55500
rect 5482 55444 5550 55500
rect 5606 55444 5674 55500
rect 5730 55444 5798 55500
rect 5854 55444 5922 55500
rect 5978 55444 6046 55500
rect 6102 55444 6170 55500
rect 6226 55444 6294 55500
rect 6350 55444 6418 55500
rect 6474 55444 6542 55500
rect 6598 55444 6666 55500
rect 6722 55444 6790 55500
rect 6846 55444 6914 55500
rect 6970 55444 7038 55500
rect 7094 55444 7161 55500
rect 5111 55429 7161 55444
rect 5111 55377 6297 55429
rect 6349 55377 6421 55429
rect 6473 55377 6545 55429
rect 6597 55377 6669 55429
rect 6721 55377 6793 55429
rect 6845 55377 6917 55429
rect 6969 55377 7041 55429
rect 7093 55377 7161 55429
rect 5111 55376 7161 55377
rect 5111 55320 5178 55376
rect 5234 55320 5302 55376
rect 5358 55320 5426 55376
rect 5482 55320 5550 55376
rect 5606 55320 5674 55376
rect 5730 55320 5798 55376
rect 5854 55320 5922 55376
rect 5978 55320 6046 55376
rect 6102 55320 6170 55376
rect 6226 55320 6294 55376
rect 6350 55320 6418 55376
rect 6474 55320 6542 55376
rect 6598 55320 6666 55376
rect 6722 55320 6790 55376
rect 6846 55320 6914 55376
rect 6970 55320 7038 55376
rect 7094 55320 7161 55376
rect 5111 55305 7161 55320
rect 5111 55253 6297 55305
rect 6349 55253 6421 55305
rect 6473 55253 6545 55305
rect 6597 55253 6669 55305
rect 6721 55253 6793 55305
rect 6845 55253 6917 55305
rect 6969 55253 7041 55305
rect 7093 55253 7161 55305
rect 5111 55252 7161 55253
rect 5111 55196 5178 55252
rect 5234 55196 5302 55252
rect 5358 55196 5426 55252
rect 5482 55196 5550 55252
rect 5606 55196 5674 55252
rect 5730 55196 5798 55252
rect 5854 55196 5922 55252
rect 5978 55196 6046 55252
rect 6102 55196 6170 55252
rect 6226 55196 6294 55252
rect 6350 55196 6418 55252
rect 6474 55196 6542 55252
rect 6598 55196 6666 55252
rect 6722 55196 6790 55252
rect 6846 55196 6914 55252
rect 6970 55196 7038 55252
rect 7094 55196 7161 55252
rect 5111 55181 7161 55196
rect 5111 55129 6297 55181
rect 6349 55129 6421 55181
rect 6473 55129 6545 55181
rect 6597 55129 6669 55181
rect 6721 55129 6793 55181
rect 6845 55129 6917 55181
rect 6969 55129 7041 55181
rect 7093 55129 7161 55181
rect 5111 55128 7161 55129
rect 5111 55072 5178 55128
rect 5234 55072 5302 55128
rect 5358 55072 5426 55128
rect 5482 55072 5550 55128
rect 5606 55072 5674 55128
rect 5730 55072 5798 55128
rect 5854 55072 5922 55128
rect 5978 55072 6046 55128
rect 6102 55072 6170 55128
rect 6226 55072 6294 55128
rect 6350 55072 6418 55128
rect 6474 55072 6542 55128
rect 6598 55072 6666 55128
rect 6722 55072 6790 55128
rect 6846 55072 6914 55128
rect 6970 55072 7038 55128
rect 7094 55072 7161 55128
rect 5111 55057 7161 55072
rect 5111 55005 6297 55057
rect 6349 55005 6421 55057
rect 6473 55005 6545 55057
rect 6597 55005 6669 55057
rect 6721 55005 6793 55057
rect 6845 55005 6917 55057
rect 6969 55005 7041 55057
rect 7093 55005 7161 55057
rect 5111 55004 7161 55005
rect 5111 54948 5178 55004
rect 5234 54948 5302 55004
rect 5358 54948 5426 55004
rect 5482 54948 5550 55004
rect 5606 54948 5674 55004
rect 5730 54948 5798 55004
rect 5854 54948 5922 55004
rect 5978 54948 6046 55004
rect 6102 54948 6170 55004
rect 6226 54948 6294 55004
rect 6350 54948 6418 55004
rect 6474 54948 6542 55004
rect 6598 54948 6666 55004
rect 6722 54948 6790 55004
rect 6846 54948 6914 55004
rect 6970 54948 7038 55004
rect 7094 54948 7161 55004
rect 5111 54933 7161 54948
rect 5111 54881 6297 54933
rect 6349 54881 6421 54933
rect 6473 54881 6545 54933
rect 6597 54881 6669 54933
rect 6721 54881 6793 54933
rect 6845 54881 6917 54933
rect 6969 54881 7041 54933
rect 7093 54881 7161 54933
rect 5111 54880 7161 54881
rect 5111 54824 5178 54880
rect 5234 54824 5302 54880
rect 5358 54824 5426 54880
rect 5482 54824 5550 54880
rect 5606 54824 5674 54880
rect 5730 54824 5798 54880
rect 5854 54824 5922 54880
rect 5978 54824 6046 54880
rect 6102 54824 6170 54880
rect 6226 54824 6294 54880
rect 6350 54824 6418 54880
rect 6474 54824 6542 54880
rect 6598 54824 6666 54880
rect 6722 54824 6790 54880
rect 6846 54824 6914 54880
rect 6970 54824 7038 54880
rect 7094 54824 7161 54880
rect 5111 54809 7161 54824
rect 5111 54757 6297 54809
rect 6349 54757 6421 54809
rect 6473 54757 6545 54809
rect 6597 54757 6669 54809
rect 6721 54757 6793 54809
rect 6845 54757 6917 54809
rect 6969 54757 7041 54809
rect 7093 54757 7161 54809
rect 5111 54756 7161 54757
rect 5111 54700 5178 54756
rect 5234 54700 5302 54756
rect 5358 54700 5426 54756
rect 5482 54700 5550 54756
rect 5606 54700 5674 54756
rect 5730 54700 5798 54756
rect 5854 54700 5922 54756
rect 5978 54700 6046 54756
rect 6102 54700 6170 54756
rect 6226 54700 6294 54756
rect 6350 54700 6418 54756
rect 6474 54700 6542 54756
rect 6598 54700 6666 54756
rect 6722 54700 6790 54756
rect 6846 54700 6914 54756
rect 6970 54700 7038 54756
rect 7094 54700 7161 54756
rect 5111 54685 7161 54700
rect 5111 54633 6297 54685
rect 6349 54633 6421 54685
rect 6473 54633 6545 54685
rect 6597 54633 6669 54685
rect 6721 54633 6793 54685
rect 6845 54633 6917 54685
rect 6969 54633 7041 54685
rect 7093 54633 7161 54685
rect 5111 54632 7161 54633
rect 5111 54576 5178 54632
rect 5234 54576 5302 54632
rect 5358 54576 5426 54632
rect 5482 54576 5550 54632
rect 5606 54576 5674 54632
rect 5730 54576 5798 54632
rect 5854 54576 5922 54632
rect 5978 54576 6046 54632
rect 6102 54576 6170 54632
rect 6226 54576 6294 54632
rect 6350 54576 6418 54632
rect 6474 54576 6542 54632
rect 6598 54576 6666 54632
rect 6722 54576 6790 54632
rect 6846 54576 6914 54632
rect 6970 54576 7038 54632
rect 7094 54576 7161 54632
rect 5111 54561 7161 54576
rect 5111 54509 6297 54561
rect 6349 54509 6421 54561
rect 6473 54509 6545 54561
rect 6597 54509 6669 54561
rect 6721 54509 6793 54561
rect 6845 54509 6917 54561
rect 6969 54509 7041 54561
rect 7093 54509 7161 54561
rect 5111 54508 7161 54509
rect 5111 54452 5178 54508
rect 5234 54452 5302 54508
rect 5358 54452 5426 54508
rect 5482 54452 5550 54508
rect 5606 54452 5674 54508
rect 5730 54452 5798 54508
rect 5854 54452 5922 54508
rect 5978 54452 6046 54508
rect 6102 54452 6170 54508
rect 6226 54452 6294 54508
rect 6350 54452 6418 54508
rect 6474 54452 6542 54508
rect 6598 54452 6666 54508
rect 6722 54452 6790 54508
rect 6846 54452 6914 54508
rect 6970 54452 7038 54508
rect 7094 54452 7161 54508
rect 5111 54437 7161 54452
rect 5111 54385 6297 54437
rect 6349 54385 6421 54437
rect 6473 54385 6545 54437
rect 6597 54385 6669 54437
rect 6721 54385 6793 54437
rect 6845 54385 6917 54437
rect 6969 54385 7041 54437
rect 7093 54385 7161 54437
rect 5111 54313 7161 54385
rect 5111 54261 6297 54313
rect 6349 54261 6421 54313
rect 6473 54261 6545 54313
rect 6597 54261 6669 54313
rect 6721 54261 6793 54313
rect 6845 54261 6917 54313
rect 6969 54261 7041 54313
rect 7093 54261 7161 54313
rect 5111 54189 7161 54261
rect 5111 54137 6297 54189
rect 6349 54137 6421 54189
rect 6473 54137 6545 54189
rect 6597 54137 6669 54189
rect 6721 54137 6793 54189
rect 6845 54137 6917 54189
rect 6969 54137 7041 54189
rect 7093 54137 7161 54189
rect 5111 54065 7161 54137
rect 5111 54013 6297 54065
rect 6349 54013 6421 54065
rect 6473 54013 6545 54065
rect 6597 54013 6669 54065
rect 6721 54013 6793 54065
rect 6845 54013 6917 54065
rect 6969 54013 7041 54065
rect 7093 54013 7161 54065
rect 5111 53941 7161 54013
rect 5111 53889 6297 53941
rect 6349 53889 6421 53941
rect 6473 53889 6545 53941
rect 6597 53889 6669 53941
rect 6721 53889 6793 53941
rect 6845 53889 6917 53941
rect 6969 53889 7041 53941
rect 7093 53889 7161 53941
rect 5111 53817 7161 53889
rect 5111 53765 6297 53817
rect 6349 53765 6421 53817
rect 6473 53765 6545 53817
rect 6597 53765 6669 53817
rect 6721 53765 6793 53817
rect 6845 53765 6917 53817
rect 6969 53765 7041 53817
rect 7093 53765 7161 53817
rect 5111 53693 7161 53765
rect 5111 53641 6297 53693
rect 6349 53641 6421 53693
rect 6473 53641 6545 53693
rect 6597 53641 6669 53693
rect 6721 53641 6793 53693
rect 6845 53641 6917 53693
rect 6969 53641 7041 53693
rect 7093 53641 7161 53693
rect 5111 52588 7161 53641
rect 5111 52536 5180 52588
rect 5232 52536 5304 52588
rect 5356 52536 5428 52588
rect 5480 52536 5552 52588
rect 5604 52536 5676 52588
rect 5728 52536 5800 52588
rect 5852 52536 5924 52588
rect 5976 52536 6048 52588
rect 6100 52536 6172 52588
rect 6224 52536 6296 52588
rect 6348 52536 6420 52588
rect 6472 52536 6544 52588
rect 6596 52536 6668 52588
rect 6720 52536 6792 52588
rect 6844 52536 6916 52588
rect 6968 52536 7040 52588
rect 7092 52536 7161 52588
rect 5111 52464 7161 52536
rect 5111 52412 5180 52464
rect 5232 52412 5304 52464
rect 5356 52412 5428 52464
rect 5480 52412 5552 52464
rect 5604 52412 5676 52464
rect 5728 52412 5800 52464
rect 5852 52412 5924 52464
rect 5976 52412 6048 52464
rect 6100 52412 6172 52464
rect 6224 52412 6296 52464
rect 6348 52412 6420 52464
rect 6472 52412 6544 52464
rect 6596 52412 6668 52464
rect 6720 52412 6792 52464
rect 6844 52412 6916 52464
rect 6968 52412 7040 52464
rect 7092 52412 7161 52464
rect 5111 52340 7161 52412
rect 5111 52288 5180 52340
rect 5232 52288 5304 52340
rect 5356 52288 5428 52340
rect 5480 52288 5552 52340
rect 5604 52288 5676 52340
rect 5728 52288 5800 52340
rect 5852 52288 5924 52340
rect 5976 52288 6048 52340
rect 6100 52288 6172 52340
rect 6224 52288 6296 52340
rect 6348 52288 6420 52340
rect 6472 52288 6544 52340
rect 6596 52288 6668 52340
rect 6720 52288 6792 52340
rect 6844 52288 6916 52340
rect 6968 52288 7040 52340
rect 7092 52288 7161 52340
rect 5111 51627 7161 52288
rect 5111 51575 5180 51627
rect 5232 51575 5304 51627
rect 5356 51575 5428 51627
rect 5480 51575 5552 51627
rect 5604 51575 5676 51627
rect 5728 51575 5800 51627
rect 5852 51575 5924 51627
rect 5976 51575 6048 51627
rect 6100 51575 6172 51627
rect 6224 51575 6296 51627
rect 6348 51575 6420 51627
rect 6472 51575 6544 51627
rect 6596 51575 6668 51627
rect 6720 51575 6792 51627
rect 6844 51575 6916 51627
rect 6968 51575 7040 51627
rect 7092 51575 7161 51627
rect 5111 51503 7161 51575
rect 5111 51451 5180 51503
rect 5232 51451 5304 51503
rect 5356 51451 5428 51503
rect 5480 51451 5552 51503
rect 5604 51451 5676 51503
rect 5728 51451 5800 51503
rect 5852 51451 5924 51503
rect 5976 51451 6048 51503
rect 6100 51451 6172 51503
rect 6224 51451 6296 51503
rect 6348 51451 6420 51503
rect 6472 51451 6544 51503
rect 6596 51451 6668 51503
rect 6720 51451 6792 51503
rect 6844 51451 6916 51503
rect 6968 51451 7040 51503
rect 7092 51451 7161 51503
rect 5111 50948 7161 51451
rect 5111 50892 5178 50948
rect 5234 50892 5302 50948
rect 5358 50892 5426 50948
rect 5482 50892 5550 50948
rect 5606 50892 5674 50948
rect 5730 50892 5798 50948
rect 5854 50892 5922 50948
rect 5978 50892 6046 50948
rect 6102 50892 6170 50948
rect 6226 50892 6294 50948
rect 6350 50892 6418 50948
rect 6474 50892 6542 50948
rect 6598 50892 6666 50948
rect 6722 50892 6790 50948
rect 6846 50892 6914 50948
rect 6970 50892 7038 50948
rect 7094 50892 7161 50948
rect 5111 50824 7161 50892
rect 5111 50768 5178 50824
rect 5234 50768 5302 50824
rect 5358 50768 5426 50824
rect 5482 50768 5550 50824
rect 5606 50768 5674 50824
rect 5730 50768 5798 50824
rect 5854 50768 5922 50824
rect 5978 50768 6046 50824
rect 6102 50768 6170 50824
rect 6226 50768 6294 50824
rect 6350 50768 6418 50824
rect 6474 50768 6542 50824
rect 6598 50768 6666 50824
rect 6722 50768 6790 50824
rect 6846 50768 6914 50824
rect 6970 50768 7038 50824
rect 7094 50768 7161 50824
rect 5111 50700 7161 50768
rect 5111 50644 5178 50700
rect 5234 50644 5302 50700
rect 5358 50644 5426 50700
rect 5482 50644 5550 50700
rect 5606 50644 5674 50700
rect 5730 50644 5798 50700
rect 5854 50644 5922 50700
rect 5978 50644 6046 50700
rect 6102 50644 6170 50700
rect 6226 50644 6294 50700
rect 6350 50644 6418 50700
rect 6474 50644 6542 50700
rect 6598 50644 6666 50700
rect 6722 50644 6790 50700
rect 6846 50644 6914 50700
rect 6970 50644 7038 50700
rect 7094 50644 7161 50700
rect 5111 50641 5180 50644
rect 5232 50641 5304 50644
rect 5356 50641 5428 50644
rect 5480 50641 5552 50644
rect 5604 50641 5676 50644
rect 5728 50641 5800 50644
rect 5852 50641 5924 50644
rect 5976 50641 6048 50644
rect 6100 50641 6172 50644
rect 6224 50641 6296 50644
rect 6348 50641 6420 50644
rect 6472 50641 6544 50644
rect 6596 50641 6668 50644
rect 6720 50641 6792 50644
rect 6844 50641 6916 50644
rect 6968 50641 7040 50644
rect 7092 50641 7161 50644
rect 5111 50576 7161 50641
rect 5111 50520 5178 50576
rect 5234 50520 5302 50576
rect 5358 50520 5426 50576
rect 5482 50520 5550 50576
rect 5606 50520 5674 50576
rect 5730 50520 5798 50576
rect 5854 50520 5922 50576
rect 5978 50520 6046 50576
rect 6102 50520 6170 50576
rect 6226 50520 6294 50576
rect 6350 50520 6418 50576
rect 6474 50520 6542 50576
rect 6598 50520 6666 50576
rect 6722 50520 6790 50576
rect 6846 50520 6914 50576
rect 6970 50520 7038 50576
rect 7094 50520 7161 50576
rect 5111 50517 5180 50520
rect 5232 50517 5304 50520
rect 5356 50517 5428 50520
rect 5480 50517 5552 50520
rect 5604 50517 5676 50520
rect 5728 50517 5800 50520
rect 5852 50517 5924 50520
rect 5976 50517 6048 50520
rect 6100 50517 6172 50520
rect 6224 50517 6296 50520
rect 6348 50517 6420 50520
rect 6472 50517 6544 50520
rect 6596 50517 6668 50520
rect 6720 50517 6792 50520
rect 6844 50517 6916 50520
rect 6968 50517 7040 50520
rect 7092 50517 7161 50520
rect 5111 50452 7161 50517
rect 5111 50396 5178 50452
rect 5234 50396 5302 50452
rect 5358 50396 5426 50452
rect 5482 50396 5550 50452
rect 5606 50396 5674 50452
rect 5730 50396 5798 50452
rect 5854 50396 5922 50452
rect 5978 50396 6046 50452
rect 6102 50396 6170 50452
rect 6226 50396 6294 50452
rect 6350 50396 6418 50452
rect 6474 50396 6542 50452
rect 6598 50396 6666 50452
rect 6722 50396 6790 50452
rect 6846 50396 6914 50452
rect 6970 50396 7038 50452
rect 7094 50396 7161 50452
rect 5111 50328 7161 50396
rect 5111 50272 5178 50328
rect 5234 50272 5302 50328
rect 5358 50272 5426 50328
rect 5482 50272 5550 50328
rect 5606 50272 5674 50328
rect 5730 50272 5798 50328
rect 5854 50272 5922 50328
rect 5978 50272 6046 50328
rect 6102 50272 6170 50328
rect 6226 50272 6294 50328
rect 6350 50272 6418 50328
rect 6474 50272 6542 50328
rect 6598 50272 6666 50328
rect 6722 50272 6790 50328
rect 6846 50272 6914 50328
rect 6970 50272 7038 50328
rect 7094 50272 7161 50328
rect 5111 50204 7161 50272
rect 5111 50148 5178 50204
rect 5234 50148 5302 50204
rect 5358 50148 5426 50204
rect 5482 50148 5550 50204
rect 5606 50148 5674 50204
rect 5730 50148 5798 50204
rect 5854 50148 5922 50204
rect 5978 50148 6046 50204
rect 6102 50148 6170 50204
rect 6226 50148 6294 50204
rect 6350 50148 6418 50204
rect 6474 50148 6542 50204
rect 6598 50148 6666 50204
rect 6722 50148 6790 50204
rect 6846 50148 6914 50204
rect 6970 50148 7038 50204
rect 7094 50148 7161 50204
rect 5111 50080 7161 50148
rect 5111 50024 5178 50080
rect 5234 50024 5302 50080
rect 5358 50024 5426 50080
rect 5482 50024 5550 50080
rect 5606 50024 5674 50080
rect 5730 50024 5798 50080
rect 5854 50024 5922 50080
rect 5978 50024 6046 50080
rect 6102 50024 6170 50080
rect 6226 50024 6294 50080
rect 6350 50024 6418 50080
rect 6474 50024 6542 50080
rect 6598 50024 6666 50080
rect 6722 50024 6790 50080
rect 6846 50024 6914 50080
rect 6970 50024 7038 50080
rect 7094 50024 7161 50080
rect 5111 49956 7161 50024
rect 5111 49900 5178 49956
rect 5234 49900 5302 49956
rect 5358 49900 5426 49956
rect 5482 49900 5550 49956
rect 5606 49900 5674 49956
rect 5730 49900 5798 49956
rect 5854 49900 5922 49956
rect 5978 49900 6046 49956
rect 6102 49900 6170 49956
rect 6226 49900 6294 49956
rect 6350 49900 6418 49956
rect 6474 49900 6542 49956
rect 6598 49900 6666 49956
rect 6722 49900 6790 49956
rect 6846 49900 6914 49956
rect 6970 49900 7038 49956
rect 7094 49900 7161 49956
rect 5111 49832 7161 49900
rect 5111 49776 5178 49832
rect 5234 49776 5302 49832
rect 5358 49776 5426 49832
rect 5482 49776 5550 49832
rect 5606 49776 5674 49832
rect 5730 49776 5798 49832
rect 5854 49776 5922 49832
rect 5978 49776 6046 49832
rect 6102 49776 6170 49832
rect 6226 49776 6294 49832
rect 6350 49776 6418 49832
rect 6474 49776 6542 49832
rect 6598 49776 6666 49832
rect 6722 49776 6790 49832
rect 6846 49776 6914 49832
rect 6970 49776 7038 49832
rect 7094 49776 7161 49832
rect 5111 49759 7161 49776
rect 5111 49708 5180 49759
rect 5232 49708 5304 49759
rect 5356 49708 5428 49759
rect 5480 49708 5552 49759
rect 5604 49708 5676 49759
rect 5728 49708 5800 49759
rect 5852 49708 5924 49759
rect 5976 49708 6048 49759
rect 6100 49708 6172 49759
rect 6224 49708 6296 49759
rect 6348 49708 6420 49759
rect 6472 49708 6544 49759
rect 6596 49708 6668 49759
rect 6720 49708 6792 49759
rect 6844 49708 6916 49759
rect 6968 49708 7040 49759
rect 7092 49708 7161 49759
rect 5111 49652 5178 49708
rect 5234 49652 5302 49708
rect 5358 49652 5426 49708
rect 5482 49652 5550 49708
rect 5606 49652 5674 49708
rect 5730 49652 5798 49708
rect 5854 49652 5922 49708
rect 5978 49652 6046 49708
rect 6102 49652 6170 49708
rect 6226 49652 6294 49708
rect 6350 49652 6418 49708
rect 6474 49652 6542 49708
rect 6598 49652 6666 49708
rect 6722 49652 6790 49708
rect 6846 49652 6914 49708
rect 6970 49652 7038 49708
rect 7094 49652 7161 49708
rect 5111 49635 7161 49652
rect 5111 49583 5180 49635
rect 5232 49583 5304 49635
rect 5356 49583 5428 49635
rect 5480 49583 5552 49635
rect 5604 49583 5676 49635
rect 5728 49583 5800 49635
rect 5852 49583 5924 49635
rect 5976 49583 6048 49635
rect 6100 49583 6172 49635
rect 6224 49583 6296 49635
rect 6348 49583 6420 49635
rect 6472 49583 6544 49635
rect 6596 49583 6668 49635
rect 6720 49583 6792 49635
rect 6844 49583 6916 49635
rect 6968 49583 7040 49635
rect 7092 49583 7161 49635
rect 5111 48825 7161 49583
rect 5111 48773 5180 48825
rect 5232 48773 5304 48825
rect 5356 48773 5428 48825
rect 5480 48773 5552 48825
rect 5604 48773 5676 48825
rect 5728 48773 5800 48825
rect 5852 48773 5924 48825
rect 5976 48773 6048 48825
rect 6100 48773 6172 48825
rect 6224 48773 6296 48825
rect 6348 48773 6420 48825
rect 6472 48773 6544 48825
rect 6596 48773 6668 48825
rect 6720 48773 6792 48825
rect 6844 48773 6916 48825
rect 6968 48773 7040 48825
rect 7092 48773 7161 48825
rect 5111 48701 7161 48773
rect 5111 48649 5180 48701
rect 5232 48649 5304 48701
rect 5356 48649 5428 48701
rect 5480 48649 5552 48701
rect 5604 48649 5676 48701
rect 5728 48649 5800 48701
rect 5852 48649 5924 48701
rect 5976 48649 6048 48701
rect 6100 48649 6172 48701
rect 6224 48649 6296 48701
rect 6348 48649 6420 48701
rect 6472 48649 6544 48701
rect 6596 48649 6668 48701
rect 6720 48649 6792 48701
rect 6844 48649 6916 48701
rect 6968 48649 7040 48701
rect 7092 48649 7161 48701
rect 5111 47988 7161 48649
rect 5111 47936 5180 47988
rect 5232 47936 5304 47988
rect 5356 47936 5428 47988
rect 5480 47936 5552 47988
rect 5604 47936 5676 47988
rect 5728 47936 5800 47988
rect 5852 47936 5924 47988
rect 5976 47936 6048 47988
rect 6100 47936 6172 47988
rect 6224 47936 6296 47988
rect 6348 47936 6420 47988
rect 6472 47936 6544 47988
rect 6596 47936 6668 47988
rect 6720 47936 6792 47988
rect 6844 47936 6916 47988
rect 6968 47936 7040 47988
rect 7092 47936 7161 47988
rect 5111 47864 7161 47936
rect 5111 47812 5180 47864
rect 5232 47812 5304 47864
rect 5356 47812 5428 47864
rect 5480 47812 5552 47864
rect 5604 47812 5676 47864
rect 5728 47812 5800 47864
rect 5852 47812 5924 47864
rect 5976 47812 6048 47864
rect 6100 47812 6172 47864
rect 6224 47812 6296 47864
rect 6348 47812 6420 47864
rect 6472 47812 6544 47864
rect 6596 47812 6668 47864
rect 6720 47812 6792 47864
rect 6844 47812 6916 47864
rect 6968 47812 7040 47864
rect 7092 47812 7161 47864
rect 5111 47748 7161 47812
rect 5111 47692 5178 47748
rect 5234 47692 5302 47748
rect 5358 47692 5426 47748
rect 5482 47692 5550 47748
rect 5606 47692 5674 47748
rect 5730 47692 5798 47748
rect 5854 47692 5922 47748
rect 5978 47692 6046 47748
rect 6102 47692 6170 47748
rect 6226 47692 6294 47748
rect 6350 47692 6418 47748
rect 6474 47692 6542 47748
rect 6598 47692 6666 47748
rect 6722 47692 6790 47748
rect 6846 47692 6914 47748
rect 6970 47692 7038 47748
rect 7094 47692 7161 47748
rect 5111 47688 5180 47692
rect 5232 47688 5304 47692
rect 5356 47688 5428 47692
rect 5480 47688 5552 47692
rect 5604 47688 5676 47692
rect 5728 47688 5800 47692
rect 5852 47688 5924 47692
rect 5976 47688 6048 47692
rect 6100 47688 6172 47692
rect 6224 47688 6296 47692
rect 6348 47688 6420 47692
rect 6472 47688 6544 47692
rect 6596 47688 6668 47692
rect 6720 47688 6792 47692
rect 6844 47688 6916 47692
rect 6968 47688 7040 47692
rect 7092 47688 7161 47692
rect 5111 47624 7161 47688
rect 5111 47568 5178 47624
rect 5234 47568 5302 47624
rect 5358 47568 5426 47624
rect 5482 47568 5550 47624
rect 5606 47568 5674 47624
rect 5730 47568 5798 47624
rect 5854 47568 5922 47624
rect 5978 47568 6046 47624
rect 6102 47568 6170 47624
rect 6226 47568 6294 47624
rect 6350 47568 6418 47624
rect 6474 47568 6542 47624
rect 6598 47568 6666 47624
rect 6722 47568 6790 47624
rect 6846 47568 6914 47624
rect 6970 47568 7038 47624
rect 7094 47568 7161 47624
rect 5111 47500 7161 47568
rect 5111 47444 5178 47500
rect 5234 47444 5302 47500
rect 5358 47444 5426 47500
rect 5482 47444 5550 47500
rect 5606 47444 5674 47500
rect 5730 47444 5798 47500
rect 5854 47444 5922 47500
rect 5978 47444 6046 47500
rect 6102 47444 6170 47500
rect 6226 47444 6294 47500
rect 6350 47444 6418 47500
rect 6474 47444 6542 47500
rect 6598 47444 6666 47500
rect 6722 47444 6790 47500
rect 6846 47444 6914 47500
rect 6970 47444 7038 47500
rect 7094 47444 7161 47500
rect 5111 47376 7161 47444
rect 5111 47320 5178 47376
rect 5234 47320 5302 47376
rect 5358 47320 5426 47376
rect 5482 47320 5550 47376
rect 5606 47320 5674 47376
rect 5730 47320 5798 47376
rect 5854 47320 5922 47376
rect 5978 47320 6046 47376
rect 6102 47320 6170 47376
rect 6226 47320 6294 47376
rect 6350 47320 6418 47376
rect 6474 47320 6542 47376
rect 6598 47320 6666 47376
rect 6722 47320 6790 47376
rect 6846 47320 6914 47376
rect 6970 47320 7038 47376
rect 7094 47320 7161 47376
rect 5111 47281 7161 47320
rect 7221 57225 7757 57278
rect 7221 57169 7275 57225
rect 7331 57169 7399 57225
rect 7455 57169 7523 57225
rect 7579 57169 7647 57225
rect 7703 57169 7757 57225
rect 7221 57108 7757 57169
rect 7221 57056 7247 57108
rect 7299 57101 7355 57108
rect 7407 57101 7463 57108
rect 7331 57056 7355 57101
rect 7455 57056 7463 57101
rect 7515 57101 7571 57108
rect 7623 57101 7679 57108
rect 7515 57056 7523 57101
rect 7623 57056 7647 57101
rect 7731 57056 7757 57108
rect 7221 57045 7275 57056
rect 7331 57045 7399 57056
rect 7455 57045 7523 57056
rect 7579 57045 7647 57056
rect 7703 57045 7757 57056
rect 7221 56977 7757 57045
rect 7221 56921 7275 56977
rect 7331 56921 7399 56977
rect 7455 56921 7523 56977
rect 7579 56921 7647 56977
rect 7703 56921 7757 56977
rect 7221 56853 7757 56921
rect 7221 56797 7275 56853
rect 7331 56797 7399 56853
rect 7455 56797 7523 56853
rect 7579 56797 7647 56853
rect 7703 56797 7757 56853
rect 7221 56729 7757 56797
rect 7221 56673 7275 56729
rect 7331 56673 7399 56729
rect 7455 56673 7523 56729
rect 7579 56673 7647 56729
rect 7703 56673 7757 56729
rect 7221 56605 7757 56673
rect 7221 56549 7275 56605
rect 7331 56549 7399 56605
rect 7455 56549 7523 56605
rect 7579 56549 7647 56605
rect 7703 56549 7757 56605
rect 7221 56481 7757 56549
rect 7221 56425 7275 56481
rect 7331 56425 7399 56481
rect 7455 56425 7523 56481
rect 7579 56425 7647 56481
rect 7703 56425 7757 56481
rect 7221 56357 7757 56425
rect 7221 56301 7275 56357
rect 7331 56301 7399 56357
rect 7455 56301 7523 56357
rect 7579 56301 7647 56357
rect 7703 56301 7757 56357
rect 7221 56233 7757 56301
rect 7221 56177 7275 56233
rect 7331 56177 7399 56233
rect 7455 56177 7523 56233
rect 7579 56177 7647 56233
rect 7703 56177 7757 56233
rect 7221 56109 7757 56177
rect 7221 56053 7275 56109
rect 7331 56053 7399 56109
rect 7455 56053 7523 56109
rect 7579 56053 7647 56109
rect 7703 56053 7757 56109
rect 7221 54148 7757 56053
rect 7221 54092 7275 54148
rect 7331 54092 7399 54148
rect 7455 54092 7523 54148
rect 7579 54092 7647 54148
rect 7703 54092 7757 54148
rect 7221 54024 7757 54092
rect 7221 53968 7275 54024
rect 7331 53968 7399 54024
rect 7455 53968 7523 54024
rect 7579 53968 7647 54024
rect 7703 53968 7757 54024
rect 7221 53900 7757 53968
rect 7221 53844 7275 53900
rect 7331 53844 7399 53900
rect 7455 53844 7523 53900
rect 7579 53844 7647 53900
rect 7703 53844 7757 53900
rect 7221 53776 7757 53844
rect 7221 53720 7275 53776
rect 7331 53720 7399 53776
rect 7455 53720 7523 53776
rect 7579 53720 7647 53776
rect 7703 53720 7757 53776
rect 7221 53652 7757 53720
rect 7221 53596 7275 53652
rect 7331 53596 7399 53652
rect 7455 53596 7523 53652
rect 7579 53596 7647 53652
rect 7703 53596 7757 53652
rect 7221 53528 7757 53596
rect 7221 53484 7275 53528
rect 7331 53484 7399 53528
rect 7455 53484 7523 53528
rect 7579 53484 7647 53528
rect 7703 53484 7757 53528
rect 7221 53432 7247 53484
rect 7331 53472 7355 53484
rect 7455 53472 7463 53484
rect 7299 53432 7355 53472
rect 7407 53432 7463 53472
rect 7515 53472 7523 53484
rect 7623 53472 7647 53484
rect 7515 53432 7571 53472
rect 7623 53432 7679 53472
rect 7731 53432 7757 53484
rect 7221 53404 7757 53432
rect 7221 53376 7275 53404
rect 7331 53376 7399 53404
rect 7455 53376 7523 53404
rect 7579 53376 7647 53404
rect 7703 53376 7757 53404
rect 7221 53324 7247 53376
rect 7331 53348 7355 53376
rect 7455 53348 7463 53376
rect 7299 53324 7355 53348
rect 7407 53324 7463 53348
rect 7515 53348 7523 53376
rect 7623 53348 7647 53376
rect 7515 53324 7571 53348
rect 7623 53324 7679 53348
rect 7731 53324 7757 53376
rect 7221 53280 7757 53324
rect 7221 53268 7275 53280
rect 7331 53268 7399 53280
rect 7455 53268 7523 53280
rect 7579 53268 7647 53280
rect 7703 53268 7757 53280
rect 7221 53216 7247 53268
rect 7331 53224 7355 53268
rect 7455 53224 7463 53268
rect 7299 53216 7355 53224
rect 7407 53216 7463 53224
rect 7515 53224 7523 53268
rect 7623 53224 7647 53268
rect 7515 53216 7571 53224
rect 7623 53216 7679 53224
rect 7731 53216 7757 53268
rect 7221 53156 7757 53216
rect 7221 53100 7275 53156
rect 7331 53100 7399 53156
rect 7455 53100 7523 53156
rect 7579 53100 7647 53156
rect 7703 53100 7757 53156
rect 7221 53032 7757 53100
rect 7221 52976 7275 53032
rect 7331 52976 7399 53032
rect 7455 52976 7523 53032
rect 7579 52976 7647 53032
rect 7703 52976 7757 53032
rect 7221 52908 7757 52976
rect 7221 52852 7275 52908
rect 7331 52852 7399 52908
rect 7455 52852 7523 52908
rect 7579 52852 7647 52908
rect 7703 52852 7757 52908
rect 7221 52017 7757 52852
rect 7221 51965 7277 52017
rect 7329 51965 7401 52017
rect 7453 51965 7525 52017
rect 7577 51965 7649 52017
rect 7701 51965 7757 52017
rect 7221 51893 7757 51965
rect 7221 51841 7277 51893
rect 7329 51841 7401 51893
rect 7453 51841 7525 51893
rect 7577 51841 7649 51893
rect 7701 51841 7757 51893
rect 7221 51222 7757 51841
rect 7221 51170 7277 51222
rect 7329 51170 7401 51222
rect 7453 51170 7525 51222
rect 7577 51170 7649 51222
rect 7701 51170 7757 51222
rect 7221 51098 7757 51170
rect 7221 51046 7277 51098
rect 7329 51046 7401 51098
rect 7453 51046 7525 51098
rect 7577 51046 7649 51098
rect 7701 51046 7757 51098
rect 7221 50974 7757 51046
rect 7221 50922 7277 50974
rect 7329 50922 7401 50974
rect 7453 50922 7525 50974
rect 7577 50922 7649 50974
rect 7701 50922 7757 50974
rect 7221 50288 7757 50922
rect 7221 50236 7277 50288
rect 7329 50236 7401 50288
rect 7453 50236 7525 50288
rect 7577 50236 7649 50288
rect 7701 50236 7757 50288
rect 7221 50164 7757 50236
rect 7221 50112 7277 50164
rect 7329 50112 7401 50164
rect 7453 50112 7525 50164
rect 7577 50112 7649 50164
rect 7701 50112 7757 50164
rect 7221 50040 7757 50112
rect 7221 49988 7277 50040
rect 7329 49988 7401 50040
rect 7453 49988 7525 50040
rect 7577 49988 7649 50040
rect 7701 49988 7757 50040
rect 7221 49354 7757 49988
rect 7221 49348 7277 49354
rect 7329 49348 7401 49354
rect 7453 49348 7525 49354
rect 7577 49348 7649 49354
rect 7701 49348 7757 49354
rect 7221 49292 7275 49348
rect 7331 49292 7399 49348
rect 7455 49292 7523 49348
rect 7579 49292 7647 49348
rect 7703 49292 7757 49348
rect 7221 49230 7757 49292
rect 7221 49224 7277 49230
rect 7329 49224 7401 49230
rect 7453 49224 7525 49230
rect 7577 49224 7649 49230
rect 7701 49224 7757 49230
rect 7221 49168 7275 49224
rect 7331 49168 7399 49224
rect 7455 49168 7523 49224
rect 7579 49168 7647 49224
rect 7703 49168 7757 49224
rect 7221 49106 7757 49168
rect 7221 49100 7277 49106
rect 7329 49100 7401 49106
rect 7453 49100 7525 49106
rect 7577 49100 7649 49106
rect 7701 49100 7757 49106
rect 7221 49044 7275 49100
rect 7331 49044 7399 49100
rect 7455 49044 7523 49100
rect 7579 49044 7647 49100
rect 7703 49044 7757 49100
rect 7221 48976 7757 49044
rect 7221 48920 7275 48976
rect 7331 48920 7399 48976
rect 7455 48920 7523 48976
rect 7579 48920 7647 48976
rect 7703 48920 7757 48976
rect 7221 48852 7757 48920
rect 7221 48796 7275 48852
rect 7331 48796 7399 48852
rect 7455 48796 7523 48852
rect 7579 48796 7647 48852
rect 7703 48796 7757 48852
rect 7221 48728 7757 48796
rect 7221 48672 7275 48728
rect 7331 48672 7399 48728
rect 7455 48672 7523 48728
rect 7579 48672 7647 48728
rect 7703 48672 7757 48728
rect 7221 48604 7757 48672
rect 7221 48548 7275 48604
rect 7331 48548 7399 48604
rect 7455 48548 7523 48604
rect 7579 48548 7647 48604
rect 7703 48548 7757 48604
rect 7221 48480 7757 48548
rect 7221 48424 7275 48480
rect 7331 48424 7399 48480
rect 7455 48424 7523 48480
rect 7579 48424 7647 48480
rect 7703 48424 7757 48480
rect 7221 48383 7277 48424
rect 7329 48383 7401 48424
rect 7453 48383 7525 48424
rect 7577 48383 7649 48424
rect 7701 48383 7757 48424
rect 7221 48356 7757 48383
rect 7221 48300 7275 48356
rect 7331 48300 7399 48356
rect 7455 48300 7523 48356
rect 7579 48300 7647 48356
rect 7703 48300 7757 48356
rect 7221 48259 7277 48300
rect 7329 48259 7401 48300
rect 7453 48259 7525 48300
rect 7577 48259 7649 48300
rect 7701 48259 7757 48300
rect 7221 48232 7757 48259
rect 7221 48176 7275 48232
rect 7331 48176 7399 48232
rect 7455 48176 7523 48232
rect 7579 48176 7647 48232
rect 7703 48176 7757 48232
rect 7221 48108 7757 48176
rect 7221 48052 7275 48108
rect 7331 48052 7399 48108
rect 7455 48052 7523 48108
rect 7579 48052 7647 48108
rect 7703 48052 7757 48108
rect 7221 47281 7757 48052
rect 7817 56669 9867 57600
rect 7817 56617 7885 56669
rect 7937 56617 8009 56669
rect 8061 56617 8133 56669
rect 8185 56617 8257 56669
rect 8309 56617 8381 56669
rect 8433 56617 8505 56669
rect 8557 56617 8629 56669
rect 8681 56617 9867 56669
rect 7817 56545 9867 56617
rect 7817 56493 7885 56545
rect 7937 56493 8009 56545
rect 8061 56493 8133 56545
rect 8185 56493 8257 56545
rect 8309 56493 8381 56545
rect 8433 56493 8505 56545
rect 8557 56493 8629 56545
rect 8681 56493 9867 56545
rect 7817 56421 9867 56493
rect 7817 56369 7885 56421
rect 7937 56369 8009 56421
rect 8061 56369 8133 56421
rect 8185 56369 8257 56421
rect 8309 56369 8381 56421
rect 8433 56369 8505 56421
rect 8557 56369 8629 56421
rect 8681 56369 9867 56421
rect 7817 56297 9867 56369
rect 7817 56245 7885 56297
rect 7937 56245 8009 56297
rect 8061 56245 8133 56297
rect 8185 56245 8257 56297
rect 8309 56245 8381 56297
rect 8433 56245 8505 56297
rect 8557 56245 8629 56297
rect 8681 56245 9867 56297
rect 7817 56173 9867 56245
rect 7817 56121 7885 56173
rect 7937 56121 8009 56173
rect 8061 56121 8133 56173
rect 8185 56121 8257 56173
rect 8309 56121 8381 56173
rect 8433 56121 8505 56173
rect 8557 56121 8629 56173
rect 8681 56121 9867 56173
rect 7817 56049 9867 56121
rect 7817 55997 7885 56049
rect 7937 55997 8009 56049
rect 8061 55997 8133 56049
rect 8185 55997 8257 56049
rect 8309 55997 8381 56049
rect 8433 55997 8505 56049
rect 8557 55997 8629 56049
rect 8681 55997 9867 56049
rect 7817 55925 9867 55997
rect 7817 55873 7885 55925
rect 7937 55873 8009 55925
rect 8061 55873 8133 55925
rect 8185 55873 8257 55925
rect 8309 55873 8381 55925
rect 8433 55873 8505 55925
rect 8557 55873 8629 55925
rect 8681 55873 9867 55925
rect 7817 55801 9867 55873
rect 7817 55749 7885 55801
rect 7937 55749 8009 55801
rect 8061 55749 8133 55801
rect 8185 55749 8257 55801
rect 8309 55749 8381 55801
rect 8433 55749 8505 55801
rect 8557 55749 8629 55801
rect 8681 55749 9867 55801
rect 7817 55748 9867 55749
rect 7817 55692 7884 55748
rect 7940 55692 8008 55748
rect 8064 55692 8132 55748
rect 8188 55692 8256 55748
rect 8312 55692 8380 55748
rect 8436 55692 8504 55748
rect 8560 55692 8628 55748
rect 8684 55692 8752 55748
rect 8808 55692 8876 55748
rect 8932 55692 9000 55748
rect 9056 55692 9124 55748
rect 9180 55692 9248 55748
rect 9304 55692 9372 55748
rect 9428 55692 9496 55748
rect 9552 55692 9620 55748
rect 9676 55692 9744 55748
rect 9800 55692 9867 55748
rect 7817 55677 9867 55692
rect 7817 55625 7885 55677
rect 7937 55625 8009 55677
rect 8061 55625 8133 55677
rect 8185 55625 8257 55677
rect 8309 55625 8381 55677
rect 8433 55625 8505 55677
rect 8557 55625 8629 55677
rect 8681 55625 9867 55677
rect 7817 55624 9867 55625
rect 7817 55568 7884 55624
rect 7940 55568 8008 55624
rect 8064 55568 8132 55624
rect 8188 55568 8256 55624
rect 8312 55568 8380 55624
rect 8436 55568 8504 55624
rect 8560 55568 8628 55624
rect 8684 55568 8752 55624
rect 8808 55568 8876 55624
rect 8932 55568 9000 55624
rect 9056 55568 9124 55624
rect 9180 55568 9248 55624
rect 9304 55568 9372 55624
rect 9428 55568 9496 55624
rect 9552 55568 9620 55624
rect 9676 55568 9744 55624
rect 9800 55568 9867 55624
rect 7817 55553 9867 55568
rect 7817 55501 7885 55553
rect 7937 55501 8009 55553
rect 8061 55501 8133 55553
rect 8185 55501 8257 55553
rect 8309 55501 8381 55553
rect 8433 55501 8505 55553
rect 8557 55501 8629 55553
rect 8681 55501 9867 55553
rect 7817 55500 9867 55501
rect 7817 55444 7884 55500
rect 7940 55444 8008 55500
rect 8064 55444 8132 55500
rect 8188 55444 8256 55500
rect 8312 55444 8380 55500
rect 8436 55444 8504 55500
rect 8560 55444 8628 55500
rect 8684 55444 8752 55500
rect 8808 55444 8876 55500
rect 8932 55444 9000 55500
rect 9056 55444 9124 55500
rect 9180 55444 9248 55500
rect 9304 55444 9372 55500
rect 9428 55444 9496 55500
rect 9552 55444 9620 55500
rect 9676 55444 9744 55500
rect 9800 55444 9867 55500
rect 7817 55429 9867 55444
rect 7817 55377 7885 55429
rect 7937 55377 8009 55429
rect 8061 55377 8133 55429
rect 8185 55377 8257 55429
rect 8309 55377 8381 55429
rect 8433 55377 8505 55429
rect 8557 55377 8629 55429
rect 8681 55377 9867 55429
rect 7817 55376 9867 55377
rect 7817 55320 7884 55376
rect 7940 55320 8008 55376
rect 8064 55320 8132 55376
rect 8188 55320 8256 55376
rect 8312 55320 8380 55376
rect 8436 55320 8504 55376
rect 8560 55320 8628 55376
rect 8684 55320 8752 55376
rect 8808 55320 8876 55376
rect 8932 55320 9000 55376
rect 9056 55320 9124 55376
rect 9180 55320 9248 55376
rect 9304 55320 9372 55376
rect 9428 55320 9496 55376
rect 9552 55320 9620 55376
rect 9676 55320 9744 55376
rect 9800 55320 9867 55376
rect 7817 55305 9867 55320
rect 7817 55253 7885 55305
rect 7937 55253 8009 55305
rect 8061 55253 8133 55305
rect 8185 55253 8257 55305
rect 8309 55253 8381 55305
rect 8433 55253 8505 55305
rect 8557 55253 8629 55305
rect 8681 55253 9867 55305
rect 7817 55252 9867 55253
rect 7817 55196 7884 55252
rect 7940 55196 8008 55252
rect 8064 55196 8132 55252
rect 8188 55196 8256 55252
rect 8312 55196 8380 55252
rect 8436 55196 8504 55252
rect 8560 55196 8628 55252
rect 8684 55196 8752 55252
rect 8808 55196 8876 55252
rect 8932 55196 9000 55252
rect 9056 55196 9124 55252
rect 9180 55196 9248 55252
rect 9304 55196 9372 55252
rect 9428 55196 9496 55252
rect 9552 55196 9620 55252
rect 9676 55196 9744 55252
rect 9800 55196 9867 55252
rect 7817 55181 9867 55196
rect 7817 55129 7885 55181
rect 7937 55129 8009 55181
rect 8061 55129 8133 55181
rect 8185 55129 8257 55181
rect 8309 55129 8381 55181
rect 8433 55129 8505 55181
rect 8557 55129 8629 55181
rect 8681 55129 9867 55181
rect 7817 55128 9867 55129
rect 7817 55072 7884 55128
rect 7940 55072 8008 55128
rect 8064 55072 8132 55128
rect 8188 55072 8256 55128
rect 8312 55072 8380 55128
rect 8436 55072 8504 55128
rect 8560 55072 8628 55128
rect 8684 55072 8752 55128
rect 8808 55072 8876 55128
rect 8932 55072 9000 55128
rect 9056 55072 9124 55128
rect 9180 55072 9248 55128
rect 9304 55072 9372 55128
rect 9428 55072 9496 55128
rect 9552 55072 9620 55128
rect 9676 55072 9744 55128
rect 9800 55072 9867 55128
rect 7817 55057 9867 55072
rect 7817 55005 7885 55057
rect 7937 55005 8009 55057
rect 8061 55005 8133 55057
rect 8185 55005 8257 55057
rect 8309 55005 8381 55057
rect 8433 55005 8505 55057
rect 8557 55005 8629 55057
rect 8681 55005 9867 55057
rect 7817 55004 9867 55005
rect 7817 54948 7884 55004
rect 7940 54948 8008 55004
rect 8064 54948 8132 55004
rect 8188 54948 8256 55004
rect 8312 54948 8380 55004
rect 8436 54948 8504 55004
rect 8560 54948 8628 55004
rect 8684 54948 8752 55004
rect 8808 54948 8876 55004
rect 8932 54948 9000 55004
rect 9056 54948 9124 55004
rect 9180 54948 9248 55004
rect 9304 54948 9372 55004
rect 9428 54948 9496 55004
rect 9552 54948 9620 55004
rect 9676 54948 9744 55004
rect 9800 54948 9867 55004
rect 7817 54933 9867 54948
rect 7817 54881 7885 54933
rect 7937 54881 8009 54933
rect 8061 54881 8133 54933
rect 8185 54881 8257 54933
rect 8309 54881 8381 54933
rect 8433 54881 8505 54933
rect 8557 54881 8629 54933
rect 8681 54881 9867 54933
rect 7817 54880 9867 54881
rect 7817 54824 7884 54880
rect 7940 54824 8008 54880
rect 8064 54824 8132 54880
rect 8188 54824 8256 54880
rect 8312 54824 8380 54880
rect 8436 54824 8504 54880
rect 8560 54824 8628 54880
rect 8684 54824 8752 54880
rect 8808 54824 8876 54880
rect 8932 54824 9000 54880
rect 9056 54824 9124 54880
rect 9180 54824 9248 54880
rect 9304 54824 9372 54880
rect 9428 54824 9496 54880
rect 9552 54824 9620 54880
rect 9676 54824 9744 54880
rect 9800 54824 9867 54880
rect 7817 54809 9867 54824
rect 7817 54757 7885 54809
rect 7937 54757 8009 54809
rect 8061 54757 8133 54809
rect 8185 54757 8257 54809
rect 8309 54757 8381 54809
rect 8433 54757 8505 54809
rect 8557 54757 8629 54809
rect 8681 54757 9867 54809
rect 7817 54756 9867 54757
rect 7817 54700 7884 54756
rect 7940 54700 8008 54756
rect 8064 54700 8132 54756
rect 8188 54700 8256 54756
rect 8312 54700 8380 54756
rect 8436 54700 8504 54756
rect 8560 54700 8628 54756
rect 8684 54700 8752 54756
rect 8808 54700 8876 54756
rect 8932 54700 9000 54756
rect 9056 54700 9124 54756
rect 9180 54700 9248 54756
rect 9304 54700 9372 54756
rect 9428 54700 9496 54756
rect 9552 54700 9620 54756
rect 9676 54700 9744 54756
rect 9800 54700 9867 54756
rect 7817 54685 9867 54700
rect 7817 54633 7885 54685
rect 7937 54633 8009 54685
rect 8061 54633 8133 54685
rect 8185 54633 8257 54685
rect 8309 54633 8381 54685
rect 8433 54633 8505 54685
rect 8557 54633 8629 54685
rect 8681 54633 9867 54685
rect 7817 54632 9867 54633
rect 7817 54576 7884 54632
rect 7940 54576 8008 54632
rect 8064 54576 8132 54632
rect 8188 54576 8256 54632
rect 8312 54576 8380 54632
rect 8436 54576 8504 54632
rect 8560 54576 8628 54632
rect 8684 54576 8752 54632
rect 8808 54576 8876 54632
rect 8932 54576 9000 54632
rect 9056 54576 9124 54632
rect 9180 54576 9248 54632
rect 9304 54576 9372 54632
rect 9428 54576 9496 54632
rect 9552 54576 9620 54632
rect 9676 54576 9744 54632
rect 9800 54576 9867 54632
rect 7817 54561 9867 54576
rect 7817 54509 7885 54561
rect 7937 54509 8009 54561
rect 8061 54509 8133 54561
rect 8185 54509 8257 54561
rect 8309 54509 8381 54561
rect 8433 54509 8505 54561
rect 8557 54509 8629 54561
rect 8681 54509 9867 54561
rect 7817 54508 9867 54509
rect 7817 54452 7884 54508
rect 7940 54452 8008 54508
rect 8064 54452 8132 54508
rect 8188 54452 8256 54508
rect 8312 54452 8380 54508
rect 8436 54452 8504 54508
rect 8560 54452 8628 54508
rect 8684 54452 8752 54508
rect 8808 54452 8876 54508
rect 8932 54452 9000 54508
rect 9056 54452 9124 54508
rect 9180 54452 9248 54508
rect 9304 54452 9372 54508
rect 9428 54452 9496 54508
rect 9552 54452 9620 54508
rect 9676 54452 9744 54508
rect 9800 54452 9867 54508
rect 7817 54437 9867 54452
rect 7817 54385 7885 54437
rect 7937 54385 8009 54437
rect 8061 54385 8133 54437
rect 8185 54385 8257 54437
rect 8309 54385 8381 54437
rect 8433 54385 8505 54437
rect 8557 54385 8629 54437
rect 8681 54385 9867 54437
rect 7817 54313 9867 54385
rect 7817 54261 7885 54313
rect 7937 54261 8009 54313
rect 8061 54261 8133 54313
rect 8185 54261 8257 54313
rect 8309 54261 8381 54313
rect 8433 54261 8505 54313
rect 8557 54261 8629 54313
rect 8681 54261 9867 54313
rect 7817 54189 9867 54261
rect 7817 54137 7885 54189
rect 7937 54137 8009 54189
rect 8061 54137 8133 54189
rect 8185 54137 8257 54189
rect 8309 54137 8381 54189
rect 8433 54137 8505 54189
rect 8557 54137 8629 54189
rect 8681 54137 9867 54189
rect 7817 54065 9867 54137
rect 7817 54013 7885 54065
rect 7937 54013 8009 54065
rect 8061 54013 8133 54065
rect 8185 54013 8257 54065
rect 8309 54013 8381 54065
rect 8433 54013 8505 54065
rect 8557 54013 8629 54065
rect 8681 54013 9867 54065
rect 7817 53941 9867 54013
rect 7817 53889 7885 53941
rect 7937 53889 8009 53941
rect 8061 53889 8133 53941
rect 8185 53889 8257 53941
rect 8309 53889 8381 53941
rect 8433 53889 8505 53941
rect 8557 53889 8629 53941
rect 8681 53889 9867 53941
rect 7817 53817 9867 53889
rect 7817 53765 7885 53817
rect 7937 53765 8009 53817
rect 8061 53765 8133 53817
rect 8185 53765 8257 53817
rect 8309 53765 8381 53817
rect 8433 53765 8505 53817
rect 8557 53765 8629 53817
rect 8681 53765 9867 53817
rect 7817 53693 9867 53765
rect 7817 53641 7885 53693
rect 7937 53641 8009 53693
rect 8061 53641 8133 53693
rect 8185 53641 8257 53693
rect 8309 53641 8381 53693
rect 8433 53641 8505 53693
rect 8557 53641 8629 53693
rect 8681 53641 9867 53693
rect 7817 52588 9867 53641
rect 7817 52536 7886 52588
rect 7938 52536 8010 52588
rect 8062 52536 8134 52588
rect 8186 52536 8258 52588
rect 8310 52536 8382 52588
rect 8434 52536 8506 52588
rect 8558 52536 8630 52588
rect 8682 52536 8754 52588
rect 8806 52536 8878 52588
rect 8930 52536 9002 52588
rect 9054 52536 9126 52588
rect 9178 52536 9250 52588
rect 9302 52536 9374 52588
rect 9426 52536 9498 52588
rect 9550 52536 9622 52588
rect 9674 52536 9746 52588
rect 9798 52536 9867 52588
rect 7817 52464 9867 52536
rect 7817 52412 7886 52464
rect 7938 52412 8010 52464
rect 8062 52412 8134 52464
rect 8186 52412 8258 52464
rect 8310 52412 8382 52464
rect 8434 52412 8506 52464
rect 8558 52412 8630 52464
rect 8682 52412 8754 52464
rect 8806 52412 8878 52464
rect 8930 52412 9002 52464
rect 9054 52412 9126 52464
rect 9178 52412 9250 52464
rect 9302 52412 9374 52464
rect 9426 52412 9498 52464
rect 9550 52412 9622 52464
rect 9674 52412 9746 52464
rect 9798 52412 9867 52464
rect 7817 52340 9867 52412
rect 7817 52288 7886 52340
rect 7938 52288 8010 52340
rect 8062 52288 8134 52340
rect 8186 52288 8258 52340
rect 8310 52288 8382 52340
rect 8434 52288 8506 52340
rect 8558 52288 8630 52340
rect 8682 52288 8754 52340
rect 8806 52288 8878 52340
rect 8930 52288 9002 52340
rect 9054 52288 9126 52340
rect 9178 52288 9250 52340
rect 9302 52288 9374 52340
rect 9426 52288 9498 52340
rect 9550 52288 9622 52340
rect 9674 52288 9746 52340
rect 9798 52288 9867 52340
rect 7817 51627 9867 52288
rect 7817 51575 7886 51627
rect 7938 51575 8010 51627
rect 8062 51575 8134 51627
rect 8186 51575 8258 51627
rect 8310 51575 8382 51627
rect 8434 51575 8506 51627
rect 8558 51575 8630 51627
rect 8682 51575 8754 51627
rect 8806 51575 8878 51627
rect 8930 51575 9002 51627
rect 9054 51575 9126 51627
rect 9178 51575 9250 51627
rect 9302 51575 9374 51627
rect 9426 51575 9498 51627
rect 9550 51575 9622 51627
rect 9674 51575 9746 51627
rect 9798 51575 9867 51627
rect 7817 51503 9867 51575
rect 7817 51451 7886 51503
rect 7938 51451 8010 51503
rect 8062 51451 8134 51503
rect 8186 51451 8258 51503
rect 8310 51451 8382 51503
rect 8434 51451 8506 51503
rect 8558 51451 8630 51503
rect 8682 51451 8754 51503
rect 8806 51451 8878 51503
rect 8930 51451 9002 51503
rect 9054 51451 9126 51503
rect 9178 51451 9250 51503
rect 9302 51451 9374 51503
rect 9426 51451 9498 51503
rect 9550 51451 9622 51503
rect 9674 51451 9746 51503
rect 9798 51451 9867 51503
rect 7817 50948 9867 51451
rect 7817 50892 7884 50948
rect 7940 50892 8008 50948
rect 8064 50892 8132 50948
rect 8188 50892 8256 50948
rect 8312 50892 8380 50948
rect 8436 50892 8504 50948
rect 8560 50892 8628 50948
rect 8684 50892 8752 50948
rect 8808 50892 8876 50948
rect 8932 50892 9000 50948
rect 9056 50892 9124 50948
rect 9180 50892 9248 50948
rect 9304 50892 9372 50948
rect 9428 50892 9496 50948
rect 9552 50892 9620 50948
rect 9676 50892 9744 50948
rect 9800 50892 9867 50948
rect 7817 50824 9867 50892
rect 7817 50768 7884 50824
rect 7940 50768 8008 50824
rect 8064 50768 8132 50824
rect 8188 50768 8256 50824
rect 8312 50768 8380 50824
rect 8436 50768 8504 50824
rect 8560 50768 8628 50824
rect 8684 50768 8752 50824
rect 8808 50768 8876 50824
rect 8932 50768 9000 50824
rect 9056 50768 9124 50824
rect 9180 50768 9248 50824
rect 9304 50768 9372 50824
rect 9428 50768 9496 50824
rect 9552 50768 9620 50824
rect 9676 50768 9744 50824
rect 9800 50768 9867 50824
rect 7817 50700 9867 50768
rect 7817 50644 7884 50700
rect 7940 50644 8008 50700
rect 8064 50644 8132 50700
rect 8188 50644 8256 50700
rect 8312 50644 8380 50700
rect 8436 50644 8504 50700
rect 8560 50644 8628 50700
rect 8684 50644 8752 50700
rect 8808 50644 8876 50700
rect 8932 50644 9000 50700
rect 9056 50644 9124 50700
rect 9180 50644 9248 50700
rect 9304 50644 9372 50700
rect 9428 50644 9496 50700
rect 9552 50644 9620 50700
rect 9676 50644 9744 50700
rect 9800 50644 9867 50700
rect 7817 50641 7886 50644
rect 7938 50641 8010 50644
rect 8062 50641 8134 50644
rect 8186 50641 8258 50644
rect 8310 50641 8382 50644
rect 8434 50641 8506 50644
rect 8558 50641 8630 50644
rect 8682 50641 8754 50644
rect 8806 50641 8878 50644
rect 8930 50641 9002 50644
rect 9054 50641 9126 50644
rect 9178 50641 9250 50644
rect 9302 50641 9374 50644
rect 9426 50641 9498 50644
rect 9550 50641 9622 50644
rect 9674 50641 9746 50644
rect 9798 50641 9867 50644
rect 7817 50576 9867 50641
rect 7817 50520 7884 50576
rect 7940 50520 8008 50576
rect 8064 50520 8132 50576
rect 8188 50520 8256 50576
rect 8312 50520 8380 50576
rect 8436 50520 8504 50576
rect 8560 50520 8628 50576
rect 8684 50520 8752 50576
rect 8808 50520 8876 50576
rect 8932 50520 9000 50576
rect 9056 50520 9124 50576
rect 9180 50520 9248 50576
rect 9304 50520 9372 50576
rect 9428 50520 9496 50576
rect 9552 50520 9620 50576
rect 9676 50520 9744 50576
rect 9800 50520 9867 50576
rect 7817 50517 7886 50520
rect 7938 50517 8010 50520
rect 8062 50517 8134 50520
rect 8186 50517 8258 50520
rect 8310 50517 8382 50520
rect 8434 50517 8506 50520
rect 8558 50517 8630 50520
rect 8682 50517 8754 50520
rect 8806 50517 8878 50520
rect 8930 50517 9002 50520
rect 9054 50517 9126 50520
rect 9178 50517 9250 50520
rect 9302 50517 9374 50520
rect 9426 50517 9498 50520
rect 9550 50517 9622 50520
rect 9674 50517 9746 50520
rect 9798 50517 9867 50520
rect 7817 50452 9867 50517
rect 7817 50396 7884 50452
rect 7940 50396 8008 50452
rect 8064 50396 8132 50452
rect 8188 50396 8256 50452
rect 8312 50396 8380 50452
rect 8436 50396 8504 50452
rect 8560 50396 8628 50452
rect 8684 50396 8752 50452
rect 8808 50396 8876 50452
rect 8932 50396 9000 50452
rect 9056 50396 9124 50452
rect 9180 50396 9248 50452
rect 9304 50396 9372 50452
rect 9428 50396 9496 50452
rect 9552 50396 9620 50452
rect 9676 50396 9744 50452
rect 9800 50396 9867 50452
rect 7817 50328 9867 50396
rect 7817 50272 7884 50328
rect 7940 50272 8008 50328
rect 8064 50272 8132 50328
rect 8188 50272 8256 50328
rect 8312 50272 8380 50328
rect 8436 50272 8504 50328
rect 8560 50272 8628 50328
rect 8684 50272 8752 50328
rect 8808 50272 8876 50328
rect 8932 50272 9000 50328
rect 9056 50272 9124 50328
rect 9180 50272 9248 50328
rect 9304 50272 9372 50328
rect 9428 50272 9496 50328
rect 9552 50272 9620 50328
rect 9676 50272 9744 50328
rect 9800 50272 9867 50328
rect 7817 50204 9867 50272
rect 7817 50148 7884 50204
rect 7940 50148 8008 50204
rect 8064 50148 8132 50204
rect 8188 50148 8256 50204
rect 8312 50148 8380 50204
rect 8436 50148 8504 50204
rect 8560 50148 8628 50204
rect 8684 50148 8752 50204
rect 8808 50148 8876 50204
rect 8932 50148 9000 50204
rect 9056 50148 9124 50204
rect 9180 50148 9248 50204
rect 9304 50148 9372 50204
rect 9428 50148 9496 50204
rect 9552 50148 9620 50204
rect 9676 50148 9744 50204
rect 9800 50148 9867 50204
rect 7817 50080 9867 50148
rect 7817 50024 7884 50080
rect 7940 50024 8008 50080
rect 8064 50024 8132 50080
rect 8188 50024 8256 50080
rect 8312 50024 8380 50080
rect 8436 50024 8504 50080
rect 8560 50024 8628 50080
rect 8684 50024 8752 50080
rect 8808 50024 8876 50080
rect 8932 50024 9000 50080
rect 9056 50024 9124 50080
rect 9180 50024 9248 50080
rect 9304 50024 9372 50080
rect 9428 50024 9496 50080
rect 9552 50024 9620 50080
rect 9676 50024 9744 50080
rect 9800 50024 9867 50080
rect 7817 49956 9867 50024
rect 7817 49900 7884 49956
rect 7940 49900 8008 49956
rect 8064 49900 8132 49956
rect 8188 49900 8256 49956
rect 8312 49900 8380 49956
rect 8436 49900 8504 49956
rect 8560 49900 8628 49956
rect 8684 49900 8752 49956
rect 8808 49900 8876 49956
rect 8932 49900 9000 49956
rect 9056 49900 9124 49956
rect 9180 49900 9248 49956
rect 9304 49900 9372 49956
rect 9428 49900 9496 49956
rect 9552 49900 9620 49956
rect 9676 49900 9744 49956
rect 9800 49900 9867 49956
rect 7817 49832 9867 49900
rect 7817 49776 7884 49832
rect 7940 49776 8008 49832
rect 8064 49776 8132 49832
rect 8188 49776 8256 49832
rect 8312 49776 8380 49832
rect 8436 49776 8504 49832
rect 8560 49776 8628 49832
rect 8684 49776 8752 49832
rect 8808 49776 8876 49832
rect 8932 49776 9000 49832
rect 9056 49776 9124 49832
rect 9180 49776 9248 49832
rect 9304 49776 9372 49832
rect 9428 49776 9496 49832
rect 9552 49776 9620 49832
rect 9676 49776 9744 49832
rect 9800 49776 9867 49832
rect 7817 49759 9867 49776
rect 7817 49708 7886 49759
rect 7938 49708 8010 49759
rect 8062 49708 8134 49759
rect 8186 49708 8258 49759
rect 8310 49708 8382 49759
rect 8434 49708 8506 49759
rect 8558 49708 8630 49759
rect 8682 49708 8754 49759
rect 8806 49708 8878 49759
rect 8930 49708 9002 49759
rect 9054 49708 9126 49759
rect 9178 49708 9250 49759
rect 9302 49708 9374 49759
rect 9426 49708 9498 49759
rect 9550 49708 9622 49759
rect 9674 49708 9746 49759
rect 9798 49708 9867 49759
rect 7817 49652 7884 49708
rect 7940 49652 8008 49708
rect 8064 49652 8132 49708
rect 8188 49652 8256 49708
rect 8312 49652 8380 49708
rect 8436 49652 8504 49708
rect 8560 49652 8628 49708
rect 8684 49652 8752 49708
rect 8808 49652 8876 49708
rect 8932 49652 9000 49708
rect 9056 49652 9124 49708
rect 9180 49652 9248 49708
rect 9304 49652 9372 49708
rect 9428 49652 9496 49708
rect 9552 49652 9620 49708
rect 9676 49652 9744 49708
rect 9800 49652 9867 49708
rect 7817 49635 9867 49652
rect 7817 49583 7886 49635
rect 7938 49583 8010 49635
rect 8062 49583 8134 49635
rect 8186 49583 8258 49635
rect 8310 49583 8382 49635
rect 8434 49583 8506 49635
rect 8558 49583 8630 49635
rect 8682 49583 8754 49635
rect 8806 49583 8878 49635
rect 8930 49583 9002 49635
rect 9054 49583 9126 49635
rect 9178 49583 9250 49635
rect 9302 49583 9374 49635
rect 9426 49583 9498 49635
rect 9550 49583 9622 49635
rect 9674 49583 9746 49635
rect 9798 49583 9867 49635
rect 7817 48825 9867 49583
rect 7817 48773 7886 48825
rect 7938 48773 8010 48825
rect 8062 48773 8134 48825
rect 8186 48773 8258 48825
rect 8310 48773 8382 48825
rect 8434 48773 8506 48825
rect 8558 48773 8630 48825
rect 8682 48773 8754 48825
rect 8806 48773 8878 48825
rect 8930 48773 9002 48825
rect 9054 48773 9126 48825
rect 9178 48773 9250 48825
rect 9302 48773 9374 48825
rect 9426 48773 9498 48825
rect 9550 48773 9622 48825
rect 9674 48773 9746 48825
rect 9798 48773 9867 48825
rect 7817 48701 9867 48773
rect 7817 48649 7886 48701
rect 7938 48649 8010 48701
rect 8062 48649 8134 48701
rect 8186 48649 8258 48701
rect 8310 48649 8382 48701
rect 8434 48649 8506 48701
rect 8558 48649 8630 48701
rect 8682 48649 8754 48701
rect 8806 48649 8878 48701
rect 8930 48649 9002 48701
rect 9054 48649 9126 48701
rect 9178 48649 9250 48701
rect 9302 48649 9374 48701
rect 9426 48649 9498 48701
rect 9550 48649 9622 48701
rect 9674 48649 9746 48701
rect 9798 48649 9867 48701
rect 7817 47988 9867 48649
rect 7817 47936 7886 47988
rect 7938 47936 8010 47988
rect 8062 47936 8134 47988
rect 8186 47936 8258 47988
rect 8310 47936 8382 47988
rect 8434 47936 8506 47988
rect 8558 47936 8630 47988
rect 8682 47936 8754 47988
rect 8806 47936 8878 47988
rect 8930 47936 9002 47988
rect 9054 47936 9126 47988
rect 9178 47936 9250 47988
rect 9302 47936 9374 47988
rect 9426 47936 9498 47988
rect 9550 47936 9622 47988
rect 9674 47936 9746 47988
rect 9798 47936 9867 47988
rect 7817 47864 9867 47936
rect 7817 47812 7886 47864
rect 7938 47812 8010 47864
rect 8062 47812 8134 47864
rect 8186 47812 8258 47864
rect 8310 47812 8382 47864
rect 8434 47812 8506 47864
rect 8558 47812 8630 47864
rect 8682 47812 8754 47864
rect 8806 47812 8878 47864
rect 8930 47812 9002 47864
rect 9054 47812 9126 47864
rect 9178 47812 9250 47864
rect 9302 47812 9374 47864
rect 9426 47812 9498 47864
rect 9550 47812 9622 47864
rect 9674 47812 9746 47864
rect 9798 47812 9867 47864
rect 7817 47748 9867 47812
rect 7817 47692 7884 47748
rect 7940 47692 8008 47748
rect 8064 47692 8132 47748
rect 8188 47692 8256 47748
rect 8312 47692 8380 47748
rect 8436 47692 8504 47748
rect 8560 47692 8628 47748
rect 8684 47692 8752 47748
rect 8808 47692 8876 47748
rect 8932 47692 9000 47748
rect 9056 47692 9124 47748
rect 9180 47692 9248 47748
rect 9304 47692 9372 47748
rect 9428 47692 9496 47748
rect 9552 47692 9620 47748
rect 9676 47692 9744 47748
rect 9800 47692 9867 47748
rect 7817 47688 7886 47692
rect 7938 47688 8010 47692
rect 8062 47688 8134 47692
rect 8186 47688 8258 47692
rect 8310 47688 8382 47692
rect 8434 47688 8506 47692
rect 8558 47688 8630 47692
rect 8682 47688 8754 47692
rect 8806 47688 8878 47692
rect 8930 47688 9002 47692
rect 9054 47688 9126 47692
rect 9178 47688 9250 47692
rect 9302 47688 9374 47692
rect 9426 47688 9498 47692
rect 9550 47688 9622 47692
rect 9674 47688 9746 47692
rect 9798 47688 9867 47692
rect 7817 47624 9867 47688
rect 7817 47568 7884 47624
rect 7940 47568 8008 47624
rect 8064 47568 8132 47624
rect 8188 47568 8256 47624
rect 8312 47568 8380 47624
rect 8436 47568 8504 47624
rect 8560 47568 8628 47624
rect 8684 47568 8752 47624
rect 8808 47568 8876 47624
rect 8932 47568 9000 47624
rect 9056 47568 9124 47624
rect 9180 47568 9248 47624
rect 9304 47568 9372 47624
rect 9428 47568 9496 47624
rect 9552 47568 9620 47624
rect 9676 47568 9744 47624
rect 9800 47568 9867 47624
rect 7817 47500 9867 47568
rect 7817 47444 7884 47500
rect 7940 47444 8008 47500
rect 8064 47444 8132 47500
rect 8188 47444 8256 47500
rect 8312 47444 8380 47500
rect 8436 47444 8504 47500
rect 8560 47444 8628 47500
rect 8684 47444 8752 47500
rect 8808 47444 8876 47500
rect 8932 47444 9000 47500
rect 9056 47444 9124 47500
rect 9180 47444 9248 47500
rect 9304 47444 9372 47500
rect 9428 47444 9496 47500
rect 9552 47444 9620 47500
rect 9676 47444 9744 47500
rect 9800 47444 9867 47500
rect 7817 47376 9867 47444
rect 7817 47320 7884 47376
rect 7940 47320 8008 47376
rect 8064 47320 8132 47376
rect 8188 47320 8256 47376
rect 8312 47320 8380 47376
rect 8436 47320 8504 47376
rect 8560 47320 8628 47376
rect 8684 47320 8752 47376
rect 8808 47320 8876 47376
rect 8932 47320 9000 47376
rect 9056 47320 9124 47376
rect 9180 47320 9248 47376
rect 9304 47320 9372 47376
rect 9428 47320 9496 47376
rect 9552 47320 9620 47376
rect 9676 47320 9744 47376
rect 9800 47320 9867 47376
rect 7817 47281 9867 47320
rect 9927 57225 10127 57278
rect 9927 57169 9937 57225
rect 9993 57169 10061 57225
rect 10117 57169 10127 57225
rect 9927 57108 10127 57169
rect 9927 57101 9947 57108
rect 9927 57045 9937 57101
rect 9999 57056 10055 57108
rect 10107 57101 10127 57108
rect 9993 57045 10061 57056
rect 10117 57045 10127 57101
rect 9927 56977 10127 57045
rect 9927 56921 9937 56977
rect 9993 56921 10061 56977
rect 10117 56921 10127 56977
rect 9927 56853 10127 56921
rect 9927 56797 9937 56853
rect 9993 56797 10061 56853
rect 10117 56797 10127 56853
rect 9927 56729 10127 56797
rect 9927 56673 9937 56729
rect 9993 56673 10061 56729
rect 10117 56673 10127 56729
rect 9927 56605 10127 56673
rect 9927 56549 9937 56605
rect 9993 56549 10061 56605
rect 10117 56549 10127 56605
rect 9927 56481 10127 56549
rect 9927 56425 9937 56481
rect 9993 56425 10061 56481
rect 10117 56425 10127 56481
rect 9927 56357 10127 56425
rect 9927 56301 9937 56357
rect 9993 56301 10061 56357
rect 10117 56301 10127 56357
rect 9927 56233 10127 56301
rect 9927 56177 9937 56233
rect 9993 56177 10061 56233
rect 10117 56177 10127 56233
rect 9927 56109 10127 56177
rect 9927 56053 9937 56109
rect 9993 56053 10061 56109
rect 10117 56053 10127 56109
rect 9927 54148 10127 56053
rect 9927 54092 9937 54148
rect 9993 54092 10061 54148
rect 10117 54092 10127 54148
rect 9927 54024 10127 54092
rect 9927 53968 9937 54024
rect 9993 53968 10061 54024
rect 10117 53968 10127 54024
rect 9927 53900 10127 53968
rect 9927 53844 9937 53900
rect 9993 53844 10061 53900
rect 10117 53844 10127 53900
rect 9927 53776 10127 53844
rect 9927 53720 9937 53776
rect 9993 53720 10061 53776
rect 10117 53720 10127 53776
rect 9927 53652 10127 53720
rect 9927 53596 9937 53652
rect 9993 53596 10061 53652
rect 10117 53596 10127 53652
rect 9927 53528 10127 53596
rect 9927 53472 9937 53528
rect 9993 53484 10061 53528
rect 9927 53432 9947 53472
rect 9999 53432 10055 53484
rect 10117 53472 10127 53528
rect 10107 53432 10127 53472
rect 9927 53404 10127 53432
rect 9927 53348 9937 53404
rect 9993 53376 10061 53404
rect 9927 53324 9947 53348
rect 9999 53324 10055 53376
rect 10117 53348 10127 53404
rect 10107 53324 10127 53348
rect 9927 53280 10127 53324
rect 9927 53224 9937 53280
rect 9993 53268 10061 53280
rect 9927 53216 9947 53224
rect 9999 53216 10055 53268
rect 10117 53224 10127 53280
rect 10107 53216 10127 53224
rect 9927 53156 10127 53216
rect 9927 53100 9937 53156
rect 9993 53100 10061 53156
rect 10117 53100 10127 53156
rect 9927 53032 10127 53100
rect 9927 52976 9937 53032
rect 9993 52976 10061 53032
rect 10117 52976 10127 53032
rect 9927 52908 10127 52976
rect 9927 52852 9937 52908
rect 9993 52852 10061 52908
rect 10117 52852 10127 52908
rect 9927 52017 10127 52852
rect 9927 51965 9939 52017
rect 9991 51965 10063 52017
rect 10115 51965 10127 52017
rect 9927 51893 10127 51965
rect 9927 51841 9939 51893
rect 9991 51841 10063 51893
rect 10115 51841 10127 51893
rect 9927 51222 10127 51841
rect 9927 51170 9939 51222
rect 9991 51170 10063 51222
rect 10115 51170 10127 51222
rect 9927 51098 10127 51170
rect 9927 51046 9939 51098
rect 9991 51046 10063 51098
rect 10115 51046 10127 51098
rect 9927 50974 10127 51046
rect 9927 50922 9939 50974
rect 9991 50922 10063 50974
rect 10115 50922 10127 50974
rect 9927 50288 10127 50922
rect 9927 50236 9939 50288
rect 9991 50236 10063 50288
rect 10115 50236 10127 50288
rect 9927 50164 10127 50236
rect 9927 50112 9939 50164
rect 9991 50112 10063 50164
rect 10115 50112 10127 50164
rect 9927 50040 10127 50112
rect 9927 49988 9939 50040
rect 9991 49988 10063 50040
rect 10115 49988 10127 50040
rect 9927 49354 10127 49988
rect 9927 49348 9939 49354
rect 9991 49348 10063 49354
rect 10115 49348 10127 49354
rect 9927 49292 9937 49348
rect 9993 49292 10061 49348
rect 10117 49292 10127 49348
rect 9927 49230 10127 49292
rect 9927 49224 9939 49230
rect 9991 49224 10063 49230
rect 10115 49224 10127 49230
rect 9927 49168 9937 49224
rect 9993 49168 10061 49224
rect 10117 49168 10127 49224
rect 9927 49106 10127 49168
rect 9927 49100 9939 49106
rect 9991 49100 10063 49106
rect 10115 49100 10127 49106
rect 9927 49044 9937 49100
rect 9993 49044 10061 49100
rect 10117 49044 10127 49100
rect 9927 48976 10127 49044
rect 9927 48920 9937 48976
rect 9993 48920 10061 48976
rect 10117 48920 10127 48976
rect 9927 48852 10127 48920
rect 9927 48796 9937 48852
rect 9993 48796 10061 48852
rect 10117 48796 10127 48852
rect 9927 48728 10127 48796
rect 9927 48672 9937 48728
rect 9993 48672 10061 48728
rect 10117 48672 10127 48728
rect 9927 48604 10127 48672
rect 9927 48548 9937 48604
rect 9993 48548 10061 48604
rect 10117 48548 10127 48604
rect 9927 48480 10127 48548
rect 9927 48424 9937 48480
rect 9993 48424 10061 48480
rect 10117 48424 10127 48480
rect 9927 48383 9939 48424
rect 9991 48383 10063 48424
rect 10115 48383 10127 48424
rect 9927 48356 10127 48383
rect 9927 48300 9937 48356
rect 9993 48300 10061 48356
rect 10117 48300 10127 48356
rect 9927 48259 9939 48300
rect 9991 48259 10063 48300
rect 10115 48259 10127 48300
rect 9927 48232 10127 48259
rect 9927 48176 9937 48232
rect 9993 48176 10061 48232
rect 10117 48176 10127 48232
rect 9927 48108 10127 48176
rect 9927 48052 9937 48108
rect 9993 48052 10061 48108
rect 10117 48052 10127 48108
rect 9927 47281 10127 48052
rect 10187 56669 12237 57600
rect 10187 56617 10214 56669
rect 10266 56617 10338 56669
rect 10390 56617 10462 56669
rect 10514 56617 10586 56669
rect 10638 56617 11225 56669
rect 11277 56617 11349 56669
rect 11401 56617 11473 56669
rect 11525 56617 11597 56669
rect 11649 56617 11721 56669
rect 11773 56617 11845 56669
rect 11897 56617 11969 56669
rect 12021 56617 12093 56669
rect 12145 56617 12237 56669
rect 10187 56545 12237 56617
rect 10187 56493 10214 56545
rect 10266 56493 10338 56545
rect 10390 56493 10462 56545
rect 10514 56493 10586 56545
rect 10638 56493 11225 56545
rect 11277 56493 11349 56545
rect 11401 56493 11473 56545
rect 11525 56493 11597 56545
rect 11649 56493 11721 56545
rect 11773 56493 11845 56545
rect 11897 56493 11969 56545
rect 12021 56493 12093 56545
rect 12145 56493 12237 56545
rect 10187 56421 12237 56493
rect 10187 56369 10214 56421
rect 10266 56369 10338 56421
rect 10390 56369 10462 56421
rect 10514 56369 10586 56421
rect 10638 56369 11225 56421
rect 11277 56369 11349 56421
rect 11401 56369 11473 56421
rect 11525 56369 11597 56421
rect 11649 56369 11721 56421
rect 11773 56369 11845 56421
rect 11897 56369 11969 56421
rect 12021 56369 12093 56421
rect 12145 56369 12237 56421
rect 10187 56297 12237 56369
rect 10187 56245 10214 56297
rect 10266 56245 10338 56297
rect 10390 56245 10462 56297
rect 10514 56245 10586 56297
rect 10638 56245 11225 56297
rect 11277 56245 11349 56297
rect 11401 56245 11473 56297
rect 11525 56245 11597 56297
rect 11649 56245 11721 56297
rect 11773 56245 11845 56297
rect 11897 56245 11969 56297
rect 12021 56245 12093 56297
rect 12145 56245 12237 56297
rect 10187 56173 12237 56245
rect 10187 56121 10214 56173
rect 10266 56121 10338 56173
rect 10390 56121 10462 56173
rect 10514 56121 10586 56173
rect 10638 56121 11225 56173
rect 11277 56121 11349 56173
rect 11401 56121 11473 56173
rect 11525 56121 11597 56173
rect 11649 56121 11721 56173
rect 11773 56121 11845 56173
rect 11897 56121 11969 56173
rect 12021 56121 12093 56173
rect 12145 56121 12237 56173
rect 10187 56049 12237 56121
rect 10187 55997 10214 56049
rect 10266 55997 10338 56049
rect 10390 55997 10462 56049
rect 10514 55997 10586 56049
rect 10638 55997 11225 56049
rect 11277 55997 11349 56049
rect 11401 55997 11473 56049
rect 11525 55997 11597 56049
rect 11649 55997 11721 56049
rect 11773 55997 11845 56049
rect 11897 55997 11969 56049
rect 12021 55997 12093 56049
rect 12145 55997 12237 56049
rect 10187 55925 12237 55997
rect 10187 55873 10214 55925
rect 10266 55873 10338 55925
rect 10390 55873 10462 55925
rect 10514 55873 10586 55925
rect 10638 55873 11225 55925
rect 11277 55873 11349 55925
rect 11401 55873 11473 55925
rect 11525 55873 11597 55925
rect 11649 55873 11721 55925
rect 11773 55873 11845 55925
rect 11897 55873 11969 55925
rect 12021 55873 12093 55925
rect 12145 55873 12237 55925
rect 10187 55801 12237 55873
rect 10187 55749 10214 55801
rect 10266 55749 10338 55801
rect 10390 55749 10462 55801
rect 10514 55749 10586 55801
rect 10638 55749 11225 55801
rect 11277 55749 11349 55801
rect 11401 55749 11473 55801
rect 11525 55749 11597 55801
rect 11649 55749 11721 55801
rect 11773 55749 11845 55801
rect 11897 55749 11969 55801
rect 12021 55749 12093 55801
rect 12145 55749 12237 55801
rect 10187 55748 12237 55749
rect 10187 55692 10254 55748
rect 10310 55692 10378 55748
rect 10434 55692 10502 55748
rect 10558 55692 10626 55748
rect 10682 55692 10750 55748
rect 10806 55692 10874 55748
rect 10930 55692 10998 55748
rect 11054 55692 11122 55748
rect 11178 55692 11246 55748
rect 11302 55692 11370 55748
rect 11426 55692 11494 55748
rect 11550 55692 11618 55748
rect 11674 55692 11742 55748
rect 11798 55692 11866 55748
rect 11922 55692 11990 55748
rect 12046 55692 12114 55748
rect 12170 55692 12237 55748
rect 10187 55677 12237 55692
rect 10187 55625 10214 55677
rect 10266 55625 10338 55677
rect 10390 55625 10462 55677
rect 10514 55625 10586 55677
rect 10638 55625 11225 55677
rect 11277 55625 11349 55677
rect 11401 55625 11473 55677
rect 11525 55625 11597 55677
rect 11649 55625 11721 55677
rect 11773 55625 11845 55677
rect 11897 55625 11969 55677
rect 12021 55625 12093 55677
rect 12145 55625 12237 55677
rect 10187 55624 12237 55625
rect 10187 55568 10254 55624
rect 10310 55568 10378 55624
rect 10434 55568 10502 55624
rect 10558 55568 10626 55624
rect 10682 55568 10750 55624
rect 10806 55568 10874 55624
rect 10930 55568 10998 55624
rect 11054 55568 11122 55624
rect 11178 55568 11246 55624
rect 11302 55568 11370 55624
rect 11426 55568 11494 55624
rect 11550 55568 11618 55624
rect 11674 55568 11742 55624
rect 11798 55568 11866 55624
rect 11922 55568 11990 55624
rect 12046 55568 12114 55624
rect 12170 55568 12237 55624
rect 10187 55553 12237 55568
rect 10187 55501 10214 55553
rect 10266 55501 10338 55553
rect 10390 55501 10462 55553
rect 10514 55501 10586 55553
rect 10638 55501 11225 55553
rect 11277 55501 11349 55553
rect 11401 55501 11473 55553
rect 11525 55501 11597 55553
rect 11649 55501 11721 55553
rect 11773 55501 11845 55553
rect 11897 55501 11969 55553
rect 12021 55501 12093 55553
rect 12145 55501 12237 55553
rect 10187 55500 12237 55501
rect 10187 55444 10254 55500
rect 10310 55444 10378 55500
rect 10434 55444 10502 55500
rect 10558 55444 10626 55500
rect 10682 55444 10750 55500
rect 10806 55444 10874 55500
rect 10930 55444 10998 55500
rect 11054 55444 11122 55500
rect 11178 55444 11246 55500
rect 11302 55444 11370 55500
rect 11426 55444 11494 55500
rect 11550 55444 11618 55500
rect 11674 55444 11742 55500
rect 11798 55444 11866 55500
rect 11922 55444 11990 55500
rect 12046 55444 12114 55500
rect 12170 55444 12237 55500
rect 10187 55429 12237 55444
rect 10187 55377 10214 55429
rect 10266 55377 10338 55429
rect 10390 55377 10462 55429
rect 10514 55377 10586 55429
rect 10638 55377 11225 55429
rect 11277 55377 11349 55429
rect 11401 55377 11473 55429
rect 11525 55377 11597 55429
rect 11649 55377 11721 55429
rect 11773 55377 11845 55429
rect 11897 55377 11969 55429
rect 12021 55377 12093 55429
rect 12145 55377 12237 55429
rect 10187 55376 12237 55377
rect 10187 55320 10254 55376
rect 10310 55320 10378 55376
rect 10434 55320 10502 55376
rect 10558 55320 10626 55376
rect 10682 55320 10750 55376
rect 10806 55320 10874 55376
rect 10930 55320 10998 55376
rect 11054 55320 11122 55376
rect 11178 55320 11246 55376
rect 11302 55320 11370 55376
rect 11426 55320 11494 55376
rect 11550 55320 11618 55376
rect 11674 55320 11742 55376
rect 11798 55320 11866 55376
rect 11922 55320 11990 55376
rect 12046 55320 12114 55376
rect 12170 55320 12237 55376
rect 10187 55305 12237 55320
rect 10187 55253 10214 55305
rect 10266 55253 10338 55305
rect 10390 55253 10462 55305
rect 10514 55253 10586 55305
rect 10638 55253 11225 55305
rect 11277 55253 11349 55305
rect 11401 55253 11473 55305
rect 11525 55253 11597 55305
rect 11649 55253 11721 55305
rect 11773 55253 11845 55305
rect 11897 55253 11969 55305
rect 12021 55253 12093 55305
rect 12145 55253 12237 55305
rect 10187 55252 12237 55253
rect 10187 55196 10254 55252
rect 10310 55196 10378 55252
rect 10434 55196 10502 55252
rect 10558 55196 10626 55252
rect 10682 55196 10750 55252
rect 10806 55196 10874 55252
rect 10930 55196 10998 55252
rect 11054 55196 11122 55252
rect 11178 55196 11246 55252
rect 11302 55196 11370 55252
rect 11426 55196 11494 55252
rect 11550 55196 11618 55252
rect 11674 55196 11742 55252
rect 11798 55196 11866 55252
rect 11922 55196 11990 55252
rect 12046 55196 12114 55252
rect 12170 55196 12237 55252
rect 10187 55181 12237 55196
rect 10187 55129 10214 55181
rect 10266 55129 10338 55181
rect 10390 55129 10462 55181
rect 10514 55129 10586 55181
rect 10638 55129 11225 55181
rect 11277 55129 11349 55181
rect 11401 55129 11473 55181
rect 11525 55129 11597 55181
rect 11649 55129 11721 55181
rect 11773 55129 11845 55181
rect 11897 55129 11969 55181
rect 12021 55129 12093 55181
rect 12145 55129 12237 55181
rect 10187 55128 12237 55129
rect 10187 55072 10254 55128
rect 10310 55072 10378 55128
rect 10434 55072 10502 55128
rect 10558 55072 10626 55128
rect 10682 55072 10750 55128
rect 10806 55072 10874 55128
rect 10930 55072 10998 55128
rect 11054 55072 11122 55128
rect 11178 55072 11246 55128
rect 11302 55072 11370 55128
rect 11426 55072 11494 55128
rect 11550 55072 11618 55128
rect 11674 55072 11742 55128
rect 11798 55072 11866 55128
rect 11922 55072 11990 55128
rect 12046 55072 12114 55128
rect 12170 55072 12237 55128
rect 10187 55057 12237 55072
rect 10187 55005 10214 55057
rect 10266 55005 10338 55057
rect 10390 55005 10462 55057
rect 10514 55005 10586 55057
rect 10638 55005 11225 55057
rect 11277 55005 11349 55057
rect 11401 55005 11473 55057
rect 11525 55005 11597 55057
rect 11649 55005 11721 55057
rect 11773 55005 11845 55057
rect 11897 55005 11969 55057
rect 12021 55005 12093 55057
rect 12145 55005 12237 55057
rect 10187 55004 12237 55005
rect 10187 54948 10254 55004
rect 10310 54948 10378 55004
rect 10434 54948 10502 55004
rect 10558 54948 10626 55004
rect 10682 54948 10750 55004
rect 10806 54948 10874 55004
rect 10930 54948 10998 55004
rect 11054 54948 11122 55004
rect 11178 54948 11246 55004
rect 11302 54948 11370 55004
rect 11426 54948 11494 55004
rect 11550 54948 11618 55004
rect 11674 54948 11742 55004
rect 11798 54948 11866 55004
rect 11922 54948 11990 55004
rect 12046 54948 12114 55004
rect 12170 54948 12237 55004
rect 10187 54933 12237 54948
rect 10187 54881 10214 54933
rect 10266 54881 10338 54933
rect 10390 54881 10462 54933
rect 10514 54881 10586 54933
rect 10638 54881 11225 54933
rect 11277 54881 11349 54933
rect 11401 54881 11473 54933
rect 11525 54881 11597 54933
rect 11649 54881 11721 54933
rect 11773 54881 11845 54933
rect 11897 54881 11969 54933
rect 12021 54881 12093 54933
rect 12145 54881 12237 54933
rect 10187 54880 12237 54881
rect 10187 54824 10254 54880
rect 10310 54824 10378 54880
rect 10434 54824 10502 54880
rect 10558 54824 10626 54880
rect 10682 54824 10750 54880
rect 10806 54824 10874 54880
rect 10930 54824 10998 54880
rect 11054 54824 11122 54880
rect 11178 54824 11246 54880
rect 11302 54824 11370 54880
rect 11426 54824 11494 54880
rect 11550 54824 11618 54880
rect 11674 54824 11742 54880
rect 11798 54824 11866 54880
rect 11922 54824 11990 54880
rect 12046 54824 12114 54880
rect 12170 54824 12237 54880
rect 10187 54809 12237 54824
rect 10187 54757 10214 54809
rect 10266 54757 10338 54809
rect 10390 54757 10462 54809
rect 10514 54757 10586 54809
rect 10638 54757 11225 54809
rect 11277 54757 11349 54809
rect 11401 54757 11473 54809
rect 11525 54757 11597 54809
rect 11649 54757 11721 54809
rect 11773 54757 11845 54809
rect 11897 54757 11969 54809
rect 12021 54757 12093 54809
rect 12145 54757 12237 54809
rect 10187 54756 12237 54757
rect 10187 54700 10254 54756
rect 10310 54700 10378 54756
rect 10434 54700 10502 54756
rect 10558 54700 10626 54756
rect 10682 54700 10750 54756
rect 10806 54700 10874 54756
rect 10930 54700 10998 54756
rect 11054 54700 11122 54756
rect 11178 54700 11246 54756
rect 11302 54700 11370 54756
rect 11426 54700 11494 54756
rect 11550 54700 11618 54756
rect 11674 54700 11742 54756
rect 11798 54700 11866 54756
rect 11922 54700 11990 54756
rect 12046 54700 12114 54756
rect 12170 54700 12237 54756
rect 10187 54685 12237 54700
rect 10187 54633 10214 54685
rect 10266 54633 10338 54685
rect 10390 54633 10462 54685
rect 10514 54633 10586 54685
rect 10638 54633 11225 54685
rect 11277 54633 11349 54685
rect 11401 54633 11473 54685
rect 11525 54633 11597 54685
rect 11649 54633 11721 54685
rect 11773 54633 11845 54685
rect 11897 54633 11969 54685
rect 12021 54633 12093 54685
rect 12145 54633 12237 54685
rect 10187 54632 12237 54633
rect 10187 54576 10254 54632
rect 10310 54576 10378 54632
rect 10434 54576 10502 54632
rect 10558 54576 10626 54632
rect 10682 54576 10750 54632
rect 10806 54576 10874 54632
rect 10930 54576 10998 54632
rect 11054 54576 11122 54632
rect 11178 54576 11246 54632
rect 11302 54576 11370 54632
rect 11426 54576 11494 54632
rect 11550 54576 11618 54632
rect 11674 54576 11742 54632
rect 11798 54576 11866 54632
rect 11922 54576 11990 54632
rect 12046 54576 12114 54632
rect 12170 54576 12237 54632
rect 10187 54561 12237 54576
rect 10187 54509 10214 54561
rect 10266 54509 10338 54561
rect 10390 54509 10462 54561
rect 10514 54509 10586 54561
rect 10638 54509 11225 54561
rect 11277 54509 11349 54561
rect 11401 54509 11473 54561
rect 11525 54509 11597 54561
rect 11649 54509 11721 54561
rect 11773 54509 11845 54561
rect 11897 54509 11969 54561
rect 12021 54509 12093 54561
rect 12145 54509 12237 54561
rect 10187 54508 12237 54509
rect 10187 54452 10254 54508
rect 10310 54452 10378 54508
rect 10434 54452 10502 54508
rect 10558 54452 10626 54508
rect 10682 54452 10750 54508
rect 10806 54452 10874 54508
rect 10930 54452 10998 54508
rect 11054 54452 11122 54508
rect 11178 54452 11246 54508
rect 11302 54452 11370 54508
rect 11426 54452 11494 54508
rect 11550 54452 11618 54508
rect 11674 54452 11742 54508
rect 11798 54452 11866 54508
rect 11922 54452 11990 54508
rect 12046 54452 12114 54508
rect 12170 54452 12237 54508
rect 10187 54437 12237 54452
rect 10187 54385 10214 54437
rect 10266 54385 10338 54437
rect 10390 54385 10462 54437
rect 10514 54385 10586 54437
rect 10638 54385 11225 54437
rect 11277 54385 11349 54437
rect 11401 54385 11473 54437
rect 11525 54385 11597 54437
rect 11649 54385 11721 54437
rect 11773 54385 11845 54437
rect 11897 54385 11969 54437
rect 12021 54385 12093 54437
rect 12145 54385 12237 54437
rect 10187 54313 12237 54385
rect 10187 54261 10214 54313
rect 10266 54261 10338 54313
rect 10390 54261 10462 54313
rect 10514 54261 10586 54313
rect 10638 54261 11225 54313
rect 11277 54261 11349 54313
rect 11401 54261 11473 54313
rect 11525 54261 11597 54313
rect 11649 54261 11721 54313
rect 11773 54261 11845 54313
rect 11897 54261 11969 54313
rect 12021 54261 12093 54313
rect 12145 54261 12237 54313
rect 10187 54189 12237 54261
rect 10187 54137 10214 54189
rect 10266 54137 10338 54189
rect 10390 54137 10462 54189
rect 10514 54137 10586 54189
rect 10638 54137 11225 54189
rect 11277 54137 11349 54189
rect 11401 54137 11473 54189
rect 11525 54137 11597 54189
rect 11649 54137 11721 54189
rect 11773 54137 11845 54189
rect 11897 54137 11969 54189
rect 12021 54137 12093 54189
rect 12145 54137 12237 54189
rect 10187 54065 12237 54137
rect 10187 54013 10214 54065
rect 10266 54013 10338 54065
rect 10390 54013 10462 54065
rect 10514 54013 10586 54065
rect 10638 54013 11225 54065
rect 11277 54013 11349 54065
rect 11401 54013 11473 54065
rect 11525 54013 11597 54065
rect 11649 54013 11721 54065
rect 11773 54013 11845 54065
rect 11897 54013 11969 54065
rect 12021 54013 12093 54065
rect 12145 54013 12237 54065
rect 10187 53941 12237 54013
rect 10187 53889 10214 53941
rect 10266 53889 10338 53941
rect 10390 53889 10462 53941
rect 10514 53889 10586 53941
rect 10638 53889 11225 53941
rect 11277 53889 11349 53941
rect 11401 53889 11473 53941
rect 11525 53889 11597 53941
rect 11649 53889 11721 53941
rect 11773 53889 11845 53941
rect 11897 53889 11969 53941
rect 12021 53889 12093 53941
rect 12145 53889 12237 53941
rect 10187 53817 12237 53889
rect 10187 53765 10214 53817
rect 10266 53765 10338 53817
rect 10390 53765 10462 53817
rect 10514 53765 10586 53817
rect 10638 53765 11225 53817
rect 11277 53765 11349 53817
rect 11401 53765 11473 53817
rect 11525 53765 11597 53817
rect 11649 53765 11721 53817
rect 11773 53765 11845 53817
rect 11897 53765 11969 53817
rect 12021 53765 12093 53817
rect 12145 53765 12237 53817
rect 10187 53693 12237 53765
rect 10187 53641 10214 53693
rect 10266 53641 10338 53693
rect 10390 53641 10462 53693
rect 10514 53641 10586 53693
rect 10638 53641 11225 53693
rect 11277 53641 11349 53693
rect 11401 53641 11473 53693
rect 11525 53641 11597 53693
rect 11649 53641 11721 53693
rect 11773 53641 11845 53693
rect 11897 53641 11969 53693
rect 12021 53641 12093 53693
rect 12145 53641 12237 53693
rect 10187 52588 12237 53641
rect 10187 52536 10256 52588
rect 10308 52536 10380 52588
rect 10432 52536 10504 52588
rect 10556 52536 10628 52588
rect 10680 52536 10752 52588
rect 10804 52536 10876 52588
rect 10928 52536 11000 52588
rect 11052 52536 11124 52588
rect 11176 52536 11248 52588
rect 11300 52536 11372 52588
rect 11424 52536 11496 52588
rect 11548 52536 11620 52588
rect 11672 52536 11744 52588
rect 11796 52536 11868 52588
rect 11920 52536 11992 52588
rect 12044 52536 12116 52588
rect 12168 52536 12237 52588
rect 10187 52464 12237 52536
rect 10187 52412 10256 52464
rect 10308 52412 10380 52464
rect 10432 52412 10504 52464
rect 10556 52412 10628 52464
rect 10680 52412 10752 52464
rect 10804 52412 10876 52464
rect 10928 52412 11000 52464
rect 11052 52412 11124 52464
rect 11176 52412 11248 52464
rect 11300 52412 11372 52464
rect 11424 52412 11496 52464
rect 11548 52412 11620 52464
rect 11672 52412 11744 52464
rect 11796 52412 11868 52464
rect 11920 52412 11992 52464
rect 12044 52412 12116 52464
rect 12168 52412 12237 52464
rect 10187 52340 12237 52412
rect 10187 52288 10256 52340
rect 10308 52288 10380 52340
rect 10432 52288 10504 52340
rect 10556 52288 10628 52340
rect 10680 52288 10752 52340
rect 10804 52288 10876 52340
rect 10928 52288 11000 52340
rect 11052 52288 11124 52340
rect 11176 52288 11248 52340
rect 11300 52288 11372 52340
rect 11424 52288 11496 52340
rect 11548 52288 11620 52340
rect 11672 52288 11744 52340
rect 11796 52288 11868 52340
rect 11920 52288 11992 52340
rect 12044 52288 12116 52340
rect 12168 52288 12237 52340
rect 10187 51627 12237 52288
rect 10187 51575 10251 51627
rect 10303 51575 10375 51627
rect 10427 51575 10499 51627
rect 10551 51575 10623 51627
rect 10675 51575 10747 51627
rect 10799 51575 10871 51627
rect 10923 51575 10995 51627
rect 11047 51575 11119 51627
rect 11171 51575 11243 51627
rect 11295 51575 11367 51627
rect 11419 51575 12237 51627
rect 10187 51503 12237 51575
rect 10187 51451 10251 51503
rect 10303 51451 10375 51503
rect 10427 51451 10499 51503
rect 10551 51451 10623 51503
rect 10675 51451 10747 51503
rect 10799 51451 10871 51503
rect 10923 51451 10995 51503
rect 11047 51451 11119 51503
rect 11171 51451 11243 51503
rect 11295 51451 11367 51503
rect 11419 51451 12237 51503
rect 10187 50948 12237 51451
rect 10187 50892 10254 50948
rect 10310 50892 10378 50948
rect 10434 50892 10502 50948
rect 10558 50892 10626 50948
rect 10682 50892 10750 50948
rect 10806 50892 10874 50948
rect 10930 50892 10998 50948
rect 11054 50892 11122 50948
rect 11178 50892 11246 50948
rect 11302 50892 11370 50948
rect 11426 50892 11494 50948
rect 11550 50892 11618 50948
rect 11674 50892 11742 50948
rect 11798 50892 11866 50948
rect 11922 50892 11990 50948
rect 12046 50892 12114 50948
rect 12170 50892 12237 50948
rect 10187 50824 12237 50892
rect 10187 50768 10254 50824
rect 10310 50768 10378 50824
rect 10434 50768 10502 50824
rect 10558 50768 10626 50824
rect 10682 50768 10750 50824
rect 10806 50768 10874 50824
rect 10930 50768 10998 50824
rect 11054 50768 11122 50824
rect 11178 50768 11246 50824
rect 11302 50768 11370 50824
rect 11426 50768 11494 50824
rect 11550 50768 11618 50824
rect 11674 50768 11742 50824
rect 11798 50768 11866 50824
rect 11922 50768 11990 50824
rect 12046 50768 12114 50824
rect 12170 50768 12237 50824
rect 10187 50700 12237 50768
rect 10187 50693 10254 50700
rect 10310 50693 10378 50700
rect 10434 50693 10502 50700
rect 10558 50693 10626 50700
rect 10682 50693 10750 50700
rect 10806 50693 10874 50700
rect 10930 50693 10998 50700
rect 11054 50693 11122 50700
rect 11178 50693 11246 50700
rect 11302 50693 11370 50700
rect 10187 50641 10251 50693
rect 10310 50644 10375 50693
rect 10434 50644 10499 50693
rect 10558 50644 10623 50693
rect 10682 50644 10747 50693
rect 10806 50644 10871 50693
rect 10930 50644 10995 50693
rect 11054 50644 11119 50693
rect 11178 50644 11243 50693
rect 11302 50644 11367 50693
rect 11426 50644 11494 50700
rect 11550 50644 11618 50700
rect 11674 50644 11742 50700
rect 11798 50644 11866 50700
rect 11922 50644 11990 50700
rect 12046 50644 12114 50700
rect 12170 50644 12237 50700
rect 10303 50641 10375 50644
rect 10427 50641 10499 50644
rect 10551 50641 10623 50644
rect 10675 50641 10747 50644
rect 10799 50641 10871 50644
rect 10923 50641 10995 50644
rect 11047 50641 11119 50644
rect 11171 50641 11243 50644
rect 11295 50641 11367 50644
rect 11419 50641 12237 50644
rect 10187 50576 12237 50641
rect 10187 50569 10254 50576
rect 10310 50569 10378 50576
rect 10434 50569 10502 50576
rect 10558 50569 10626 50576
rect 10682 50569 10750 50576
rect 10806 50569 10874 50576
rect 10930 50569 10998 50576
rect 11054 50569 11122 50576
rect 11178 50569 11246 50576
rect 11302 50569 11370 50576
rect 10187 50517 10251 50569
rect 10310 50520 10375 50569
rect 10434 50520 10499 50569
rect 10558 50520 10623 50569
rect 10682 50520 10747 50569
rect 10806 50520 10871 50569
rect 10930 50520 10995 50569
rect 11054 50520 11119 50569
rect 11178 50520 11243 50569
rect 11302 50520 11367 50569
rect 11426 50520 11494 50576
rect 11550 50520 11618 50576
rect 11674 50520 11742 50576
rect 11798 50520 11866 50576
rect 11922 50520 11990 50576
rect 12046 50520 12114 50576
rect 12170 50520 12237 50576
rect 10303 50517 10375 50520
rect 10427 50517 10499 50520
rect 10551 50517 10623 50520
rect 10675 50517 10747 50520
rect 10799 50517 10871 50520
rect 10923 50517 10995 50520
rect 11047 50517 11119 50520
rect 11171 50517 11243 50520
rect 11295 50517 11367 50520
rect 11419 50517 12237 50520
rect 10187 50452 12237 50517
rect 10187 50396 10254 50452
rect 10310 50396 10378 50452
rect 10434 50396 10502 50452
rect 10558 50396 10626 50452
rect 10682 50396 10750 50452
rect 10806 50396 10874 50452
rect 10930 50396 10998 50452
rect 11054 50396 11122 50452
rect 11178 50396 11246 50452
rect 11302 50396 11370 50452
rect 11426 50396 11494 50452
rect 11550 50396 11618 50452
rect 11674 50396 11742 50452
rect 11798 50396 11866 50452
rect 11922 50396 11990 50452
rect 12046 50396 12114 50452
rect 12170 50396 12237 50452
rect 10187 50328 12237 50396
rect 10187 50272 10254 50328
rect 10310 50272 10378 50328
rect 10434 50272 10502 50328
rect 10558 50272 10626 50328
rect 10682 50272 10750 50328
rect 10806 50272 10874 50328
rect 10930 50272 10998 50328
rect 11054 50272 11122 50328
rect 11178 50272 11246 50328
rect 11302 50272 11370 50328
rect 11426 50272 11494 50328
rect 11550 50272 11618 50328
rect 11674 50272 11742 50328
rect 11798 50272 11866 50328
rect 11922 50272 11990 50328
rect 12046 50272 12114 50328
rect 12170 50272 12237 50328
rect 10187 50204 12237 50272
rect 10187 50148 10254 50204
rect 10310 50148 10378 50204
rect 10434 50148 10502 50204
rect 10558 50148 10626 50204
rect 10682 50148 10750 50204
rect 10806 50148 10874 50204
rect 10930 50148 10998 50204
rect 11054 50148 11122 50204
rect 11178 50148 11246 50204
rect 11302 50148 11370 50204
rect 11426 50148 11494 50204
rect 11550 50148 11618 50204
rect 11674 50148 11742 50204
rect 11798 50148 11866 50204
rect 11922 50148 11990 50204
rect 12046 50148 12114 50204
rect 12170 50148 12237 50204
rect 10187 50080 12237 50148
rect 10187 50024 10254 50080
rect 10310 50024 10378 50080
rect 10434 50024 10502 50080
rect 10558 50024 10626 50080
rect 10682 50024 10750 50080
rect 10806 50024 10874 50080
rect 10930 50024 10998 50080
rect 11054 50024 11122 50080
rect 11178 50024 11246 50080
rect 11302 50024 11370 50080
rect 11426 50024 11494 50080
rect 11550 50024 11618 50080
rect 11674 50024 11742 50080
rect 11798 50024 11866 50080
rect 11922 50024 11990 50080
rect 12046 50024 12114 50080
rect 12170 50024 12237 50080
rect 10187 49956 12237 50024
rect 10187 49900 10254 49956
rect 10310 49900 10378 49956
rect 10434 49900 10502 49956
rect 10558 49900 10626 49956
rect 10682 49900 10750 49956
rect 10806 49900 10874 49956
rect 10930 49900 10998 49956
rect 11054 49900 11122 49956
rect 11178 49900 11246 49956
rect 11302 49900 11370 49956
rect 11426 49900 11494 49956
rect 11550 49900 11618 49956
rect 11674 49900 11742 49956
rect 11798 49900 11866 49956
rect 11922 49900 11990 49956
rect 12046 49900 12114 49956
rect 12170 49900 12237 49956
rect 10187 49832 12237 49900
rect 10187 49776 10254 49832
rect 10310 49776 10378 49832
rect 10434 49776 10502 49832
rect 10558 49776 10626 49832
rect 10682 49776 10750 49832
rect 10806 49776 10874 49832
rect 10930 49776 10998 49832
rect 11054 49776 11122 49832
rect 11178 49776 11246 49832
rect 11302 49776 11370 49832
rect 11426 49776 11494 49832
rect 11550 49776 11618 49832
rect 11674 49776 11742 49832
rect 11798 49776 11866 49832
rect 11922 49776 11990 49832
rect 12046 49776 12114 49832
rect 12170 49776 12237 49832
rect 10187 49759 12237 49776
rect 10187 49707 10251 49759
rect 10303 49708 10375 49759
rect 10427 49708 10499 49759
rect 10551 49708 10623 49759
rect 10675 49708 10747 49759
rect 10799 49708 10871 49759
rect 10923 49708 10995 49759
rect 11047 49708 11119 49759
rect 11171 49708 11243 49759
rect 11295 49708 11367 49759
rect 11419 49708 12237 49759
rect 10310 49707 10375 49708
rect 10434 49707 10499 49708
rect 10558 49707 10623 49708
rect 10682 49707 10747 49708
rect 10806 49707 10871 49708
rect 10930 49707 10995 49708
rect 11054 49707 11119 49708
rect 11178 49707 11243 49708
rect 11302 49707 11367 49708
rect 10187 49652 10254 49707
rect 10310 49652 10378 49707
rect 10434 49652 10502 49707
rect 10558 49652 10626 49707
rect 10682 49652 10750 49707
rect 10806 49652 10874 49707
rect 10930 49652 10998 49707
rect 11054 49652 11122 49707
rect 11178 49652 11246 49707
rect 11302 49652 11370 49707
rect 11426 49652 11494 49708
rect 11550 49652 11618 49708
rect 11674 49652 11742 49708
rect 11798 49652 11866 49708
rect 11922 49652 11990 49708
rect 12046 49652 12114 49708
rect 12170 49652 12237 49708
rect 10187 49635 12237 49652
rect 10187 49583 10251 49635
rect 10303 49583 10375 49635
rect 10427 49583 10499 49635
rect 10551 49583 10623 49635
rect 10675 49583 10747 49635
rect 10799 49583 10871 49635
rect 10923 49583 10995 49635
rect 11047 49583 11119 49635
rect 11171 49583 11243 49635
rect 11295 49583 11367 49635
rect 11419 49583 12237 49635
rect 10187 48825 12237 49583
rect 10187 48773 10251 48825
rect 10303 48773 10375 48825
rect 10427 48773 10499 48825
rect 10551 48773 10623 48825
rect 10675 48773 10747 48825
rect 10799 48773 10871 48825
rect 10923 48773 10995 48825
rect 11047 48773 11119 48825
rect 11171 48773 11243 48825
rect 11295 48773 11367 48825
rect 11419 48773 12237 48825
rect 10187 48701 12237 48773
rect 10187 48649 10251 48701
rect 10303 48649 10375 48701
rect 10427 48649 10499 48701
rect 10551 48649 10623 48701
rect 10675 48649 10747 48701
rect 10799 48649 10871 48701
rect 10923 48649 10995 48701
rect 11047 48649 11119 48701
rect 11171 48649 11243 48701
rect 11295 48649 11367 48701
rect 11419 48649 12237 48701
rect 10187 47988 12237 48649
rect 10187 47936 10256 47988
rect 10308 47936 10380 47988
rect 10432 47936 10504 47988
rect 10556 47936 10628 47988
rect 10680 47936 10752 47988
rect 10804 47936 10876 47988
rect 10928 47936 11000 47988
rect 11052 47936 11124 47988
rect 11176 47936 11248 47988
rect 11300 47936 11372 47988
rect 11424 47936 11496 47988
rect 11548 47936 11620 47988
rect 11672 47936 11744 47988
rect 11796 47936 11868 47988
rect 11920 47936 11992 47988
rect 12044 47936 12116 47988
rect 12168 47936 12237 47988
rect 10187 47864 12237 47936
rect 10187 47812 10256 47864
rect 10308 47812 10380 47864
rect 10432 47812 10504 47864
rect 10556 47812 10628 47864
rect 10680 47812 10752 47864
rect 10804 47812 10876 47864
rect 10928 47812 11000 47864
rect 11052 47812 11124 47864
rect 11176 47812 11248 47864
rect 11300 47812 11372 47864
rect 11424 47812 11496 47864
rect 11548 47812 11620 47864
rect 11672 47812 11744 47864
rect 11796 47812 11868 47864
rect 11920 47812 11992 47864
rect 12044 47812 12116 47864
rect 12168 47812 12237 47864
rect 10187 47748 12237 47812
rect 10187 47692 10254 47748
rect 10310 47692 10378 47748
rect 10434 47692 10502 47748
rect 10558 47692 10626 47748
rect 10682 47692 10750 47748
rect 10806 47692 10874 47748
rect 10930 47692 10998 47748
rect 11054 47692 11122 47748
rect 11178 47692 11246 47748
rect 11302 47692 11370 47748
rect 11426 47692 11494 47748
rect 11550 47692 11618 47748
rect 11674 47692 11742 47748
rect 11798 47692 11866 47748
rect 11922 47692 11990 47748
rect 12046 47692 12114 47748
rect 12170 47692 12237 47748
rect 10187 47688 10256 47692
rect 10308 47688 10380 47692
rect 10432 47688 10504 47692
rect 10556 47688 10628 47692
rect 10680 47688 10752 47692
rect 10804 47688 10876 47692
rect 10928 47688 11000 47692
rect 11052 47688 11124 47692
rect 11176 47688 11248 47692
rect 11300 47688 11372 47692
rect 11424 47688 11496 47692
rect 11548 47688 11620 47692
rect 11672 47688 11744 47692
rect 11796 47688 11868 47692
rect 11920 47688 11992 47692
rect 12044 47688 12116 47692
rect 12168 47688 12237 47692
rect 10187 47624 12237 47688
rect 10187 47568 10254 47624
rect 10310 47568 10378 47624
rect 10434 47568 10502 47624
rect 10558 47568 10626 47624
rect 10682 47568 10750 47624
rect 10806 47568 10874 47624
rect 10930 47568 10998 47624
rect 11054 47568 11122 47624
rect 11178 47568 11246 47624
rect 11302 47568 11370 47624
rect 11426 47568 11494 47624
rect 11550 47568 11618 47624
rect 11674 47568 11742 47624
rect 11798 47568 11866 47624
rect 11922 47568 11990 47624
rect 12046 47568 12114 47624
rect 12170 47568 12237 47624
rect 10187 47500 12237 47568
rect 10187 47444 10254 47500
rect 10310 47444 10378 47500
rect 10434 47444 10502 47500
rect 10558 47444 10626 47500
rect 10682 47444 10750 47500
rect 10806 47444 10874 47500
rect 10930 47444 10998 47500
rect 11054 47444 11122 47500
rect 11178 47444 11246 47500
rect 11302 47444 11370 47500
rect 11426 47444 11494 47500
rect 11550 47444 11618 47500
rect 11674 47444 11742 47500
rect 11798 47444 11866 47500
rect 11922 47444 11990 47500
rect 12046 47444 12114 47500
rect 12170 47444 12237 47500
rect 10187 47376 12237 47444
rect 10187 47320 10254 47376
rect 10310 47320 10378 47376
rect 10434 47320 10502 47376
rect 10558 47320 10626 47376
rect 10682 47320 10750 47376
rect 10806 47320 10874 47376
rect 10930 47320 10998 47376
rect 11054 47320 11122 47376
rect 11178 47320 11246 47376
rect 11302 47320 11370 47376
rect 11426 47320 11494 47376
rect 11550 47320 11618 47376
rect 11674 47320 11742 47376
rect 11798 47320 11866 47376
rect 11922 47320 11990 47376
rect 12046 47320 12114 47376
rect 12170 47320 12237 47376
rect 10187 47281 12237 47320
rect 12297 57225 12497 57278
rect 12297 57169 12307 57225
rect 12363 57169 12431 57225
rect 12487 57169 12497 57225
rect 12297 57108 12497 57169
rect 12297 57101 12317 57108
rect 12297 57045 12307 57101
rect 12369 57056 12425 57108
rect 12477 57101 12497 57108
rect 12363 57045 12431 57056
rect 12487 57045 12497 57101
rect 12297 56977 12497 57045
rect 12297 56921 12307 56977
rect 12363 56921 12431 56977
rect 12487 56921 12497 56977
rect 12297 56853 12497 56921
rect 12297 56797 12307 56853
rect 12363 56797 12431 56853
rect 12487 56797 12497 56853
rect 12297 56729 12497 56797
rect 12297 56673 12307 56729
rect 12363 56673 12431 56729
rect 12487 56673 12497 56729
rect 12297 56605 12497 56673
rect 12297 56549 12307 56605
rect 12363 56549 12431 56605
rect 12487 56549 12497 56605
rect 12297 56481 12497 56549
rect 12297 56425 12307 56481
rect 12363 56425 12431 56481
rect 12487 56425 12497 56481
rect 12297 56357 12497 56425
rect 12297 56301 12307 56357
rect 12363 56301 12431 56357
rect 12487 56301 12497 56357
rect 12297 56233 12497 56301
rect 12297 56177 12307 56233
rect 12363 56177 12431 56233
rect 12487 56177 12497 56233
rect 12297 56109 12497 56177
rect 12297 56053 12307 56109
rect 12363 56053 12431 56109
rect 12487 56053 12497 56109
rect 12297 54148 12497 56053
rect 12297 54092 12307 54148
rect 12363 54092 12431 54148
rect 12487 54092 12497 54148
rect 12297 54024 12497 54092
rect 12297 53968 12307 54024
rect 12363 53968 12431 54024
rect 12487 53968 12497 54024
rect 12297 53900 12497 53968
rect 12297 53844 12307 53900
rect 12363 53844 12431 53900
rect 12487 53844 12497 53900
rect 12297 53776 12497 53844
rect 12297 53720 12307 53776
rect 12363 53720 12431 53776
rect 12487 53720 12497 53776
rect 12297 53652 12497 53720
rect 12297 53596 12307 53652
rect 12363 53596 12431 53652
rect 12487 53596 12497 53652
rect 12297 53528 12497 53596
rect 12297 53472 12307 53528
rect 12363 53484 12431 53528
rect 12297 53432 12317 53472
rect 12369 53432 12425 53484
rect 12487 53472 12497 53528
rect 12477 53432 12497 53472
rect 12297 53404 12497 53432
rect 12297 53348 12307 53404
rect 12363 53376 12431 53404
rect 12297 53324 12317 53348
rect 12369 53324 12425 53376
rect 12487 53348 12497 53404
rect 12477 53324 12497 53348
rect 12297 53280 12497 53324
rect 12297 53224 12307 53280
rect 12363 53268 12431 53280
rect 12297 53216 12317 53224
rect 12369 53216 12425 53268
rect 12487 53224 12497 53280
rect 12477 53216 12497 53224
rect 12297 53156 12497 53216
rect 12297 53100 12307 53156
rect 12363 53100 12431 53156
rect 12487 53100 12497 53156
rect 12297 53032 12497 53100
rect 12297 52976 12307 53032
rect 12363 52976 12431 53032
rect 12487 52976 12497 53032
rect 12297 52908 12497 52976
rect 12297 52852 12307 52908
rect 12363 52852 12431 52908
rect 12487 52852 12497 52908
rect 12297 49348 12497 52852
rect 12297 49292 12307 49348
rect 12363 49292 12431 49348
rect 12487 49292 12497 49348
rect 12297 49224 12497 49292
rect 12297 49168 12307 49224
rect 12363 49168 12431 49224
rect 12487 49168 12497 49224
rect 12297 49100 12497 49168
rect 12297 49044 12307 49100
rect 12363 49044 12431 49100
rect 12487 49044 12497 49100
rect 12297 48976 12497 49044
rect 12297 48920 12307 48976
rect 12363 48920 12431 48976
rect 12487 48920 12497 48976
rect 12297 48852 12497 48920
rect 12297 48796 12307 48852
rect 12363 48796 12431 48852
rect 12487 48796 12497 48852
rect 12297 48728 12497 48796
rect 12297 48672 12307 48728
rect 12363 48672 12431 48728
rect 12487 48672 12497 48728
rect 12297 48604 12497 48672
rect 12297 48548 12307 48604
rect 12363 48548 12431 48604
rect 12487 48548 12497 48604
rect 12297 48480 12497 48548
rect 12297 48424 12307 48480
rect 12363 48424 12431 48480
rect 12487 48424 12497 48480
rect 12297 48356 12497 48424
rect 12297 48300 12307 48356
rect 12363 48300 12431 48356
rect 12487 48300 12497 48356
rect 12297 48232 12497 48300
rect 12297 48176 12307 48232
rect 12363 48176 12431 48232
rect 12487 48176 12497 48232
rect 12297 48108 12497 48176
rect 12297 48052 12307 48108
rect 12363 48052 12431 48108
rect 12487 48052 12497 48108
rect 12297 47281 12497 48052
rect 12817 56669 14717 57600
rect 12817 56617 13141 56669
rect 13193 56617 13265 56669
rect 13317 56617 13389 56669
rect 13441 56617 13513 56669
rect 13565 56617 13637 56669
rect 13689 56617 13761 56669
rect 13813 56617 13885 56669
rect 13937 56617 14009 56669
rect 14061 56617 14717 56669
rect 12817 56545 14717 56617
rect 12817 56493 13141 56545
rect 13193 56493 13265 56545
rect 13317 56493 13389 56545
rect 13441 56493 13513 56545
rect 13565 56493 13637 56545
rect 13689 56493 13761 56545
rect 13813 56493 13885 56545
rect 13937 56493 14009 56545
rect 14061 56493 14717 56545
rect 12817 56421 14717 56493
rect 12817 56369 13141 56421
rect 13193 56369 13265 56421
rect 13317 56369 13389 56421
rect 13441 56369 13513 56421
rect 13565 56369 13637 56421
rect 13689 56369 13761 56421
rect 13813 56369 13885 56421
rect 13937 56369 14009 56421
rect 14061 56369 14717 56421
rect 12817 56297 14717 56369
rect 12817 56245 13141 56297
rect 13193 56245 13265 56297
rect 13317 56245 13389 56297
rect 13441 56245 13513 56297
rect 13565 56245 13637 56297
rect 13689 56245 13761 56297
rect 13813 56245 13885 56297
rect 13937 56245 14009 56297
rect 14061 56245 14717 56297
rect 12817 56173 14717 56245
rect 12817 56121 13141 56173
rect 13193 56121 13265 56173
rect 13317 56121 13389 56173
rect 13441 56121 13513 56173
rect 13565 56121 13637 56173
rect 13689 56121 13761 56173
rect 13813 56121 13885 56173
rect 13937 56121 14009 56173
rect 14061 56121 14717 56173
rect 12817 56049 14717 56121
rect 12817 55997 13141 56049
rect 13193 55997 13265 56049
rect 13317 55997 13389 56049
rect 13441 55997 13513 56049
rect 13565 55997 13637 56049
rect 13689 55997 13761 56049
rect 13813 55997 13885 56049
rect 13937 55997 14009 56049
rect 14061 55997 14717 56049
rect 12817 55925 14717 55997
rect 12817 55873 13141 55925
rect 13193 55873 13265 55925
rect 13317 55873 13389 55925
rect 13441 55873 13513 55925
rect 13565 55873 13637 55925
rect 13689 55873 13761 55925
rect 13813 55873 13885 55925
rect 13937 55873 14009 55925
rect 14061 55873 14717 55925
rect 12817 55801 14717 55873
rect 12817 55749 13141 55801
rect 13193 55749 13265 55801
rect 13317 55749 13389 55801
rect 13441 55749 13513 55801
rect 13565 55749 13637 55801
rect 13689 55749 13761 55801
rect 13813 55749 13885 55801
rect 13937 55749 14009 55801
rect 14061 55749 14717 55801
rect 12817 55748 14717 55749
rect 12817 55692 12871 55748
rect 12927 55692 12995 55748
rect 13051 55692 13119 55748
rect 13175 55692 13243 55748
rect 13299 55692 13367 55748
rect 13423 55692 13491 55748
rect 13547 55692 13615 55748
rect 13671 55692 13739 55748
rect 13795 55692 13863 55748
rect 13919 55692 13987 55748
rect 14043 55692 14111 55748
rect 14167 55692 14235 55748
rect 14291 55692 14359 55748
rect 14415 55692 14483 55748
rect 14539 55692 14607 55748
rect 14663 55692 14717 55748
rect 12817 55677 14717 55692
rect 12817 55625 13141 55677
rect 13193 55625 13265 55677
rect 13317 55625 13389 55677
rect 13441 55625 13513 55677
rect 13565 55625 13637 55677
rect 13689 55625 13761 55677
rect 13813 55625 13885 55677
rect 13937 55625 14009 55677
rect 14061 55625 14717 55677
rect 12817 55624 14717 55625
rect 12817 55568 12871 55624
rect 12927 55568 12995 55624
rect 13051 55568 13119 55624
rect 13175 55568 13243 55624
rect 13299 55568 13367 55624
rect 13423 55568 13491 55624
rect 13547 55568 13615 55624
rect 13671 55568 13739 55624
rect 13795 55568 13863 55624
rect 13919 55568 13987 55624
rect 14043 55568 14111 55624
rect 14167 55568 14235 55624
rect 14291 55568 14359 55624
rect 14415 55568 14483 55624
rect 14539 55568 14607 55624
rect 14663 55568 14717 55624
rect 12817 55553 14717 55568
rect 12817 55501 13141 55553
rect 13193 55501 13265 55553
rect 13317 55501 13389 55553
rect 13441 55501 13513 55553
rect 13565 55501 13637 55553
rect 13689 55501 13761 55553
rect 13813 55501 13885 55553
rect 13937 55501 14009 55553
rect 14061 55501 14717 55553
rect 12817 55500 14717 55501
rect 12817 55444 12871 55500
rect 12927 55444 12995 55500
rect 13051 55444 13119 55500
rect 13175 55444 13243 55500
rect 13299 55444 13367 55500
rect 13423 55444 13491 55500
rect 13547 55444 13615 55500
rect 13671 55444 13739 55500
rect 13795 55444 13863 55500
rect 13919 55444 13987 55500
rect 14043 55444 14111 55500
rect 14167 55444 14235 55500
rect 14291 55444 14359 55500
rect 14415 55444 14483 55500
rect 14539 55444 14607 55500
rect 14663 55444 14717 55500
rect 12817 55429 14717 55444
rect 12817 55377 13141 55429
rect 13193 55377 13265 55429
rect 13317 55377 13389 55429
rect 13441 55377 13513 55429
rect 13565 55377 13637 55429
rect 13689 55377 13761 55429
rect 13813 55377 13885 55429
rect 13937 55377 14009 55429
rect 14061 55377 14717 55429
rect 12817 55376 14717 55377
rect 12817 55320 12871 55376
rect 12927 55320 12995 55376
rect 13051 55320 13119 55376
rect 13175 55320 13243 55376
rect 13299 55320 13367 55376
rect 13423 55320 13491 55376
rect 13547 55320 13615 55376
rect 13671 55320 13739 55376
rect 13795 55320 13863 55376
rect 13919 55320 13987 55376
rect 14043 55320 14111 55376
rect 14167 55320 14235 55376
rect 14291 55320 14359 55376
rect 14415 55320 14483 55376
rect 14539 55320 14607 55376
rect 14663 55320 14717 55376
rect 12817 55305 14717 55320
rect 12817 55253 13141 55305
rect 13193 55253 13265 55305
rect 13317 55253 13389 55305
rect 13441 55253 13513 55305
rect 13565 55253 13637 55305
rect 13689 55253 13761 55305
rect 13813 55253 13885 55305
rect 13937 55253 14009 55305
rect 14061 55253 14717 55305
rect 12817 55252 14717 55253
rect 12817 55196 12871 55252
rect 12927 55196 12995 55252
rect 13051 55196 13119 55252
rect 13175 55196 13243 55252
rect 13299 55196 13367 55252
rect 13423 55196 13491 55252
rect 13547 55196 13615 55252
rect 13671 55196 13739 55252
rect 13795 55196 13863 55252
rect 13919 55196 13987 55252
rect 14043 55196 14111 55252
rect 14167 55196 14235 55252
rect 14291 55196 14359 55252
rect 14415 55196 14483 55252
rect 14539 55196 14607 55252
rect 14663 55196 14717 55252
rect 12817 55181 14717 55196
rect 12817 55129 13141 55181
rect 13193 55129 13265 55181
rect 13317 55129 13389 55181
rect 13441 55129 13513 55181
rect 13565 55129 13637 55181
rect 13689 55129 13761 55181
rect 13813 55129 13885 55181
rect 13937 55129 14009 55181
rect 14061 55129 14717 55181
rect 12817 55128 14717 55129
rect 12817 55072 12871 55128
rect 12927 55072 12995 55128
rect 13051 55072 13119 55128
rect 13175 55072 13243 55128
rect 13299 55072 13367 55128
rect 13423 55072 13491 55128
rect 13547 55072 13615 55128
rect 13671 55072 13739 55128
rect 13795 55072 13863 55128
rect 13919 55072 13987 55128
rect 14043 55072 14111 55128
rect 14167 55072 14235 55128
rect 14291 55072 14359 55128
rect 14415 55072 14483 55128
rect 14539 55072 14607 55128
rect 14663 55072 14717 55128
rect 12817 55057 14717 55072
rect 12817 55005 13141 55057
rect 13193 55005 13265 55057
rect 13317 55005 13389 55057
rect 13441 55005 13513 55057
rect 13565 55005 13637 55057
rect 13689 55005 13761 55057
rect 13813 55005 13885 55057
rect 13937 55005 14009 55057
rect 14061 55005 14717 55057
rect 12817 55004 14717 55005
rect 12817 54948 12871 55004
rect 12927 54948 12995 55004
rect 13051 54948 13119 55004
rect 13175 54948 13243 55004
rect 13299 54948 13367 55004
rect 13423 54948 13491 55004
rect 13547 54948 13615 55004
rect 13671 54948 13739 55004
rect 13795 54948 13863 55004
rect 13919 54948 13987 55004
rect 14043 54948 14111 55004
rect 14167 54948 14235 55004
rect 14291 54948 14359 55004
rect 14415 54948 14483 55004
rect 14539 54948 14607 55004
rect 14663 54948 14717 55004
rect 12817 54933 14717 54948
rect 12817 54881 13141 54933
rect 13193 54881 13265 54933
rect 13317 54881 13389 54933
rect 13441 54881 13513 54933
rect 13565 54881 13637 54933
rect 13689 54881 13761 54933
rect 13813 54881 13885 54933
rect 13937 54881 14009 54933
rect 14061 54881 14717 54933
rect 12817 54880 14717 54881
rect 12817 54824 12871 54880
rect 12927 54824 12995 54880
rect 13051 54824 13119 54880
rect 13175 54824 13243 54880
rect 13299 54824 13367 54880
rect 13423 54824 13491 54880
rect 13547 54824 13615 54880
rect 13671 54824 13739 54880
rect 13795 54824 13863 54880
rect 13919 54824 13987 54880
rect 14043 54824 14111 54880
rect 14167 54824 14235 54880
rect 14291 54824 14359 54880
rect 14415 54824 14483 54880
rect 14539 54824 14607 54880
rect 14663 54824 14717 54880
rect 12817 54809 14717 54824
rect 12817 54757 13141 54809
rect 13193 54757 13265 54809
rect 13317 54757 13389 54809
rect 13441 54757 13513 54809
rect 13565 54757 13637 54809
rect 13689 54757 13761 54809
rect 13813 54757 13885 54809
rect 13937 54757 14009 54809
rect 14061 54757 14717 54809
rect 12817 54756 14717 54757
rect 12817 54700 12871 54756
rect 12927 54700 12995 54756
rect 13051 54700 13119 54756
rect 13175 54700 13243 54756
rect 13299 54700 13367 54756
rect 13423 54700 13491 54756
rect 13547 54700 13615 54756
rect 13671 54700 13739 54756
rect 13795 54700 13863 54756
rect 13919 54700 13987 54756
rect 14043 54700 14111 54756
rect 14167 54700 14235 54756
rect 14291 54700 14359 54756
rect 14415 54700 14483 54756
rect 14539 54700 14607 54756
rect 14663 54700 14717 54756
rect 12817 54685 14717 54700
rect 12817 54633 13141 54685
rect 13193 54633 13265 54685
rect 13317 54633 13389 54685
rect 13441 54633 13513 54685
rect 13565 54633 13637 54685
rect 13689 54633 13761 54685
rect 13813 54633 13885 54685
rect 13937 54633 14009 54685
rect 14061 54633 14717 54685
rect 12817 54632 14717 54633
rect 12817 54576 12871 54632
rect 12927 54576 12995 54632
rect 13051 54576 13119 54632
rect 13175 54576 13243 54632
rect 13299 54576 13367 54632
rect 13423 54576 13491 54632
rect 13547 54576 13615 54632
rect 13671 54576 13739 54632
rect 13795 54576 13863 54632
rect 13919 54576 13987 54632
rect 14043 54576 14111 54632
rect 14167 54576 14235 54632
rect 14291 54576 14359 54632
rect 14415 54576 14483 54632
rect 14539 54576 14607 54632
rect 14663 54576 14717 54632
rect 12817 54561 14717 54576
rect 12817 54509 13141 54561
rect 13193 54509 13265 54561
rect 13317 54509 13389 54561
rect 13441 54509 13513 54561
rect 13565 54509 13637 54561
rect 13689 54509 13761 54561
rect 13813 54509 13885 54561
rect 13937 54509 14009 54561
rect 14061 54509 14717 54561
rect 12817 54508 14717 54509
rect 12817 54452 12871 54508
rect 12927 54452 12995 54508
rect 13051 54452 13119 54508
rect 13175 54452 13243 54508
rect 13299 54452 13367 54508
rect 13423 54452 13491 54508
rect 13547 54452 13615 54508
rect 13671 54452 13739 54508
rect 13795 54452 13863 54508
rect 13919 54452 13987 54508
rect 14043 54452 14111 54508
rect 14167 54452 14235 54508
rect 14291 54452 14359 54508
rect 14415 54452 14483 54508
rect 14539 54452 14607 54508
rect 14663 54452 14717 54508
rect 12817 54437 14717 54452
rect 12817 54385 13141 54437
rect 13193 54385 13265 54437
rect 13317 54385 13389 54437
rect 13441 54385 13513 54437
rect 13565 54385 13637 54437
rect 13689 54385 13761 54437
rect 13813 54385 13885 54437
rect 13937 54385 14009 54437
rect 14061 54385 14717 54437
rect 12817 54313 14717 54385
rect 12817 54261 13141 54313
rect 13193 54261 13265 54313
rect 13317 54261 13389 54313
rect 13441 54261 13513 54313
rect 13565 54261 13637 54313
rect 13689 54261 13761 54313
rect 13813 54261 13885 54313
rect 13937 54261 14009 54313
rect 14061 54261 14717 54313
rect 12817 54189 14717 54261
rect 12817 54137 13141 54189
rect 13193 54137 13265 54189
rect 13317 54137 13389 54189
rect 13441 54137 13513 54189
rect 13565 54137 13637 54189
rect 13689 54137 13761 54189
rect 13813 54137 13885 54189
rect 13937 54137 14009 54189
rect 14061 54137 14717 54189
rect 12817 54065 14717 54137
rect 12817 54013 13141 54065
rect 13193 54013 13265 54065
rect 13317 54013 13389 54065
rect 13441 54013 13513 54065
rect 13565 54013 13637 54065
rect 13689 54013 13761 54065
rect 13813 54013 13885 54065
rect 13937 54013 14009 54065
rect 14061 54013 14717 54065
rect 12817 53941 14717 54013
rect 12817 53889 13141 53941
rect 13193 53889 13265 53941
rect 13317 53889 13389 53941
rect 13441 53889 13513 53941
rect 13565 53889 13637 53941
rect 13689 53889 13761 53941
rect 13813 53889 13885 53941
rect 13937 53889 14009 53941
rect 14061 53889 14717 53941
rect 12817 53817 14717 53889
rect 12817 53765 13141 53817
rect 13193 53765 13265 53817
rect 13317 53765 13389 53817
rect 13441 53765 13513 53817
rect 13565 53765 13637 53817
rect 13689 53765 13761 53817
rect 13813 53765 13885 53817
rect 13937 53765 14009 53817
rect 14061 53765 14717 53817
rect 12817 53693 14717 53765
rect 12817 53641 13141 53693
rect 13193 53641 13265 53693
rect 13317 53641 13389 53693
rect 13441 53641 13513 53693
rect 13565 53641 13637 53693
rect 13689 53641 13761 53693
rect 13813 53641 13885 53693
rect 13937 53641 14009 53693
rect 14061 53641 14717 53693
rect 12817 50948 14717 53641
rect 14892 52576 14989 52600
rect 14892 51224 14902 52576
rect 14958 51224 14989 52576
rect 14892 51200 14989 51224
rect 12817 50892 12871 50948
rect 12927 50892 12995 50948
rect 13051 50892 13119 50948
rect 13175 50892 13243 50948
rect 13299 50892 13367 50948
rect 13423 50892 13491 50948
rect 13547 50892 13615 50948
rect 13671 50892 13739 50948
rect 13795 50892 13863 50948
rect 13919 50892 13987 50948
rect 14043 50892 14111 50948
rect 14167 50892 14235 50948
rect 14291 50892 14359 50948
rect 14415 50892 14483 50948
rect 14539 50892 14607 50948
rect 14663 50892 14717 50948
rect 12817 50824 14717 50892
rect 12817 50768 12871 50824
rect 12927 50768 12995 50824
rect 13051 50768 13119 50824
rect 13175 50768 13243 50824
rect 13299 50768 13367 50824
rect 13423 50768 13491 50824
rect 13547 50768 13615 50824
rect 13671 50768 13739 50824
rect 13795 50768 13863 50824
rect 13919 50768 13987 50824
rect 14043 50768 14111 50824
rect 14167 50768 14235 50824
rect 14291 50768 14359 50824
rect 14415 50768 14483 50824
rect 14539 50768 14607 50824
rect 14663 50768 14717 50824
rect 12817 50700 14717 50768
rect 12817 50644 12871 50700
rect 12927 50644 12995 50700
rect 13051 50644 13119 50700
rect 13175 50644 13243 50700
rect 13299 50644 13367 50700
rect 13423 50644 13491 50700
rect 13547 50644 13615 50700
rect 13671 50644 13739 50700
rect 13795 50644 13863 50700
rect 13919 50644 13987 50700
rect 14043 50644 14111 50700
rect 14167 50644 14235 50700
rect 14291 50644 14359 50700
rect 14415 50644 14483 50700
rect 14539 50644 14607 50700
rect 14663 50644 14717 50700
rect 12817 50576 14717 50644
rect 12817 50520 12871 50576
rect 12927 50520 12995 50576
rect 13051 50520 13119 50576
rect 13175 50520 13243 50576
rect 13299 50520 13367 50576
rect 13423 50520 13491 50576
rect 13547 50520 13615 50576
rect 13671 50520 13739 50576
rect 13795 50520 13863 50576
rect 13919 50520 13987 50576
rect 14043 50520 14111 50576
rect 14167 50520 14235 50576
rect 14291 50520 14359 50576
rect 14415 50520 14483 50576
rect 14539 50520 14607 50576
rect 14663 50520 14717 50576
rect 12817 50452 14717 50520
rect 12817 50396 12871 50452
rect 12927 50396 12995 50452
rect 13051 50396 13119 50452
rect 13175 50396 13243 50452
rect 13299 50396 13367 50452
rect 13423 50396 13491 50452
rect 13547 50396 13615 50452
rect 13671 50396 13739 50452
rect 13795 50396 13863 50452
rect 13919 50396 13987 50452
rect 14043 50396 14111 50452
rect 14167 50396 14235 50452
rect 14291 50396 14359 50452
rect 14415 50396 14483 50452
rect 14539 50396 14607 50452
rect 14663 50396 14717 50452
rect 12817 50328 14717 50396
rect 12817 50272 12871 50328
rect 12927 50272 12995 50328
rect 13051 50272 13119 50328
rect 13175 50272 13243 50328
rect 13299 50272 13367 50328
rect 13423 50272 13491 50328
rect 13547 50272 13615 50328
rect 13671 50272 13739 50328
rect 13795 50272 13863 50328
rect 13919 50272 13987 50328
rect 14043 50272 14111 50328
rect 14167 50272 14235 50328
rect 14291 50272 14359 50328
rect 14415 50272 14483 50328
rect 14539 50272 14607 50328
rect 14663 50272 14717 50328
rect 12817 50204 14717 50272
rect 12817 50148 12871 50204
rect 12927 50148 12995 50204
rect 13051 50148 13119 50204
rect 13175 50148 13243 50204
rect 13299 50148 13367 50204
rect 13423 50148 13491 50204
rect 13547 50148 13615 50204
rect 13671 50148 13739 50204
rect 13795 50148 13863 50204
rect 13919 50148 13987 50204
rect 14043 50148 14111 50204
rect 14167 50148 14235 50204
rect 14291 50148 14359 50204
rect 14415 50148 14483 50204
rect 14539 50148 14607 50204
rect 14663 50148 14717 50204
rect 12817 50080 14717 50148
rect 12817 50024 12871 50080
rect 12927 50024 12995 50080
rect 13051 50024 13119 50080
rect 13175 50024 13243 50080
rect 13299 50024 13367 50080
rect 13423 50024 13491 50080
rect 13547 50024 13615 50080
rect 13671 50024 13739 50080
rect 13795 50024 13863 50080
rect 13919 50024 13987 50080
rect 14043 50024 14111 50080
rect 14167 50024 14235 50080
rect 14291 50024 14359 50080
rect 14415 50024 14483 50080
rect 14539 50024 14607 50080
rect 14663 50024 14717 50080
rect 12817 49956 14717 50024
rect 12817 49900 12871 49956
rect 12927 49900 12995 49956
rect 13051 49900 13119 49956
rect 13175 49900 13243 49956
rect 13299 49900 13367 49956
rect 13423 49900 13491 49956
rect 13547 49900 13615 49956
rect 13671 49900 13739 49956
rect 13795 49900 13863 49956
rect 13919 49900 13987 49956
rect 14043 49900 14111 49956
rect 14167 49900 14235 49956
rect 14291 49900 14359 49956
rect 14415 49900 14483 49956
rect 14539 49900 14607 49956
rect 14663 49900 14717 49956
rect 12817 49832 14717 49900
rect 12817 49776 12871 49832
rect 12927 49776 12995 49832
rect 13051 49776 13119 49832
rect 13175 49776 13243 49832
rect 13299 49776 13367 49832
rect 13423 49776 13491 49832
rect 13547 49776 13615 49832
rect 13671 49776 13739 49832
rect 13795 49776 13863 49832
rect 13919 49776 13987 49832
rect 14043 49776 14111 49832
rect 14167 49776 14235 49832
rect 14291 49776 14359 49832
rect 14415 49776 14483 49832
rect 14539 49776 14607 49832
rect 14663 49776 14717 49832
rect 12817 49708 14717 49776
rect 12817 49652 12871 49708
rect 12927 49652 12995 49708
rect 13051 49652 13119 49708
rect 13175 49652 13243 49708
rect 13299 49652 13367 49708
rect 13423 49652 13491 49708
rect 13547 49652 13615 49708
rect 13671 49652 13739 49708
rect 13795 49652 13863 49708
rect 13919 49652 13987 49708
rect 14043 49652 14111 49708
rect 14167 49652 14235 49708
rect 14291 49652 14359 49708
rect 14415 49652 14483 49708
rect 14539 49652 14607 49708
rect 14663 49652 14717 49708
rect 12817 47748 14717 49652
rect 12817 47692 12871 47748
rect 12927 47692 12995 47748
rect 13051 47692 13119 47748
rect 13175 47692 13243 47748
rect 13299 47692 13367 47748
rect 13423 47692 13491 47748
rect 13547 47692 13615 47748
rect 13671 47692 13739 47748
rect 13795 47692 13863 47748
rect 13919 47692 13987 47748
rect 14043 47692 14111 47748
rect 14167 47692 14235 47748
rect 14291 47692 14359 47748
rect 14415 47692 14483 47748
rect 14539 47692 14607 47748
rect 14663 47692 14717 47748
rect 12817 47624 14717 47692
rect 12817 47568 12871 47624
rect 12927 47568 12995 47624
rect 13051 47568 13119 47624
rect 13175 47568 13243 47624
rect 13299 47568 13367 47624
rect 13423 47568 13491 47624
rect 13547 47568 13615 47624
rect 13671 47568 13739 47624
rect 13795 47568 13863 47624
rect 13919 47568 13987 47624
rect 14043 47568 14111 47624
rect 14167 47568 14235 47624
rect 14291 47568 14359 47624
rect 14415 47568 14483 47624
rect 14539 47568 14607 47624
rect 14663 47568 14717 47624
rect 12817 47500 14717 47568
rect 12817 47444 12871 47500
rect 12927 47444 12995 47500
rect 13051 47444 13119 47500
rect 13175 47444 13243 47500
rect 13299 47444 13367 47500
rect 13423 47444 13491 47500
rect 13547 47444 13615 47500
rect 13671 47444 13739 47500
rect 13795 47444 13863 47500
rect 13919 47444 13987 47500
rect 14043 47444 14111 47500
rect 14167 47444 14235 47500
rect 14291 47444 14359 47500
rect 14415 47444 14483 47500
rect 14539 47444 14607 47500
rect 14663 47444 14717 47500
rect 12817 47376 14717 47444
rect 12817 47320 12871 47376
rect 12927 47320 12995 47376
rect 13051 47320 13119 47376
rect 13175 47320 13243 47376
rect 13299 47320 13367 47376
rect 13423 47320 13491 47376
rect 13547 47320 13615 47376
rect 13671 47320 13739 47376
rect 13795 47320 13863 47376
rect 13919 47320 13987 47376
rect 14043 47320 14111 47376
rect 14167 47320 14235 47376
rect 14291 47320 14359 47376
rect 14415 47320 14483 47376
rect 14539 47320 14607 47376
rect 14663 47320 14717 47376
rect 12817 47281 14717 47320
rect 2798 47252 4734 47281
rect 2798 47196 2808 47252
rect 2864 47196 2932 47252
rect 2988 47196 3056 47252
rect 3112 47196 3180 47252
rect 3236 47196 3304 47252
rect 3360 47196 3428 47252
rect 3484 47196 3552 47252
rect 3608 47196 3676 47252
rect 3732 47196 3800 47252
rect 3856 47196 3924 47252
rect 3980 47196 4048 47252
rect 4104 47196 4172 47252
rect 4228 47196 4296 47252
rect 4352 47196 4420 47252
rect 4476 47196 4544 47252
rect 4600 47196 4668 47252
rect 4724 47196 4734 47252
rect 2798 47128 4734 47196
rect 2798 47072 2808 47128
rect 2864 47072 2932 47128
rect 2988 47072 3056 47128
rect 3112 47072 3180 47128
rect 3236 47072 3304 47128
rect 3360 47072 3428 47128
rect 3484 47072 3552 47128
rect 3608 47072 3676 47128
rect 3732 47072 3800 47128
rect 3856 47072 3924 47128
rect 3980 47072 4048 47128
rect 4104 47072 4172 47128
rect 4228 47072 4296 47128
rect 4352 47072 4420 47128
rect 4476 47072 4544 47128
rect 4600 47072 4668 47128
rect 4724 47072 4734 47128
rect 2798 47004 4734 47072
rect 2798 46948 2808 47004
rect 2864 46948 2932 47004
rect 2988 46948 3056 47004
rect 3112 46948 3180 47004
rect 3236 46948 3304 47004
rect 3360 46948 3428 47004
rect 3484 46948 3552 47004
rect 3608 46948 3676 47004
rect 3732 46948 3800 47004
rect 3856 46948 3924 47004
rect 3980 46948 4048 47004
rect 4104 46948 4172 47004
rect 4228 46948 4296 47004
rect 4352 46948 4420 47004
rect 4476 46948 4544 47004
rect 4600 46948 4668 47004
rect 4724 46948 4734 47004
rect 2798 46880 4734 46948
rect 2798 46824 2808 46880
rect 2864 46824 2932 46880
rect 2988 46824 3056 46880
rect 3112 46824 3180 46880
rect 3236 46824 3304 46880
rect 3360 46824 3428 46880
rect 3484 46824 3552 46880
rect 3608 46824 3676 46880
rect 3732 46824 3800 46880
rect 3856 46824 3924 46880
rect 3980 46824 4048 46880
rect 4104 46824 4172 46880
rect 4228 46824 4296 46880
rect 4352 46824 4420 46880
rect 4476 46824 4544 46880
rect 4600 46824 4668 46880
rect 4724 46824 4734 46880
rect 2798 46756 4734 46824
rect 2798 46700 2808 46756
rect 2864 46700 2932 46756
rect 2988 46700 3056 46756
rect 3112 46700 3180 46756
rect 3236 46700 3304 46756
rect 3360 46700 3428 46756
rect 3484 46700 3552 46756
rect 3608 46700 3676 46756
rect 3732 46700 3800 46756
rect 3856 46700 3924 46756
rect 3980 46700 4048 46756
rect 4104 46700 4172 46756
rect 4228 46700 4296 46756
rect 4352 46700 4420 46756
rect 4476 46700 4544 46756
rect 4600 46700 4668 46756
rect 4724 46700 4734 46756
rect 2798 46632 4734 46700
rect 2798 46576 2808 46632
rect 2864 46576 2932 46632
rect 2988 46576 3056 46632
rect 3112 46576 3180 46632
rect 3236 46576 3304 46632
rect 3360 46576 3428 46632
rect 3484 46576 3552 46632
rect 3608 46576 3676 46632
rect 3732 46576 3800 46632
rect 3856 46576 3924 46632
rect 3980 46576 4048 46632
rect 4104 46576 4172 46632
rect 4228 46576 4296 46632
rect 4352 46576 4420 46632
rect 4476 46576 4544 46632
rect 4600 46576 4668 46632
rect 4724 46576 4734 46632
rect 2798 46508 4734 46576
rect 2798 46452 2808 46508
rect 2864 46452 2932 46508
rect 2988 46452 3056 46508
rect 3112 46452 3180 46508
rect 3236 46452 3304 46508
rect 3360 46452 3428 46508
rect 3484 46452 3552 46508
rect 3608 46452 3676 46508
rect 3732 46452 3800 46508
rect 3856 46452 3924 46508
rect 3980 46452 4048 46508
rect 4104 46452 4172 46508
rect 4228 46452 4296 46508
rect 4352 46452 4420 46508
rect 4476 46452 4544 46508
rect 4600 46452 4668 46508
rect 4724 46452 4734 46508
rect 2798 46442 4734 46452
rect 5168 47252 7104 47281
rect 5168 47196 5178 47252
rect 5234 47196 5302 47252
rect 5358 47196 5426 47252
rect 5482 47196 5550 47252
rect 5606 47196 5674 47252
rect 5730 47196 5798 47252
rect 5854 47196 5922 47252
rect 5978 47196 6046 47252
rect 6102 47196 6170 47252
rect 6226 47196 6294 47252
rect 6350 47196 6418 47252
rect 6474 47196 6542 47252
rect 6598 47196 6666 47252
rect 6722 47196 6790 47252
rect 6846 47196 6914 47252
rect 6970 47196 7038 47252
rect 7094 47196 7104 47252
rect 5168 47128 7104 47196
rect 5168 47072 5178 47128
rect 5234 47072 5302 47128
rect 5358 47072 5426 47128
rect 5482 47072 5550 47128
rect 5606 47072 5674 47128
rect 5730 47072 5798 47128
rect 5854 47072 5922 47128
rect 5978 47072 6046 47128
rect 6102 47072 6170 47128
rect 6226 47072 6294 47128
rect 6350 47072 6418 47128
rect 6474 47072 6542 47128
rect 6598 47072 6666 47128
rect 6722 47072 6790 47128
rect 6846 47072 6914 47128
rect 6970 47072 7038 47128
rect 7094 47072 7104 47128
rect 5168 47004 7104 47072
rect 5168 46948 5178 47004
rect 5234 46948 5302 47004
rect 5358 46948 5426 47004
rect 5482 46948 5550 47004
rect 5606 46948 5674 47004
rect 5730 46948 5798 47004
rect 5854 46948 5922 47004
rect 5978 46948 6046 47004
rect 6102 46948 6170 47004
rect 6226 46948 6294 47004
rect 6350 46948 6418 47004
rect 6474 46948 6542 47004
rect 6598 46948 6666 47004
rect 6722 46948 6790 47004
rect 6846 46948 6914 47004
rect 6970 46948 7038 47004
rect 7094 46948 7104 47004
rect 5168 46880 7104 46948
rect 5168 46824 5178 46880
rect 5234 46824 5302 46880
rect 5358 46824 5426 46880
rect 5482 46824 5550 46880
rect 5606 46824 5674 46880
rect 5730 46824 5798 46880
rect 5854 46824 5922 46880
rect 5978 46824 6046 46880
rect 6102 46824 6170 46880
rect 6226 46824 6294 46880
rect 6350 46824 6418 46880
rect 6474 46824 6542 46880
rect 6598 46824 6666 46880
rect 6722 46824 6790 46880
rect 6846 46824 6914 46880
rect 6970 46824 7038 46880
rect 7094 46824 7104 46880
rect 5168 46756 7104 46824
rect 5168 46700 5178 46756
rect 5234 46700 5302 46756
rect 5358 46700 5426 46756
rect 5482 46700 5550 46756
rect 5606 46700 5674 46756
rect 5730 46700 5798 46756
rect 5854 46700 5922 46756
rect 5978 46700 6046 46756
rect 6102 46700 6170 46756
rect 6226 46700 6294 46756
rect 6350 46700 6418 46756
rect 6474 46700 6542 46756
rect 6598 46700 6666 46756
rect 6722 46700 6790 46756
rect 6846 46700 6914 46756
rect 6970 46700 7038 46756
rect 7094 46700 7104 46756
rect 5168 46632 7104 46700
rect 5168 46576 5178 46632
rect 5234 46576 5302 46632
rect 5358 46576 5426 46632
rect 5482 46576 5550 46632
rect 5606 46576 5674 46632
rect 5730 46576 5798 46632
rect 5854 46576 5922 46632
rect 5978 46576 6046 46632
rect 6102 46576 6170 46632
rect 6226 46576 6294 46632
rect 6350 46576 6418 46632
rect 6474 46576 6542 46632
rect 6598 46576 6666 46632
rect 6722 46576 6790 46632
rect 6846 46576 6914 46632
rect 6970 46576 7038 46632
rect 7094 46576 7104 46632
rect 5168 46508 7104 46576
rect 5168 46452 5178 46508
rect 5234 46452 5302 46508
rect 5358 46452 5426 46508
rect 5482 46452 5550 46508
rect 5606 46452 5674 46508
rect 5730 46452 5798 46508
rect 5854 46452 5922 46508
rect 5978 46452 6046 46508
rect 6102 46452 6170 46508
rect 6226 46452 6294 46508
rect 6350 46452 6418 46508
rect 6474 46452 6542 46508
rect 6598 46452 6666 46508
rect 6722 46452 6790 46508
rect 6846 46452 6914 46508
rect 6970 46452 7038 46508
rect 7094 46452 7104 46508
rect 5168 46442 7104 46452
rect 7874 47252 9810 47281
rect 7874 47196 7884 47252
rect 7940 47196 8008 47252
rect 8064 47196 8132 47252
rect 8188 47196 8256 47252
rect 8312 47196 8380 47252
rect 8436 47196 8504 47252
rect 8560 47196 8628 47252
rect 8684 47196 8752 47252
rect 8808 47196 8876 47252
rect 8932 47196 9000 47252
rect 9056 47196 9124 47252
rect 9180 47196 9248 47252
rect 9304 47196 9372 47252
rect 9428 47196 9496 47252
rect 9552 47196 9620 47252
rect 9676 47196 9744 47252
rect 9800 47196 9810 47252
rect 7874 47128 9810 47196
rect 7874 47072 7884 47128
rect 7940 47072 8008 47128
rect 8064 47072 8132 47128
rect 8188 47072 8256 47128
rect 8312 47072 8380 47128
rect 8436 47072 8504 47128
rect 8560 47072 8628 47128
rect 8684 47072 8752 47128
rect 8808 47072 8876 47128
rect 8932 47072 9000 47128
rect 9056 47072 9124 47128
rect 9180 47072 9248 47128
rect 9304 47072 9372 47128
rect 9428 47072 9496 47128
rect 9552 47072 9620 47128
rect 9676 47072 9744 47128
rect 9800 47072 9810 47128
rect 7874 47004 9810 47072
rect 7874 46948 7884 47004
rect 7940 46948 8008 47004
rect 8064 46948 8132 47004
rect 8188 46948 8256 47004
rect 8312 46948 8380 47004
rect 8436 46948 8504 47004
rect 8560 46948 8628 47004
rect 8684 46948 8752 47004
rect 8808 46948 8876 47004
rect 8932 46948 9000 47004
rect 9056 46948 9124 47004
rect 9180 46948 9248 47004
rect 9304 46948 9372 47004
rect 9428 46948 9496 47004
rect 9552 46948 9620 47004
rect 9676 46948 9744 47004
rect 9800 46948 9810 47004
rect 7874 46880 9810 46948
rect 7874 46824 7884 46880
rect 7940 46824 8008 46880
rect 8064 46824 8132 46880
rect 8188 46824 8256 46880
rect 8312 46824 8380 46880
rect 8436 46824 8504 46880
rect 8560 46824 8628 46880
rect 8684 46824 8752 46880
rect 8808 46824 8876 46880
rect 8932 46824 9000 46880
rect 9056 46824 9124 46880
rect 9180 46824 9248 46880
rect 9304 46824 9372 46880
rect 9428 46824 9496 46880
rect 9552 46824 9620 46880
rect 9676 46824 9744 46880
rect 9800 46824 9810 46880
rect 7874 46756 9810 46824
rect 7874 46700 7884 46756
rect 7940 46700 8008 46756
rect 8064 46700 8132 46756
rect 8188 46700 8256 46756
rect 8312 46700 8380 46756
rect 8436 46700 8504 46756
rect 8560 46700 8628 46756
rect 8684 46700 8752 46756
rect 8808 46700 8876 46756
rect 8932 46700 9000 46756
rect 9056 46700 9124 46756
rect 9180 46700 9248 46756
rect 9304 46700 9372 46756
rect 9428 46700 9496 46756
rect 9552 46700 9620 46756
rect 9676 46700 9744 46756
rect 9800 46700 9810 46756
rect 7874 46632 9810 46700
rect 7874 46576 7884 46632
rect 7940 46576 8008 46632
rect 8064 46576 8132 46632
rect 8188 46576 8256 46632
rect 8312 46576 8380 46632
rect 8436 46576 8504 46632
rect 8560 46576 8628 46632
rect 8684 46576 8752 46632
rect 8808 46576 8876 46632
rect 8932 46576 9000 46632
rect 9056 46576 9124 46632
rect 9180 46576 9248 46632
rect 9304 46576 9372 46632
rect 9428 46576 9496 46632
rect 9552 46576 9620 46632
rect 9676 46576 9744 46632
rect 9800 46576 9810 46632
rect 7874 46508 9810 46576
rect 7874 46452 7884 46508
rect 7940 46452 8008 46508
rect 8064 46452 8132 46508
rect 8188 46452 8256 46508
rect 8312 46452 8380 46508
rect 8436 46452 8504 46508
rect 8560 46452 8628 46508
rect 8684 46452 8752 46508
rect 8808 46452 8876 46508
rect 8932 46452 9000 46508
rect 9056 46452 9124 46508
rect 9180 46452 9248 46508
rect 9304 46452 9372 46508
rect 9428 46452 9496 46508
rect 9552 46452 9620 46508
rect 9676 46452 9744 46508
rect 9800 46452 9810 46508
rect 7874 46442 9810 46452
rect 10244 47252 12180 47281
rect 10244 47196 10254 47252
rect 10310 47196 10378 47252
rect 10434 47196 10502 47252
rect 10558 47196 10626 47252
rect 10682 47196 10750 47252
rect 10806 47196 10874 47252
rect 10930 47196 10998 47252
rect 11054 47196 11122 47252
rect 11178 47196 11246 47252
rect 11302 47196 11370 47252
rect 11426 47196 11494 47252
rect 11550 47196 11618 47252
rect 11674 47196 11742 47252
rect 11798 47196 11866 47252
rect 11922 47196 11990 47252
rect 12046 47196 12114 47252
rect 12170 47196 12180 47252
rect 10244 47128 12180 47196
rect 10244 47072 10254 47128
rect 10310 47072 10378 47128
rect 10434 47072 10502 47128
rect 10558 47072 10626 47128
rect 10682 47072 10750 47128
rect 10806 47072 10874 47128
rect 10930 47072 10998 47128
rect 11054 47072 11122 47128
rect 11178 47072 11246 47128
rect 11302 47072 11370 47128
rect 11426 47072 11494 47128
rect 11550 47072 11618 47128
rect 11674 47072 11742 47128
rect 11798 47072 11866 47128
rect 11922 47072 11990 47128
rect 12046 47072 12114 47128
rect 12170 47072 12180 47128
rect 10244 47004 12180 47072
rect 10244 46948 10254 47004
rect 10310 46948 10378 47004
rect 10434 46948 10502 47004
rect 10558 46948 10626 47004
rect 10682 46948 10750 47004
rect 10806 46948 10874 47004
rect 10930 46948 10998 47004
rect 11054 46948 11122 47004
rect 11178 46948 11246 47004
rect 11302 46948 11370 47004
rect 11426 46948 11494 47004
rect 11550 46948 11618 47004
rect 11674 46948 11742 47004
rect 11798 46948 11866 47004
rect 11922 46948 11990 47004
rect 12046 46948 12114 47004
rect 12170 46948 12180 47004
rect 10244 46880 12180 46948
rect 10244 46824 10254 46880
rect 10310 46824 10378 46880
rect 10434 46824 10502 46880
rect 10558 46824 10626 46880
rect 10682 46824 10750 46880
rect 10806 46824 10874 46880
rect 10930 46824 10998 46880
rect 11054 46824 11122 46880
rect 11178 46824 11246 46880
rect 11302 46824 11370 46880
rect 11426 46824 11494 46880
rect 11550 46824 11618 46880
rect 11674 46824 11742 46880
rect 11798 46824 11866 46880
rect 11922 46824 11990 46880
rect 12046 46824 12114 46880
rect 12170 46824 12180 46880
rect 10244 46756 12180 46824
rect 10244 46700 10254 46756
rect 10310 46700 10378 46756
rect 10434 46700 10502 46756
rect 10558 46700 10626 46756
rect 10682 46700 10750 46756
rect 10806 46700 10874 46756
rect 10930 46700 10998 46756
rect 11054 46700 11122 46756
rect 11178 46700 11246 46756
rect 11302 46700 11370 46756
rect 11426 46700 11494 46756
rect 11550 46700 11618 46756
rect 11674 46700 11742 46756
rect 11798 46700 11866 46756
rect 11922 46700 11990 46756
rect 12046 46700 12114 46756
rect 12170 46700 12180 46756
rect 10244 46632 12180 46700
rect 10244 46576 10254 46632
rect 10310 46576 10378 46632
rect 10434 46576 10502 46632
rect 10558 46576 10626 46632
rect 10682 46576 10750 46632
rect 10806 46576 10874 46632
rect 10930 46576 10998 46632
rect 11054 46576 11122 46632
rect 11178 46576 11246 46632
rect 11302 46576 11370 46632
rect 11426 46576 11494 46632
rect 11550 46576 11618 46632
rect 11674 46576 11742 46632
rect 11798 46576 11866 46632
rect 11922 46576 11990 46632
rect 12046 46576 12114 46632
rect 12170 46576 12180 46632
rect 10244 46508 12180 46576
rect 10244 46452 10254 46508
rect 10310 46452 10378 46508
rect 10434 46452 10502 46508
rect 10558 46452 10626 46508
rect 10682 46452 10750 46508
rect 10806 46452 10874 46508
rect 10930 46452 10998 46508
rect 11054 46452 11122 46508
rect 11178 46452 11246 46508
rect 11302 46452 11370 46508
rect 11426 46452 11494 46508
rect 11550 46452 11618 46508
rect 11674 46452 11742 46508
rect 11798 46452 11866 46508
rect 11922 46452 11990 46508
rect 12046 46452 12114 46508
rect 12170 46452 12180 46508
rect 10244 46442 12180 46452
rect 12861 47252 14673 47281
rect 12861 47196 12871 47252
rect 12927 47196 12995 47252
rect 13051 47196 13119 47252
rect 13175 47196 13243 47252
rect 13299 47196 13367 47252
rect 13423 47196 13491 47252
rect 13547 47196 13615 47252
rect 13671 47196 13739 47252
rect 13795 47196 13863 47252
rect 13919 47196 13987 47252
rect 14043 47196 14111 47252
rect 14167 47196 14235 47252
rect 14291 47196 14359 47252
rect 14415 47196 14483 47252
rect 14539 47196 14607 47252
rect 14663 47196 14673 47252
rect 12861 47128 14673 47196
rect 12861 47072 12871 47128
rect 12927 47072 12995 47128
rect 13051 47072 13119 47128
rect 13175 47072 13243 47128
rect 13299 47072 13367 47128
rect 13423 47072 13491 47128
rect 13547 47072 13615 47128
rect 13671 47072 13739 47128
rect 13795 47072 13863 47128
rect 13919 47072 13987 47128
rect 14043 47072 14111 47128
rect 14167 47072 14235 47128
rect 14291 47072 14359 47128
rect 14415 47072 14483 47128
rect 14539 47072 14607 47128
rect 14663 47072 14673 47128
rect 12861 47004 14673 47072
rect 12861 46948 12871 47004
rect 12927 46948 12995 47004
rect 13051 46948 13119 47004
rect 13175 46948 13243 47004
rect 13299 46948 13367 47004
rect 13423 46948 13491 47004
rect 13547 46948 13615 47004
rect 13671 46948 13739 47004
rect 13795 46948 13863 47004
rect 13919 46948 13987 47004
rect 14043 46948 14111 47004
rect 14167 46948 14235 47004
rect 14291 46948 14359 47004
rect 14415 46948 14483 47004
rect 14539 46948 14607 47004
rect 14663 46948 14673 47004
rect 12861 46880 14673 46948
rect 12861 46824 12871 46880
rect 12927 46824 12995 46880
rect 13051 46824 13119 46880
rect 13175 46824 13243 46880
rect 13299 46824 13367 46880
rect 13423 46824 13491 46880
rect 13547 46824 13615 46880
rect 13671 46824 13739 46880
rect 13795 46824 13863 46880
rect 13919 46824 13987 46880
rect 14043 46824 14111 46880
rect 14167 46824 14235 46880
rect 14291 46824 14359 46880
rect 14415 46824 14483 46880
rect 14539 46824 14607 46880
rect 14663 46824 14673 46880
rect 12861 46756 14673 46824
rect 12861 46700 12871 46756
rect 12927 46700 12995 46756
rect 13051 46700 13119 46756
rect 13175 46700 13243 46756
rect 13299 46700 13367 46756
rect 13423 46700 13491 46756
rect 13547 46700 13615 46756
rect 13671 46700 13739 46756
rect 13795 46700 13863 46756
rect 13919 46700 13987 46756
rect 14043 46700 14111 46756
rect 14167 46700 14235 46756
rect 14291 46700 14359 46756
rect 14415 46700 14483 46756
rect 14539 46700 14607 46756
rect 14663 46700 14673 46756
rect 12861 46632 14673 46700
rect 12861 46576 12871 46632
rect 12927 46576 12995 46632
rect 13051 46576 13119 46632
rect 13175 46576 13243 46632
rect 13299 46576 13367 46632
rect 13423 46576 13491 46632
rect 13547 46576 13615 46632
rect 13671 46576 13739 46632
rect 13795 46576 13863 46632
rect 13919 46576 13987 46632
rect 14043 46576 14111 46632
rect 14167 46576 14235 46632
rect 14291 46576 14359 46632
rect 14415 46576 14483 46632
rect 14539 46576 14607 46632
rect 14663 46576 14673 46632
rect 12861 46508 14673 46576
rect 12861 46452 12871 46508
rect 12927 46452 12995 46508
rect 13051 46452 13119 46508
rect 13175 46452 13243 46508
rect 13299 46452 13367 46508
rect 13423 46452 13491 46508
rect 13547 46452 13615 46508
rect 13671 46452 13739 46508
rect 13795 46452 13863 46508
rect 13919 46452 13987 46508
rect 14043 46452 14111 46508
rect 14167 46452 14235 46508
rect 14291 46452 14359 46508
rect 14415 46452 14483 46508
rect 14539 46452 14607 46508
rect 14663 46452 14673 46508
rect 12861 46442 14673 46452
rect 2481 46148 2681 46158
rect 2481 46092 2491 46148
rect 2547 46092 2615 46148
rect 2671 46092 2681 46148
rect 2481 46024 2681 46092
rect 2481 45968 2491 46024
rect 2547 45968 2615 46024
rect 2671 45968 2681 46024
rect 2481 45900 2681 45968
rect 2481 45844 2491 45900
rect 2547 45844 2615 45900
rect 2671 45844 2681 45900
rect 2481 45776 2681 45844
rect 2481 45720 2491 45776
rect 2547 45720 2615 45776
rect 2671 45720 2681 45776
rect 2481 45652 2681 45720
rect 2481 45596 2491 45652
rect 2547 45596 2615 45652
rect 2671 45596 2681 45652
rect 2481 45528 2681 45596
rect 2481 45472 2491 45528
rect 2547 45472 2615 45528
rect 2671 45472 2681 45528
rect 2481 45404 2681 45472
rect 2481 45348 2491 45404
rect 2547 45348 2615 45404
rect 2671 45348 2681 45404
rect 2481 45280 2681 45348
rect 2481 45224 2491 45280
rect 2547 45224 2615 45280
rect 2671 45224 2681 45280
rect 2481 45156 2681 45224
rect 2481 45100 2491 45156
rect 2547 45100 2615 45156
rect 2671 45100 2681 45156
rect 2481 45032 2681 45100
rect 2481 44976 2491 45032
rect 2547 44976 2615 45032
rect 2671 44976 2681 45032
rect 2481 44908 2681 44976
rect 2481 44852 2491 44908
rect 2547 44852 2615 44908
rect 2671 44852 2681 44908
rect 2481 44842 2681 44852
rect 4851 46148 5051 46158
rect 4851 46092 4861 46148
rect 4917 46092 4985 46148
rect 5041 46092 5051 46148
rect 4851 46024 5051 46092
rect 4851 45968 4861 46024
rect 4917 45968 4985 46024
rect 5041 45968 5051 46024
rect 4851 45900 5051 45968
rect 4851 45844 4861 45900
rect 4917 45844 4985 45900
rect 5041 45844 5051 45900
rect 4851 45776 5051 45844
rect 4851 45720 4861 45776
rect 4917 45720 4985 45776
rect 5041 45720 5051 45776
rect 4851 45652 5051 45720
rect 4851 45596 4861 45652
rect 4917 45596 4985 45652
rect 5041 45596 5051 45652
rect 4851 45528 5051 45596
rect 4851 45472 4861 45528
rect 4917 45472 4985 45528
rect 5041 45472 5051 45528
rect 4851 45404 5051 45472
rect 4851 45348 4861 45404
rect 4917 45348 4985 45404
rect 5041 45348 5051 45404
rect 4851 45280 5051 45348
rect 4851 45224 4861 45280
rect 4917 45224 4985 45280
rect 5041 45224 5051 45280
rect 4851 45156 5051 45224
rect 4851 45100 4861 45156
rect 4917 45100 4985 45156
rect 5041 45100 5051 45156
rect 4851 45032 5051 45100
rect 4851 44976 4861 45032
rect 4917 44976 4985 45032
rect 5041 44976 5051 45032
rect 4851 44908 5051 44976
rect 4851 44852 4861 44908
rect 4917 44852 4985 44908
rect 5041 44852 5051 44908
rect 4851 44842 5051 44852
rect 7265 46148 7713 46158
rect 7265 46092 7275 46148
rect 7331 46092 7399 46148
rect 7455 46092 7523 46148
rect 7579 46092 7647 46148
rect 7703 46092 7713 46148
rect 7265 46024 7713 46092
rect 7265 45968 7275 46024
rect 7331 45968 7399 46024
rect 7455 45968 7523 46024
rect 7579 45968 7647 46024
rect 7703 45968 7713 46024
rect 7265 45900 7713 45968
rect 7265 45844 7275 45900
rect 7331 45844 7399 45900
rect 7455 45844 7523 45900
rect 7579 45844 7647 45900
rect 7703 45844 7713 45900
rect 7265 45776 7713 45844
rect 7265 45720 7275 45776
rect 7331 45720 7399 45776
rect 7455 45720 7523 45776
rect 7579 45720 7647 45776
rect 7703 45720 7713 45776
rect 7265 45652 7713 45720
rect 7265 45596 7275 45652
rect 7331 45596 7399 45652
rect 7455 45596 7523 45652
rect 7579 45596 7647 45652
rect 7703 45596 7713 45652
rect 7265 45528 7713 45596
rect 7265 45472 7275 45528
rect 7331 45472 7399 45528
rect 7455 45472 7523 45528
rect 7579 45472 7647 45528
rect 7703 45472 7713 45528
rect 7265 45404 7713 45472
rect 7265 45348 7275 45404
rect 7331 45348 7399 45404
rect 7455 45348 7523 45404
rect 7579 45348 7647 45404
rect 7703 45348 7713 45404
rect 7265 45280 7713 45348
rect 7265 45224 7275 45280
rect 7331 45224 7399 45280
rect 7455 45224 7523 45280
rect 7579 45224 7647 45280
rect 7703 45224 7713 45280
rect 7265 45156 7713 45224
rect 7265 45100 7275 45156
rect 7331 45100 7399 45156
rect 7455 45100 7523 45156
rect 7579 45100 7647 45156
rect 7703 45100 7713 45156
rect 7265 45032 7713 45100
rect 7265 44976 7275 45032
rect 7331 44976 7399 45032
rect 7455 44976 7523 45032
rect 7579 44976 7647 45032
rect 7703 44976 7713 45032
rect 7265 44908 7713 44976
rect 7265 44852 7275 44908
rect 7331 44852 7399 44908
rect 7455 44852 7523 44908
rect 7579 44852 7647 44908
rect 7703 44852 7713 44908
rect 7265 44842 7713 44852
rect 9927 46148 10127 46158
rect 9927 46092 9937 46148
rect 9993 46092 10061 46148
rect 10117 46092 10127 46148
rect 9927 46024 10127 46092
rect 9927 45968 9937 46024
rect 9993 45968 10061 46024
rect 10117 45968 10127 46024
rect 9927 45900 10127 45968
rect 9927 45844 9937 45900
rect 9993 45844 10061 45900
rect 10117 45844 10127 45900
rect 9927 45776 10127 45844
rect 9927 45720 9937 45776
rect 9993 45720 10061 45776
rect 10117 45720 10127 45776
rect 9927 45652 10127 45720
rect 9927 45596 9937 45652
rect 9993 45596 10061 45652
rect 10117 45596 10127 45652
rect 9927 45528 10127 45596
rect 9927 45472 9937 45528
rect 9993 45472 10061 45528
rect 10117 45472 10127 45528
rect 9927 45404 10127 45472
rect 9927 45348 9937 45404
rect 9993 45348 10061 45404
rect 10117 45348 10127 45404
rect 9927 45280 10127 45348
rect 9927 45224 9937 45280
rect 9993 45224 10061 45280
rect 10117 45224 10127 45280
rect 9927 45156 10127 45224
rect 9927 45100 9937 45156
rect 9993 45100 10061 45156
rect 10117 45100 10127 45156
rect 9927 45032 10127 45100
rect 9927 44976 9937 45032
rect 9993 44976 10061 45032
rect 10117 44976 10127 45032
rect 9927 44908 10127 44976
rect 9927 44852 9937 44908
rect 9993 44852 10061 44908
rect 10117 44852 10127 44908
rect 9927 44842 10127 44852
rect 12297 46148 12497 46158
rect 12297 46092 12307 46148
rect 12363 46092 12431 46148
rect 12487 46092 12497 46148
rect 12297 46024 12497 46092
rect 12297 45968 12307 46024
rect 12363 45968 12431 46024
rect 12487 45968 12497 46024
rect 12297 45900 12497 45968
rect 12297 45844 12307 45900
rect 12363 45844 12431 45900
rect 12487 45844 12497 45900
rect 12297 45776 12497 45844
rect 12297 45720 12307 45776
rect 12363 45720 12431 45776
rect 12487 45720 12497 45776
rect 12297 45652 12497 45720
rect 12297 45596 12307 45652
rect 12363 45596 12431 45652
rect 12487 45596 12497 45652
rect 12297 45528 12497 45596
rect 12297 45472 12307 45528
rect 12363 45472 12431 45528
rect 12487 45472 12497 45528
rect 12297 45404 12497 45472
rect 12297 45348 12307 45404
rect 12363 45348 12431 45404
rect 12487 45348 12497 45404
rect 12297 45280 12497 45348
rect 12297 45224 12307 45280
rect 12363 45224 12431 45280
rect 12487 45224 12497 45280
rect 12297 45156 12497 45224
rect 12297 45100 12307 45156
rect 12363 45100 12431 45156
rect 12487 45100 12497 45156
rect 12297 45032 12497 45100
rect 12297 44976 12307 45032
rect 12363 44976 12431 45032
rect 12487 44976 12497 45032
rect 12297 44908 12497 44976
rect 12297 44852 12307 44908
rect 12363 44852 12431 44908
rect 12487 44852 12497 44908
rect 12297 44842 12497 44852
rect 2798 44548 4734 44558
rect 2798 44492 2808 44548
rect 2864 44492 2932 44548
rect 2988 44492 3056 44548
rect 3112 44492 3180 44548
rect 3236 44492 3304 44548
rect 3360 44492 3428 44548
rect 3484 44492 3552 44548
rect 3608 44492 3676 44548
rect 3732 44492 3800 44548
rect 3856 44492 3924 44548
rect 3980 44492 4048 44548
rect 4104 44492 4172 44548
rect 4228 44492 4296 44548
rect 4352 44492 4420 44548
rect 4476 44492 4544 44548
rect 4600 44492 4668 44548
rect 4724 44492 4734 44548
rect 2798 44424 4734 44492
rect 2798 44368 2808 44424
rect 2864 44368 2932 44424
rect 2988 44368 3056 44424
rect 3112 44368 3180 44424
rect 3236 44368 3304 44424
rect 3360 44368 3428 44424
rect 3484 44368 3552 44424
rect 3608 44368 3676 44424
rect 3732 44368 3800 44424
rect 3856 44368 3924 44424
rect 3980 44368 4048 44424
rect 4104 44368 4172 44424
rect 4228 44368 4296 44424
rect 4352 44368 4420 44424
rect 4476 44368 4544 44424
rect 4600 44368 4668 44424
rect 4724 44368 4734 44424
rect 2798 44300 4734 44368
rect 2798 44244 2808 44300
rect 2864 44244 2932 44300
rect 2988 44244 3056 44300
rect 3112 44244 3180 44300
rect 3236 44244 3304 44300
rect 3360 44244 3428 44300
rect 3484 44244 3552 44300
rect 3608 44244 3676 44300
rect 3732 44244 3800 44300
rect 3856 44244 3924 44300
rect 3980 44244 4048 44300
rect 4104 44244 4172 44300
rect 4228 44244 4296 44300
rect 4352 44244 4420 44300
rect 4476 44244 4544 44300
rect 4600 44244 4668 44300
rect 4724 44244 4734 44300
rect 2798 44176 4734 44244
rect 2798 44120 2808 44176
rect 2864 44120 2932 44176
rect 2988 44120 3056 44176
rect 3112 44120 3180 44176
rect 3236 44120 3304 44176
rect 3360 44120 3428 44176
rect 3484 44120 3552 44176
rect 3608 44120 3676 44176
rect 3732 44120 3800 44176
rect 3856 44120 3924 44176
rect 3980 44120 4048 44176
rect 4104 44120 4172 44176
rect 4228 44120 4296 44176
rect 4352 44120 4420 44176
rect 4476 44120 4544 44176
rect 4600 44120 4668 44176
rect 4724 44120 4734 44176
rect 2798 44052 4734 44120
rect 2798 43996 2808 44052
rect 2864 43996 2932 44052
rect 2988 43996 3056 44052
rect 3112 43996 3180 44052
rect 3236 43996 3304 44052
rect 3360 43996 3428 44052
rect 3484 43996 3552 44052
rect 3608 43996 3676 44052
rect 3732 43996 3800 44052
rect 3856 43996 3924 44052
rect 3980 43996 4048 44052
rect 4104 43996 4172 44052
rect 4228 43996 4296 44052
rect 4352 43996 4420 44052
rect 4476 43996 4544 44052
rect 4600 43996 4668 44052
rect 4724 43996 4734 44052
rect 2798 43928 4734 43996
rect 2798 43872 2808 43928
rect 2864 43872 2932 43928
rect 2988 43872 3056 43928
rect 3112 43872 3180 43928
rect 3236 43872 3304 43928
rect 3360 43872 3428 43928
rect 3484 43872 3552 43928
rect 3608 43872 3676 43928
rect 3732 43872 3800 43928
rect 3856 43872 3924 43928
rect 3980 43872 4048 43928
rect 4104 43872 4172 43928
rect 4228 43872 4296 43928
rect 4352 43872 4420 43928
rect 4476 43872 4544 43928
rect 4600 43872 4668 43928
rect 4724 43872 4734 43928
rect 2798 43804 4734 43872
rect 2798 43748 2808 43804
rect 2864 43748 2932 43804
rect 2988 43748 3056 43804
rect 3112 43748 3180 43804
rect 3236 43748 3304 43804
rect 3360 43748 3428 43804
rect 3484 43748 3552 43804
rect 3608 43748 3676 43804
rect 3732 43748 3800 43804
rect 3856 43748 3924 43804
rect 3980 43748 4048 43804
rect 4104 43748 4172 43804
rect 4228 43748 4296 43804
rect 4352 43748 4420 43804
rect 4476 43748 4544 43804
rect 4600 43748 4668 43804
rect 4724 43748 4734 43804
rect 2798 43680 4734 43748
rect 2798 43624 2808 43680
rect 2864 43624 2932 43680
rect 2988 43624 3056 43680
rect 3112 43624 3180 43680
rect 3236 43624 3304 43680
rect 3360 43624 3428 43680
rect 3484 43624 3552 43680
rect 3608 43624 3676 43680
rect 3732 43624 3800 43680
rect 3856 43624 3924 43680
rect 3980 43624 4048 43680
rect 4104 43624 4172 43680
rect 4228 43624 4296 43680
rect 4352 43624 4420 43680
rect 4476 43624 4544 43680
rect 4600 43624 4668 43680
rect 4724 43624 4734 43680
rect 2798 43556 4734 43624
rect 2798 43500 2808 43556
rect 2864 43500 2932 43556
rect 2988 43500 3056 43556
rect 3112 43500 3180 43556
rect 3236 43500 3304 43556
rect 3360 43500 3428 43556
rect 3484 43500 3552 43556
rect 3608 43500 3676 43556
rect 3732 43500 3800 43556
rect 3856 43500 3924 43556
rect 3980 43500 4048 43556
rect 4104 43500 4172 43556
rect 4228 43500 4296 43556
rect 4352 43500 4420 43556
rect 4476 43500 4544 43556
rect 4600 43500 4668 43556
rect 4724 43500 4734 43556
rect 2798 43432 4734 43500
rect 2798 43376 2808 43432
rect 2864 43376 2932 43432
rect 2988 43376 3056 43432
rect 3112 43376 3180 43432
rect 3236 43376 3304 43432
rect 3360 43376 3428 43432
rect 3484 43376 3552 43432
rect 3608 43376 3676 43432
rect 3732 43376 3800 43432
rect 3856 43376 3924 43432
rect 3980 43376 4048 43432
rect 4104 43376 4172 43432
rect 4228 43376 4296 43432
rect 4352 43376 4420 43432
rect 4476 43376 4544 43432
rect 4600 43376 4668 43432
rect 4724 43376 4734 43432
rect 2798 43308 4734 43376
rect 2798 43252 2808 43308
rect 2864 43252 2932 43308
rect 2988 43252 3056 43308
rect 3112 43252 3180 43308
rect 3236 43252 3304 43308
rect 3360 43252 3428 43308
rect 3484 43252 3552 43308
rect 3608 43252 3676 43308
rect 3732 43252 3800 43308
rect 3856 43252 3924 43308
rect 3980 43252 4048 43308
rect 4104 43252 4172 43308
rect 4228 43252 4296 43308
rect 4352 43252 4420 43308
rect 4476 43252 4544 43308
rect 4600 43252 4668 43308
rect 4724 43252 4734 43308
rect 2798 43242 4734 43252
rect 5168 44548 7104 44558
rect 5168 44492 5178 44548
rect 5234 44492 5302 44548
rect 5358 44492 5426 44548
rect 5482 44492 5550 44548
rect 5606 44492 5674 44548
rect 5730 44492 5798 44548
rect 5854 44492 5922 44548
rect 5978 44492 6046 44548
rect 6102 44492 6170 44548
rect 6226 44492 6294 44548
rect 6350 44492 6418 44548
rect 6474 44492 6542 44548
rect 6598 44492 6666 44548
rect 6722 44492 6790 44548
rect 6846 44492 6914 44548
rect 6970 44492 7038 44548
rect 7094 44492 7104 44548
rect 5168 44424 7104 44492
rect 5168 44368 5178 44424
rect 5234 44368 5302 44424
rect 5358 44368 5426 44424
rect 5482 44368 5550 44424
rect 5606 44368 5674 44424
rect 5730 44368 5798 44424
rect 5854 44368 5922 44424
rect 5978 44368 6046 44424
rect 6102 44368 6170 44424
rect 6226 44368 6294 44424
rect 6350 44368 6418 44424
rect 6474 44368 6542 44424
rect 6598 44368 6666 44424
rect 6722 44368 6790 44424
rect 6846 44368 6914 44424
rect 6970 44368 7038 44424
rect 7094 44368 7104 44424
rect 5168 44300 7104 44368
rect 5168 44244 5178 44300
rect 5234 44244 5302 44300
rect 5358 44244 5426 44300
rect 5482 44244 5550 44300
rect 5606 44244 5674 44300
rect 5730 44244 5798 44300
rect 5854 44244 5922 44300
rect 5978 44244 6046 44300
rect 6102 44244 6170 44300
rect 6226 44244 6294 44300
rect 6350 44244 6418 44300
rect 6474 44244 6542 44300
rect 6598 44244 6666 44300
rect 6722 44244 6790 44300
rect 6846 44244 6914 44300
rect 6970 44244 7038 44300
rect 7094 44244 7104 44300
rect 5168 44176 7104 44244
rect 5168 44120 5178 44176
rect 5234 44120 5302 44176
rect 5358 44120 5426 44176
rect 5482 44120 5550 44176
rect 5606 44120 5674 44176
rect 5730 44120 5798 44176
rect 5854 44120 5922 44176
rect 5978 44120 6046 44176
rect 6102 44120 6170 44176
rect 6226 44120 6294 44176
rect 6350 44120 6418 44176
rect 6474 44120 6542 44176
rect 6598 44120 6666 44176
rect 6722 44120 6790 44176
rect 6846 44120 6914 44176
rect 6970 44120 7038 44176
rect 7094 44120 7104 44176
rect 5168 44052 7104 44120
rect 5168 43996 5178 44052
rect 5234 43996 5302 44052
rect 5358 43996 5426 44052
rect 5482 43996 5550 44052
rect 5606 43996 5674 44052
rect 5730 43996 5798 44052
rect 5854 43996 5922 44052
rect 5978 43996 6046 44052
rect 6102 43996 6170 44052
rect 6226 43996 6294 44052
rect 6350 43996 6418 44052
rect 6474 43996 6542 44052
rect 6598 43996 6666 44052
rect 6722 43996 6790 44052
rect 6846 43996 6914 44052
rect 6970 43996 7038 44052
rect 7094 43996 7104 44052
rect 5168 43928 7104 43996
rect 5168 43872 5178 43928
rect 5234 43872 5302 43928
rect 5358 43872 5426 43928
rect 5482 43872 5550 43928
rect 5606 43872 5674 43928
rect 5730 43872 5798 43928
rect 5854 43872 5922 43928
rect 5978 43872 6046 43928
rect 6102 43872 6170 43928
rect 6226 43872 6294 43928
rect 6350 43872 6418 43928
rect 6474 43872 6542 43928
rect 6598 43872 6666 43928
rect 6722 43872 6790 43928
rect 6846 43872 6914 43928
rect 6970 43872 7038 43928
rect 7094 43872 7104 43928
rect 5168 43804 7104 43872
rect 5168 43748 5178 43804
rect 5234 43748 5302 43804
rect 5358 43748 5426 43804
rect 5482 43748 5550 43804
rect 5606 43748 5674 43804
rect 5730 43748 5798 43804
rect 5854 43748 5922 43804
rect 5978 43748 6046 43804
rect 6102 43748 6170 43804
rect 6226 43748 6294 43804
rect 6350 43748 6418 43804
rect 6474 43748 6542 43804
rect 6598 43748 6666 43804
rect 6722 43748 6790 43804
rect 6846 43748 6914 43804
rect 6970 43748 7038 43804
rect 7094 43748 7104 43804
rect 5168 43680 7104 43748
rect 5168 43624 5178 43680
rect 5234 43624 5302 43680
rect 5358 43624 5426 43680
rect 5482 43624 5550 43680
rect 5606 43624 5674 43680
rect 5730 43624 5798 43680
rect 5854 43624 5922 43680
rect 5978 43624 6046 43680
rect 6102 43624 6170 43680
rect 6226 43624 6294 43680
rect 6350 43624 6418 43680
rect 6474 43624 6542 43680
rect 6598 43624 6666 43680
rect 6722 43624 6790 43680
rect 6846 43624 6914 43680
rect 6970 43624 7038 43680
rect 7094 43624 7104 43680
rect 5168 43556 7104 43624
rect 5168 43500 5178 43556
rect 5234 43500 5302 43556
rect 5358 43500 5426 43556
rect 5482 43500 5550 43556
rect 5606 43500 5674 43556
rect 5730 43500 5798 43556
rect 5854 43500 5922 43556
rect 5978 43500 6046 43556
rect 6102 43500 6170 43556
rect 6226 43500 6294 43556
rect 6350 43500 6418 43556
rect 6474 43500 6542 43556
rect 6598 43500 6666 43556
rect 6722 43500 6790 43556
rect 6846 43500 6914 43556
rect 6970 43500 7038 43556
rect 7094 43500 7104 43556
rect 5168 43432 7104 43500
rect 5168 43376 5178 43432
rect 5234 43376 5302 43432
rect 5358 43376 5426 43432
rect 5482 43376 5550 43432
rect 5606 43376 5674 43432
rect 5730 43376 5798 43432
rect 5854 43376 5922 43432
rect 5978 43376 6046 43432
rect 6102 43376 6170 43432
rect 6226 43376 6294 43432
rect 6350 43376 6418 43432
rect 6474 43376 6542 43432
rect 6598 43376 6666 43432
rect 6722 43376 6790 43432
rect 6846 43376 6914 43432
rect 6970 43376 7038 43432
rect 7094 43376 7104 43432
rect 5168 43308 7104 43376
rect 5168 43252 5178 43308
rect 5234 43252 5302 43308
rect 5358 43252 5426 43308
rect 5482 43252 5550 43308
rect 5606 43252 5674 43308
rect 5730 43252 5798 43308
rect 5854 43252 5922 43308
rect 5978 43252 6046 43308
rect 6102 43252 6170 43308
rect 6226 43252 6294 43308
rect 6350 43252 6418 43308
rect 6474 43252 6542 43308
rect 6598 43252 6666 43308
rect 6722 43252 6790 43308
rect 6846 43252 6914 43308
rect 6970 43252 7038 43308
rect 7094 43252 7104 43308
rect 5168 43242 7104 43252
rect 7874 44548 9810 44558
rect 7874 44492 7884 44548
rect 7940 44492 8008 44548
rect 8064 44492 8132 44548
rect 8188 44492 8256 44548
rect 8312 44492 8380 44548
rect 8436 44492 8504 44548
rect 8560 44492 8628 44548
rect 8684 44492 8752 44548
rect 8808 44492 8876 44548
rect 8932 44492 9000 44548
rect 9056 44492 9124 44548
rect 9180 44492 9248 44548
rect 9304 44492 9372 44548
rect 9428 44492 9496 44548
rect 9552 44492 9620 44548
rect 9676 44492 9744 44548
rect 9800 44492 9810 44548
rect 7874 44424 9810 44492
rect 7874 44368 7884 44424
rect 7940 44368 8008 44424
rect 8064 44368 8132 44424
rect 8188 44368 8256 44424
rect 8312 44368 8380 44424
rect 8436 44368 8504 44424
rect 8560 44368 8628 44424
rect 8684 44368 8752 44424
rect 8808 44368 8876 44424
rect 8932 44368 9000 44424
rect 9056 44368 9124 44424
rect 9180 44368 9248 44424
rect 9304 44368 9372 44424
rect 9428 44368 9496 44424
rect 9552 44368 9620 44424
rect 9676 44368 9744 44424
rect 9800 44368 9810 44424
rect 7874 44300 9810 44368
rect 7874 44244 7884 44300
rect 7940 44244 8008 44300
rect 8064 44244 8132 44300
rect 8188 44244 8256 44300
rect 8312 44244 8380 44300
rect 8436 44244 8504 44300
rect 8560 44244 8628 44300
rect 8684 44244 8752 44300
rect 8808 44244 8876 44300
rect 8932 44244 9000 44300
rect 9056 44244 9124 44300
rect 9180 44244 9248 44300
rect 9304 44244 9372 44300
rect 9428 44244 9496 44300
rect 9552 44244 9620 44300
rect 9676 44244 9744 44300
rect 9800 44244 9810 44300
rect 7874 44176 9810 44244
rect 7874 44120 7884 44176
rect 7940 44120 8008 44176
rect 8064 44120 8132 44176
rect 8188 44120 8256 44176
rect 8312 44120 8380 44176
rect 8436 44120 8504 44176
rect 8560 44120 8628 44176
rect 8684 44120 8752 44176
rect 8808 44120 8876 44176
rect 8932 44120 9000 44176
rect 9056 44120 9124 44176
rect 9180 44120 9248 44176
rect 9304 44120 9372 44176
rect 9428 44120 9496 44176
rect 9552 44120 9620 44176
rect 9676 44120 9744 44176
rect 9800 44120 9810 44176
rect 7874 44052 9810 44120
rect 7874 43996 7884 44052
rect 7940 43996 8008 44052
rect 8064 43996 8132 44052
rect 8188 43996 8256 44052
rect 8312 43996 8380 44052
rect 8436 43996 8504 44052
rect 8560 43996 8628 44052
rect 8684 43996 8752 44052
rect 8808 43996 8876 44052
rect 8932 43996 9000 44052
rect 9056 43996 9124 44052
rect 9180 43996 9248 44052
rect 9304 43996 9372 44052
rect 9428 43996 9496 44052
rect 9552 43996 9620 44052
rect 9676 43996 9744 44052
rect 9800 43996 9810 44052
rect 7874 43928 9810 43996
rect 7874 43872 7884 43928
rect 7940 43872 8008 43928
rect 8064 43872 8132 43928
rect 8188 43872 8256 43928
rect 8312 43872 8380 43928
rect 8436 43872 8504 43928
rect 8560 43872 8628 43928
rect 8684 43872 8752 43928
rect 8808 43872 8876 43928
rect 8932 43872 9000 43928
rect 9056 43872 9124 43928
rect 9180 43872 9248 43928
rect 9304 43872 9372 43928
rect 9428 43872 9496 43928
rect 9552 43872 9620 43928
rect 9676 43872 9744 43928
rect 9800 43872 9810 43928
rect 7874 43804 9810 43872
rect 7874 43748 7884 43804
rect 7940 43748 8008 43804
rect 8064 43748 8132 43804
rect 8188 43748 8256 43804
rect 8312 43748 8380 43804
rect 8436 43748 8504 43804
rect 8560 43748 8628 43804
rect 8684 43748 8752 43804
rect 8808 43748 8876 43804
rect 8932 43748 9000 43804
rect 9056 43748 9124 43804
rect 9180 43748 9248 43804
rect 9304 43748 9372 43804
rect 9428 43748 9496 43804
rect 9552 43748 9620 43804
rect 9676 43748 9744 43804
rect 9800 43748 9810 43804
rect 7874 43680 9810 43748
rect 7874 43624 7884 43680
rect 7940 43624 8008 43680
rect 8064 43624 8132 43680
rect 8188 43624 8256 43680
rect 8312 43624 8380 43680
rect 8436 43624 8504 43680
rect 8560 43624 8628 43680
rect 8684 43624 8752 43680
rect 8808 43624 8876 43680
rect 8932 43624 9000 43680
rect 9056 43624 9124 43680
rect 9180 43624 9248 43680
rect 9304 43624 9372 43680
rect 9428 43624 9496 43680
rect 9552 43624 9620 43680
rect 9676 43624 9744 43680
rect 9800 43624 9810 43680
rect 7874 43556 9810 43624
rect 7874 43500 7884 43556
rect 7940 43500 8008 43556
rect 8064 43500 8132 43556
rect 8188 43500 8256 43556
rect 8312 43500 8380 43556
rect 8436 43500 8504 43556
rect 8560 43500 8628 43556
rect 8684 43500 8752 43556
rect 8808 43500 8876 43556
rect 8932 43500 9000 43556
rect 9056 43500 9124 43556
rect 9180 43500 9248 43556
rect 9304 43500 9372 43556
rect 9428 43500 9496 43556
rect 9552 43500 9620 43556
rect 9676 43500 9744 43556
rect 9800 43500 9810 43556
rect 7874 43432 9810 43500
rect 7874 43376 7884 43432
rect 7940 43376 8008 43432
rect 8064 43376 8132 43432
rect 8188 43376 8256 43432
rect 8312 43376 8380 43432
rect 8436 43376 8504 43432
rect 8560 43376 8628 43432
rect 8684 43376 8752 43432
rect 8808 43376 8876 43432
rect 8932 43376 9000 43432
rect 9056 43376 9124 43432
rect 9180 43376 9248 43432
rect 9304 43376 9372 43432
rect 9428 43376 9496 43432
rect 9552 43376 9620 43432
rect 9676 43376 9744 43432
rect 9800 43376 9810 43432
rect 7874 43308 9810 43376
rect 7874 43252 7884 43308
rect 7940 43252 8008 43308
rect 8064 43252 8132 43308
rect 8188 43252 8256 43308
rect 8312 43252 8380 43308
rect 8436 43252 8504 43308
rect 8560 43252 8628 43308
rect 8684 43252 8752 43308
rect 8808 43252 8876 43308
rect 8932 43252 9000 43308
rect 9056 43252 9124 43308
rect 9180 43252 9248 43308
rect 9304 43252 9372 43308
rect 9428 43252 9496 43308
rect 9552 43252 9620 43308
rect 9676 43252 9744 43308
rect 9800 43252 9810 43308
rect 7874 43242 9810 43252
rect 10244 44548 12180 44558
rect 10244 44492 10254 44548
rect 10310 44492 10378 44548
rect 10434 44492 10502 44548
rect 10558 44492 10626 44548
rect 10682 44492 10750 44548
rect 10806 44492 10874 44548
rect 10930 44492 10998 44548
rect 11054 44492 11122 44548
rect 11178 44492 11246 44548
rect 11302 44492 11370 44548
rect 11426 44492 11494 44548
rect 11550 44492 11618 44548
rect 11674 44492 11742 44548
rect 11798 44492 11866 44548
rect 11922 44492 11990 44548
rect 12046 44492 12114 44548
rect 12170 44492 12180 44548
rect 10244 44424 12180 44492
rect 10244 44368 10254 44424
rect 10310 44368 10378 44424
rect 10434 44368 10502 44424
rect 10558 44368 10626 44424
rect 10682 44368 10750 44424
rect 10806 44368 10874 44424
rect 10930 44368 10998 44424
rect 11054 44368 11122 44424
rect 11178 44368 11246 44424
rect 11302 44368 11370 44424
rect 11426 44368 11494 44424
rect 11550 44368 11618 44424
rect 11674 44368 11742 44424
rect 11798 44368 11866 44424
rect 11922 44368 11990 44424
rect 12046 44368 12114 44424
rect 12170 44368 12180 44424
rect 10244 44300 12180 44368
rect 10244 44244 10254 44300
rect 10310 44244 10378 44300
rect 10434 44244 10502 44300
rect 10558 44244 10626 44300
rect 10682 44244 10750 44300
rect 10806 44244 10874 44300
rect 10930 44244 10998 44300
rect 11054 44244 11122 44300
rect 11178 44244 11246 44300
rect 11302 44244 11370 44300
rect 11426 44244 11494 44300
rect 11550 44244 11618 44300
rect 11674 44244 11742 44300
rect 11798 44244 11866 44300
rect 11922 44244 11990 44300
rect 12046 44244 12114 44300
rect 12170 44244 12180 44300
rect 10244 44176 12180 44244
rect 10244 44120 10254 44176
rect 10310 44120 10378 44176
rect 10434 44120 10502 44176
rect 10558 44120 10626 44176
rect 10682 44120 10750 44176
rect 10806 44120 10874 44176
rect 10930 44120 10998 44176
rect 11054 44120 11122 44176
rect 11178 44120 11246 44176
rect 11302 44120 11370 44176
rect 11426 44120 11494 44176
rect 11550 44120 11618 44176
rect 11674 44120 11742 44176
rect 11798 44120 11866 44176
rect 11922 44120 11990 44176
rect 12046 44120 12114 44176
rect 12170 44120 12180 44176
rect 10244 44052 12180 44120
rect 10244 43996 10254 44052
rect 10310 43996 10378 44052
rect 10434 43996 10502 44052
rect 10558 43996 10626 44052
rect 10682 43996 10750 44052
rect 10806 43996 10874 44052
rect 10930 43996 10998 44052
rect 11054 43996 11122 44052
rect 11178 43996 11246 44052
rect 11302 43996 11370 44052
rect 11426 43996 11494 44052
rect 11550 43996 11618 44052
rect 11674 43996 11742 44052
rect 11798 43996 11866 44052
rect 11922 43996 11990 44052
rect 12046 43996 12114 44052
rect 12170 43996 12180 44052
rect 10244 43928 12180 43996
rect 10244 43872 10254 43928
rect 10310 43872 10378 43928
rect 10434 43872 10502 43928
rect 10558 43872 10626 43928
rect 10682 43872 10750 43928
rect 10806 43872 10874 43928
rect 10930 43872 10998 43928
rect 11054 43872 11122 43928
rect 11178 43872 11246 43928
rect 11302 43872 11370 43928
rect 11426 43872 11494 43928
rect 11550 43872 11618 43928
rect 11674 43872 11742 43928
rect 11798 43872 11866 43928
rect 11922 43872 11990 43928
rect 12046 43872 12114 43928
rect 12170 43872 12180 43928
rect 10244 43804 12180 43872
rect 10244 43748 10254 43804
rect 10310 43748 10378 43804
rect 10434 43748 10502 43804
rect 10558 43748 10626 43804
rect 10682 43748 10750 43804
rect 10806 43748 10874 43804
rect 10930 43748 10998 43804
rect 11054 43748 11122 43804
rect 11178 43748 11246 43804
rect 11302 43748 11370 43804
rect 11426 43748 11494 43804
rect 11550 43748 11618 43804
rect 11674 43748 11742 43804
rect 11798 43748 11866 43804
rect 11922 43748 11990 43804
rect 12046 43748 12114 43804
rect 12170 43748 12180 43804
rect 10244 43680 12180 43748
rect 10244 43624 10254 43680
rect 10310 43624 10378 43680
rect 10434 43624 10502 43680
rect 10558 43624 10626 43680
rect 10682 43624 10750 43680
rect 10806 43624 10874 43680
rect 10930 43624 10998 43680
rect 11054 43624 11122 43680
rect 11178 43624 11246 43680
rect 11302 43624 11370 43680
rect 11426 43624 11494 43680
rect 11550 43624 11618 43680
rect 11674 43624 11742 43680
rect 11798 43624 11866 43680
rect 11922 43624 11990 43680
rect 12046 43624 12114 43680
rect 12170 43624 12180 43680
rect 10244 43556 12180 43624
rect 10244 43500 10254 43556
rect 10310 43500 10378 43556
rect 10434 43500 10502 43556
rect 10558 43500 10626 43556
rect 10682 43500 10750 43556
rect 10806 43500 10874 43556
rect 10930 43500 10998 43556
rect 11054 43500 11122 43556
rect 11178 43500 11246 43556
rect 11302 43500 11370 43556
rect 11426 43500 11494 43556
rect 11550 43500 11618 43556
rect 11674 43500 11742 43556
rect 11798 43500 11866 43556
rect 11922 43500 11990 43556
rect 12046 43500 12114 43556
rect 12170 43500 12180 43556
rect 10244 43432 12180 43500
rect 10244 43376 10254 43432
rect 10310 43376 10378 43432
rect 10434 43376 10502 43432
rect 10558 43376 10626 43432
rect 10682 43376 10750 43432
rect 10806 43376 10874 43432
rect 10930 43376 10998 43432
rect 11054 43376 11122 43432
rect 11178 43376 11246 43432
rect 11302 43376 11370 43432
rect 11426 43376 11494 43432
rect 11550 43376 11618 43432
rect 11674 43376 11742 43432
rect 11798 43376 11866 43432
rect 11922 43376 11990 43432
rect 12046 43376 12114 43432
rect 12170 43376 12180 43432
rect 10244 43308 12180 43376
rect 10244 43252 10254 43308
rect 10310 43252 10378 43308
rect 10434 43252 10502 43308
rect 10558 43252 10626 43308
rect 10682 43252 10750 43308
rect 10806 43252 10874 43308
rect 10930 43252 10998 43308
rect 11054 43252 11122 43308
rect 11178 43252 11246 43308
rect 11302 43252 11370 43308
rect 11426 43252 11494 43308
rect 11550 43252 11618 43308
rect 11674 43252 11742 43308
rect 11798 43252 11866 43308
rect 11922 43252 11990 43308
rect 12046 43252 12114 43308
rect 12170 43252 12180 43308
rect 10244 43242 12180 43252
rect 12861 44548 14673 44558
rect 12861 44492 12871 44548
rect 12927 44492 12995 44548
rect 13051 44492 13119 44548
rect 13175 44492 13243 44548
rect 13299 44492 13367 44548
rect 13423 44492 13491 44548
rect 13547 44492 13615 44548
rect 13671 44492 13739 44548
rect 13795 44492 13863 44548
rect 13919 44492 13987 44548
rect 14043 44492 14111 44548
rect 14167 44492 14235 44548
rect 14291 44492 14359 44548
rect 14415 44492 14483 44548
rect 14539 44492 14607 44548
rect 14663 44492 14673 44548
rect 12861 44424 14673 44492
rect 12861 44368 12871 44424
rect 12927 44368 12995 44424
rect 13051 44368 13119 44424
rect 13175 44368 13243 44424
rect 13299 44368 13367 44424
rect 13423 44368 13491 44424
rect 13547 44368 13615 44424
rect 13671 44368 13739 44424
rect 13795 44368 13863 44424
rect 13919 44368 13987 44424
rect 14043 44368 14111 44424
rect 14167 44368 14235 44424
rect 14291 44368 14359 44424
rect 14415 44368 14483 44424
rect 14539 44368 14607 44424
rect 14663 44368 14673 44424
rect 12861 44300 14673 44368
rect 12861 44244 12871 44300
rect 12927 44244 12995 44300
rect 13051 44244 13119 44300
rect 13175 44244 13243 44300
rect 13299 44244 13367 44300
rect 13423 44244 13491 44300
rect 13547 44244 13615 44300
rect 13671 44244 13739 44300
rect 13795 44244 13863 44300
rect 13919 44244 13987 44300
rect 14043 44244 14111 44300
rect 14167 44244 14235 44300
rect 14291 44244 14359 44300
rect 14415 44244 14483 44300
rect 14539 44244 14607 44300
rect 14663 44244 14673 44300
rect 12861 44176 14673 44244
rect 12861 44120 12871 44176
rect 12927 44120 12995 44176
rect 13051 44120 13119 44176
rect 13175 44120 13243 44176
rect 13299 44120 13367 44176
rect 13423 44120 13491 44176
rect 13547 44120 13615 44176
rect 13671 44120 13739 44176
rect 13795 44120 13863 44176
rect 13919 44120 13987 44176
rect 14043 44120 14111 44176
rect 14167 44120 14235 44176
rect 14291 44120 14359 44176
rect 14415 44120 14483 44176
rect 14539 44120 14607 44176
rect 14663 44120 14673 44176
rect 12861 44052 14673 44120
rect 12861 43996 12871 44052
rect 12927 43996 12995 44052
rect 13051 43996 13119 44052
rect 13175 43996 13243 44052
rect 13299 43996 13367 44052
rect 13423 43996 13491 44052
rect 13547 43996 13615 44052
rect 13671 43996 13739 44052
rect 13795 43996 13863 44052
rect 13919 43996 13987 44052
rect 14043 43996 14111 44052
rect 14167 43996 14235 44052
rect 14291 43996 14359 44052
rect 14415 43996 14483 44052
rect 14539 43996 14607 44052
rect 14663 43996 14673 44052
rect 12861 43928 14673 43996
rect 12861 43872 12871 43928
rect 12927 43872 12995 43928
rect 13051 43872 13119 43928
rect 13175 43872 13243 43928
rect 13299 43872 13367 43928
rect 13423 43872 13491 43928
rect 13547 43872 13615 43928
rect 13671 43872 13739 43928
rect 13795 43872 13863 43928
rect 13919 43872 13987 43928
rect 14043 43872 14111 43928
rect 14167 43872 14235 43928
rect 14291 43872 14359 43928
rect 14415 43872 14483 43928
rect 14539 43872 14607 43928
rect 14663 43872 14673 43928
rect 12861 43804 14673 43872
rect 12861 43748 12871 43804
rect 12927 43748 12995 43804
rect 13051 43748 13119 43804
rect 13175 43748 13243 43804
rect 13299 43748 13367 43804
rect 13423 43748 13491 43804
rect 13547 43748 13615 43804
rect 13671 43748 13739 43804
rect 13795 43748 13863 43804
rect 13919 43748 13987 43804
rect 14043 43748 14111 43804
rect 14167 43748 14235 43804
rect 14291 43748 14359 43804
rect 14415 43748 14483 43804
rect 14539 43748 14607 43804
rect 14663 43748 14673 43804
rect 12861 43680 14673 43748
rect 12861 43624 12871 43680
rect 12927 43624 12995 43680
rect 13051 43624 13119 43680
rect 13175 43624 13243 43680
rect 13299 43624 13367 43680
rect 13423 43624 13491 43680
rect 13547 43624 13615 43680
rect 13671 43624 13739 43680
rect 13795 43624 13863 43680
rect 13919 43624 13987 43680
rect 14043 43624 14111 43680
rect 14167 43624 14235 43680
rect 14291 43624 14359 43680
rect 14415 43624 14483 43680
rect 14539 43624 14607 43680
rect 14663 43624 14673 43680
rect 12861 43556 14673 43624
rect 12861 43500 12871 43556
rect 12927 43500 12995 43556
rect 13051 43500 13119 43556
rect 13175 43500 13243 43556
rect 13299 43500 13367 43556
rect 13423 43500 13491 43556
rect 13547 43500 13615 43556
rect 13671 43500 13739 43556
rect 13795 43500 13863 43556
rect 13919 43500 13987 43556
rect 14043 43500 14111 43556
rect 14167 43500 14235 43556
rect 14291 43500 14359 43556
rect 14415 43500 14483 43556
rect 14539 43500 14607 43556
rect 14663 43500 14673 43556
rect 12861 43432 14673 43500
rect 12861 43376 12871 43432
rect 12927 43376 12995 43432
rect 13051 43376 13119 43432
rect 13175 43376 13243 43432
rect 13299 43376 13367 43432
rect 13423 43376 13491 43432
rect 13547 43376 13615 43432
rect 13671 43376 13739 43432
rect 13795 43376 13863 43432
rect 13919 43376 13987 43432
rect 14043 43376 14111 43432
rect 14167 43376 14235 43432
rect 14291 43376 14359 43432
rect 14415 43376 14483 43432
rect 14539 43376 14607 43432
rect 14663 43376 14673 43432
rect 12861 43308 14673 43376
rect 12861 43252 12871 43308
rect 12927 43252 12995 43308
rect 13051 43252 13119 43308
rect 13175 43252 13243 43308
rect 13299 43252 13367 43308
rect 13423 43252 13491 43308
rect 13547 43252 13615 43308
rect 13671 43252 13739 43308
rect 13795 43252 13863 43308
rect 13919 43252 13987 43308
rect 14043 43252 14111 43308
rect 14167 43252 14235 43308
rect 14291 43252 14359 43308
rect 14415 43252 14483 43308
rect 14539 43252 14607 43308
rect 14663 43252 14673 43308
rect 12861 43242 14673 43252
rect 2798 42948 4734 42958
rect 2798 42892 2808 42948
rect 2864 42892 2932 42948
rect 2988 42892 3056 42948
rect 3112 42892 3180 42948
rect 3236 42892 3304 42948
rect 3360 42892 3428 42948
rect 3484 42892 3552 42948
rect 3608 42892 3676 42948
rect 3732 42892 3800 42948
rect 3856 42892 3924 42948
rect 3980 42892 4048 42948
rect 4104 42892 4172 42948
rect 4228 42892 4296 42948
rect 4352 42892 4420 42948
rect 4476 42892 4544 42948
rect 4600 42892 4668 42948
rect 4724 42892 4734 42948
rect 2798 42824 4734 42892
rect 2798 42768 2808 42824
rect 2864 42768 2932 42824
rect 2988 42768 3056 42824
rect 3112 42768 3180 42824
rect 3236 42768 3304 42824
rect 3360 42768 3428 42824
rect 3484 42768 3552 42824
rect 3608 42768 3676 42824
rect 3732 42768 3800 42824
rect 3856 42768 3924 42824
rect 3980 42768 4048 42824
rect 4104 42768 4172 42824
rect 4228 42768 4296 42824
rect 4352 42768 4420 42824
rect 4476 42768 4544 42824
rect 4600 42768 4668 42824
rect 4724 42768 4734 42824
rect 2798 42700 4734 42768
rect 2798 42644 2808 42700
rect 2864 42644 2932 42700
rect 2988 42644 3056 42700
rect 3112 42644 3180 42700
rect 3236 42644 3304 42700
rect 3360 42644 3428 42700
rect 3484 42644 3552 42700
rect 3608 42644 3676 42700
rect 3732 42644 3800 42700
rect 3856 42644 3924 42700
rect 3980 42644 4048 42700
rect 4104 42644 4172 42700
rect 4228 42644 4296 42700
rect 4352 42644 4420 42700
rect 4476 42644 4544 42700
rect 4600 42644 4668 42700
rect 4724 42644 4734 42700
rect 2798 42576 4734 42644
rect 2798 42520 2808 42576
rect 2864 42520 2932 42576
rect 2988 42520 3056 42576
rect 3112 42520 3180 42576
rect 3236 42520 3304 42576
rect 3360 42520 3428 42576
rect 3484 42520 3552 42576
rect 3608 42520 3676 42576
rect 3732 42520 3800 42576
rect 3856 42520 3924 42576
rect 3980 42520 4048 42576
rect 4104 42520 4172 42576
rect 4228 42520 4296 42576
rect 4352 42520 4420 42576
rect 4476 42520 4544 42576
rect 4600 42520 4668 42576
rect 4724 42520 4734 42576
rect 2798 42452 4734 42520
rect 2798 42396 2808 42452
rect 2864 42396 2932 42452
rect 2988 42396 3056 42452
rect 3112 42396 3180 42452
rect 3236 42396 3304 42452
rect 3360 42396 3428 42452
rect 3484 42396 3552 42452
rect 3608 42396 3676 42452
rect 3732 42396 3800 42452
rect 3856 42396 3924 42452
rect 3980 42396 4048 42452
rect 4104 42396 4172 42452
rect 4228 42396 4296 42452
rect 4352 42396 4420 42452
rect 4476 42396 4544 42452
rect 4600 42396 4668 42452
rect 4724 42396 4734 42452
rect 2798 42328 4734 42396
rect 2798 42272 2808 42328
rect 2864 42272 2932 42328
rect 2988 42272 3056 42328
rect 3112 42272 3180 42328
rect 3236 42272 3304 42328
rect 3360 42272 3428 42328
rect 3484 42272 3552 42328
rect 3608 42272 3676 42328
rect 3732 42272 3800 42328
rect 3856 42272 3924 42328
rect 3980 42272 4048 42328
rect 4104 42272 4172 42328
rect 4228 42272 4296 42328
rect 4352 42272 4420 42328
rect 4476 42272 4544 42328
rect 4600 42272 4668 42328
rect 4724 42272 4734 42328
rect 2798 42204 4734 42272
rect 2798 42148 2808 42204
rect 2864 42148 2932 42204
rect 2988 42148 3056 42204
rect 3112 42148 3180 42204
rect 3236 42148 3304 42204
rect 3360 42148 3428 42204
rect 3484 42148 3552 42204
rect 3608 42148 3676 42204
rect 3732 42148 3800 42204
rect 3856 42148 3924 42204
rect 3980 42148 4048 42204
rect 4104 42148 4172 42204
rect 4228 42148 4296 42204
rect 4352 42148 4420 42204
rect 4476 42148 4544 42204
rect 4600 42148 4668 42204
rect 4724 42148 4734 42204
rect 2798 42080 4734 42148
rect 2798 42024 2808 42080
rect 2864 42024 2932 42080
rect 2988 42024 3056 42080
rect 3112 42024 3180 42080
rect 3236 42024 3304 42080
rect 3360 42024 3428 42080
rect 3484 42024 3552 42080
rect 3608 42024 3676 42080
rect 3732 42024 3800 42080
rect 3856 42024 3924 42080
rect 3980 42024 4048 42080
rect 4104 42024 4172 42080
rect 4228 42024 4296 42080
rect 4352 42024 4420 42080
rect 4476 42024 4544 42080
rect 4600 42024 4668 42080
rect 4724 42024 4734 42080
rect 2798 41956 4734 42024
rect 2798 41900 2808 41956
rect 2864 41900 2932 41956
rect 2988 41900 3056 41956
rect 3112 41900 3180 41956
rect 3236 41900 3304 41956
rect 3360 41900 3428 41956
rect 3484 41900 3552 41956
rect 3608 41900 3676 41956
rect 3732 41900 3800 41956
rect 3856 41900 3924 41956
rect 3980 41900 4048 41956
rect 4104 41900 4172 41956
rect 4228 41900 4296 41956
rect 4352 41900 4420 41956
rect 4476 41900 4544 41956
rect 4600 41900 4668 41956
rect 4724 41900 4734 41956
rect 2798 41832 4734 41900
rect 2798 41776 2808 41832
rect 2864 41776 2932 41832
rect 2988 41776 3056 41832
rect 3112 41776 3180 41832
rect 3236 41776 3304 41832
rect 3360 41776 3428 41832
rect 3484 41776 3552 41832
rect 3608 41776 3676 41832
rect 3732 41776 3800 41832
rect 3856 41776 3924 41832
rect 3980 41776 4048 41832
rect 4104 41776 4172 41832
rect 4228 41776 4296 41832
rect 4352 41776 4420 41832
rect 4476 41776 4544 41832
rect 4600 41776 4668 41832
rect 4724 41776 4734 41832
rect 2798 41708 4734 41776
rect 2798 41652 2808 41708
rect 2864 41652 2932 41708
rect 2988 41652 3056 41708
rect 3112 41652 3180 41708
rect 3236 41652 3304 41708
rect 3360 41652 3428 41708
rect 3484 41652 3552 41708
rect 3608 41652 3676 41708
rect 3732 41652 3800 41708
rect 3856 41652 3924 41708
rect 3980 41652 4048 41708
rect 4104 41652 4172 41708
rect 4228 41652 4296 41708
rect 4352 41652 4420 41708
rect 4476 41652 4544 41708
rect 4600 41652 4668 41708
rect 4724 41652 4734 41708
rect 2798 41642 4734 41652
rect 5168 42948 7104 42958
rect 5168 42892 5178 42948
rect 5234 42892 5302 42948
rect 5358 42892 5426 42948
rect 5482 42892 5550 42948
rect 5606 42892 5674 42948
rect 5730 42892 5798 42948
rect 5854 42892 5922 42948
rect 5978 42892 6046 42948
rect 6102 42892 6170 42948
rect 6226 42892 6294 42948
rect 6350 42892 6418 42948
rect 6474 42892 6542 42948
rect 6598 42892 6666 42948
rect 6722 42892 6790 42948
rect 6846 42892 6914 42948
rect 6970 42892 7038 42948
rect 7094 42892 7104 42948
rect 5168 42824 7104 42892
rect 5168 42768 5178 42824
rect 5234 42768 5302 42824
rect 5358 42768 5426 42824
rect 5482 42768 5550 42824
rect 5606 42768 5674 42824
rect 5730 42768 5798 42824
rect 5854 42768 5922 42824
rect 5978 42768 6046 42824
rect 6102 42768 6170 42824
rect 6226 42768 6294 42824
rect 6350 42768 6418 42824
rect 6474 42768 6542 42824
rect 6598 42768 6666 42824
rect 6722 42768 6790 42824
rect 6846 42768 6914 42824
rect 6970 42768 7038 42824
rect 7094 42768 7104 42824
rect 5168 42700 7104 42768
rect 5168 42644 5178 42700
rect 5234 42644 5302 42700
rect 5358 42644 5426 42700
rect 5482 42644 5550 42700
rect 5606 42644 5674 42700
rect 5730 42644 5798 42700
rect 5854 42644 5922 42700
rect 5978 42644 6046 42700
rect 6102 42644 6170 42700
rect 6226 42644 6294 42700
rect 6350 42644 6418 42700
rect 6474 42644 6542 42700
rect 6598 42644 6666 42700
rect 6722 42644 6790 42700
rect 6846 42644 6914 42700
rect 6970 42644 7038 42700
rect 7094 42644 7104 42700
rect 5168 42576 7104 42644
rect 5168 42520 5178 42576
rect 5234 42520 5302 42576
rect 5358 42520 5426 42576
rect 5482 42520 5550 42576
rect 5606 42520 5674 42576
rect 5730 42520 5798 42576
rect 5854 42520 5922 42576
rect 5978 42520 6046 42576
rect 6102 42520 6170 42576
rect 6226 42520 6294 42576
rect 6350 42520 6418 42576
rect 6474 42520 6542 42576
rect 6598 42520 6666 42576
rect 6722 42520 6790 42576
rect 6846 42520 6914 42576
rect 6970 42520 7038 42576
rect 7094 42520 7104 42576
rect 5168 42452 7104 42520
rect 5168 42396 5178 42452
rect 5234 42396 5302 42452
rect 5358 42396 5426 42452
rect 5482 42396 5550 42452
rect 5606 42396 5674 42452
rect 5730 42396 5798 42452
rect 5854 42396 5922 42452
rect 5978 42396 6046 42452
rect 6102 42396 6170 42452
rect 6226 42396 6294 42452
rect 6350 42396 6418 42452
rect 6474 42396 6542 42452
rect 6598 42396 6666 42452
rect 6722 42396 6790 42452
rect 6846 42396 6914 42452
rect 6970 42396 7038 42452
rect 7094 42396 7104 42452
rect 5168 42328 7104 42396
rect 5168 42272 5178 42328
rect 5234 42272 5302 42328
rect 5358 42272 5426 42328
rect 5482 42272 5550 42328
rect 5606 42272 5674 42328
rect 5730 42272 5798 42328
rect 5854 42272 5922 42328
rect 5978 42272 6046 42328
rect 6102 42272 6170 42328
rect 6226 42272 6294 42328
rect 6350 42272 6418 42328
rect 6474 42272 6542 42328
rect 6598 42272 6666 42328
rect 6722 42272 6790 42328
rect 6846 42272 6914 42328
rect 6970 42272 7038 42328
rect 7094 42272 7104 42328
rect 5168 42204 7104 42272
rect 5168 42148 5178 42204
rect 5234 42148 5302 42204
rect 5358 42148 5426 42204
rect 5482 42148 5550 42204
rect 5606 42148 5674 42204
rect 5730 42148 5798 42204
rect 5854 42148 5922 42204
rect 5978 42148 6046 42204
rect 6102 42148 6170 42204
rect 6226 42148 6294 42204
rect 6350 42148 6418 42204
rect 6474 42148 6542 42204
rect 6598 42148 6666 42204
rect 6722 42148 6790 42204
rect 6846 42148 6914 42204
rect 6970 42148 7038 42204
rect 7094 42148 7104 42204
rect 5168 42080 7104 42148
rect 5168 42024 5178 42080
rect 5234 42024 5302 42080
rect 5358 42024 5426 42080
rect 5482 42024 5550 42080
rect 5606 42024 5674 42080
rect 5730 42024 5798 42080
rect 5854 42024 5922 42080
rect 5978 42024 6046 42080
rect 6102 42024 6170 42080
rect 6226 42024 6294 42080
rect 6350 42024 6418 42080
rect 6474 42024 6542 42080
rect 6598 42024 6666 42080
rect 6722 42024 6790 42080
rect 6846 42024 6914 42080
rect 6970 42024 7038 42080
rect 7094 42024 7104 42080
rect 5168 41956 7104 42024
rect 5168 41900 5178 41956
rect 5234 41900 5302 41956
rect 5358 41900 5426 41956
rect 5482 41900 5550 41956
rect 5606 41900 5674 41956
rect 5730 41900 5798 41956
rect 5854 41900 5922 41956
rect 5978 41900 6046 41956
rect 6102 41900 6170 41956
rect 6226 41900 6294 41956
rect 6350 41900 6418 41956
rect 6474 41900 6542 41956
rect 6598 41900 6666 41956
rect 6722 41900 6790 41956
rect 6846 41900 6914 41956
rect 6970 41900 7038 41956
rect 7094 41900 7104 41956
rect 5168 41832 7104 41900
rect 5168 41776 5178 41832
rect 5234 41776 5302 41832
rect 5358 41776 5426 41832
rect 5482 41776 5550 41832
rect 5606 41776 5674 41832
rect 5730 41776 5798 41832
rect 5854 41776 5922 41832
rect 5978 41776 6046 41832
rect 6102 41776 6170 41832
rect 6226 41776 6294 41832
rect 6350 41776 6418 41832
rect 6474 41776 6542 41832
rect 6598 41776 6666 41832
rect 6722 41776 6790 41832
rect 6846 41776 6914 41832
rect 6970 41776 7038 41832
rect 7094 41776 7104 41832
rect 5168 41708 7104 41776
rect 5168 41652 5178 41708
rect 5234 41652 5302 41708
rect 5358 41652 5426 41708
rect 5482 41652 5550 41708
rect 5606 41652 5674 41708
rect 5730 41652 5798 41708
rect 5854 41652 5922 41708
rect 5978 41652 6046 41708
rect 6102 41652 6170 41708
rect 6226 41652 6294 41708
rect 6350 41652 6418 41708
rect 6474 41652 6542 41708
rect 6598 41652 6666 41708
rect 6722 41652 6790 41708
rect 6846 41652 6914 41708
rect 6970 41652 7038 41708
rect 7094 41652 7104 41708
rect 5168 41642 7104 41652
rect 7874 42948 9810 42958
rect 7874 42892 7884 42948
rect 7940 42892 8008 42948
rect 8064 42892 8132 42948
rect 8188 42892 8256 42948
rect 8312 42892 8380 42948
rect 8436 42892 8504 42948
rect 8560 42892 8628 42948
rect 8684 42892 8752 42948
rect 8808 42892 8876 42948
rect 8932 42892 9000 42948
rect 9056 42892 9124 42948
rect 9180 42892 9248 42948
rect 9304 42892 9372 42948
rect 9428 42892 9496 42948
rect 9552 42892 9620 42948
rect 9676 42892 9744 42948
rect 9800 42892 9810 42948
rect 7874 42824 9810 42892
rect 7874 42768 7884 42824
rect 7940 42768 8008 42824
rect 8064 42768 8132 42824
rect 8188 42768 8256 42824
rect 8312 42768 8380 42824
rect 8436 42768 8504 42824
rect 8560 42768 8628 42824
rect 8684 42768 8752 42824
rect 8808 42768 8876 42824
rect 8932 42768 9000 42824
rect 9056 42768 9124 42824
rect 9180 42768 9248 42824
rect 9304 42768 9372 42824
rect 9428 42768 9496 42824
rect 9552 42768 9620 42824
rect 9676 42768 9744 42824
rect 9800 42768 9810 42824
rect 7874 42700 9810 42768
rect 7874 42644 7884 42700
rect 7940 42644 8008 42700
rect 8064 42644 8132 42700
rect 8188 42644 8256 42700
rect 8312 42644 8380 42700
rect 8436 42644 8504 42700
rect 8560 42644 8628 42700
rect 8684 42644 8752 42700
rect 8808 42644 8876 42700
rect 8932 42644 9000 42700
rect 9056 42644 9124 42700
rect 9180 42644 9248 42700
rect 9304 42644 9372 42700
rect 9428 42644 9496 42700
rect 9552 42644 9620 42700
rect 9676 42644 9744 42700
rect 9800 42644 9810 42700
rect 7874 42576 9810 42644
rect 7874 42520 7884 42576
rect 7940 42520 8008 42576
rect 8064 42520 8132 42576
rect 8188 42520 8256 42576
rect 8312 42520 8380 42576
rect 8436 42520 8504 42576
rect 8560 42520 8628 42576
rect 8684 42520 8752 42576
rect 8808 42520 8876 42576
rect 8932 42520 9000 42576
rect 9056 42520 9124 42576
rect 9180 42520 9248 42576
rect 9304 42520 9372 42576
rect 9428 42520 9496 42576
rect 9552 42520 9620 42576
rect 9676 42520 9744 42576
rect 9800 42520 9810 42576
rect 7874 42452 9810 42520
rect 7874 42396 7884 42452
rect 7940 42396 8008 42452
rect 8064 42396 8132 42452
rect 8188 42396 8256 42452
rect 8312 42396 8380 42452
rect 8436 42396 8504 42452
rect 8560 42396 8628 42452
rect 8684 42396 8752 42452
rect 8808 42396 8876 42452
rect 8932 42396 9000 42452
rect 9056 42396 9124 42452
rect 9180 42396 9248 42452
rect 9304 42396 9372 42452
rect 9428 42396 9496 42452
rect 9552 42396 9620 42452
rect 9676 42396 9744 42452
rect 9800 42396 9810 42452
rect 7874 42328 9810 42396
rect 7874 42272 7884 42328
rect 7940 42272 8008 42328
rect 8064 42272 8132 42328
rect 8188 42272 8256 42328
rect 8312 42272 8380 42328
rect 8436 42272 8504 42328
rect 8560 42272 8628 42328
rect 8684 42272 8752 42328
rect 8808 42272 8876 42328
rect 8932 42272 9000 42328
rect 9056 42272 9124 42328
rect 9180 42272 9248 42328
rect 9304 42272 9372 42328
rect 9428 42272 9496 42328
rect 9552 42272 9620 42328
rect 9676 42272 9744 42328
rect 9800 42272 9810 42328
rect 7874 42204 9810 42272
rect 7874 42148 7884 42204
rect 7940 42148 8008 42204
rect 8064 42148 8132 42204
rect 8188 42148 8256 42204
rect 8312 42148 8380 42204
rect 8436 42148 8504 42204
rect 8560 42148 8628 42204
rect 8684 42148 8752 42204
rect 8808 42148 8876 42204
rect 8932 42148 9000 42204
rect 9056 42148 9124 42204
rect 9180 42148 9248 42204
rect 9304 42148 9372 42204
rect 9428 42148 9496 42204
rect 9552 42148 9620 42204
rect 9676 42148 9744 42204
rect 9800 42148 9810 42204
rect 7874 42080 9810 42148
rect 7874 42024 7884 42080
rect 7940 42024 8008 42080
rect 8064 42024 8132 42080
rect 8188 42024 8256 42080
rect 8312 42024 8380 42080
rect 8436 42024 8504 42080
rect 8560 42024 8628 42080
rect 8684 42024 8752 42080
rect 8808 42024 8876 42080
rect 8932 42024 9000 42080
rect 9056 42024 9124 42080
rect 9180 42024 9248 42080
rect 9304 42024 9372 42080
rect 9428 42024 9496 42080
rect 9552 42024 9620 42080
rect 9676 42024 9744 42080
rect 9800 42024 9810 42080
rect 7874 41956 9810 42024
rect 7874 41900 7884 41956
rect 7940 41900 8008 41956
rect 8064 41900 8132 41956
rect 8188 41900 8256 41956
rect 8312 41900 8380 41956
rect 8436 41900 8504 41956
rect 8560 41900 8628 41956
rect 8684 41900 8752 41956
rect 8808 41900 8876 41956
rect 8932 41900 9000 41956
rect 9056 41900 9124 41956
rect 9180 41900 9248 41956
rect 9304 41900 9372 41956
rect 9428 41900 9496 41956
rect 9552 41900 9620 41956
rect 9676 41900 9744 41956
rect 9800 41900 9810 41956
rect 7874 41832 9810 41900
rect 7874 41776 7884 41832
rect 7940 41776 8008 41832
rect 8064 41776 8132 41832
rect 8188 41776 8256 41832
rect 8312 41776 8380 41832
rect 8436 41776 8504 41832
rect 8560 41776 8628 41832
rect 8684 41776 8752 41832
rect 8808 41776 8876 41832
rect 8932 41776 9000 41832
rect 9056 41776 9124 41832
rect 9180 41776 9248 41832
rect 9304 41776 9372 41832
rect 9428 41776 9496 41832
rect 9552 41776 9620 41832
rect 9676 41776 9744 41832
rect 9800 41776 9810 41832
rect 7874 41708 9810 41776
rect 7874 41652 7884 41708
rect 7940 41652 8008 41708
rect 8064 41652 8132 41708
rect 8188 41652 8256 41708
rect 8312 41652 8380 41708
rect 8436 41652 8504 41708
rect 8560 41652 8628 41708
rect 8684 41652 8752 41708
rect 8808 41652 8876 41708
rect 8932 41652 9000 41708
rect 9056 41652 9124 41708
rect 9180 41652 9248 41708
rect 9304 41652 9372 41708
rect 9428 41652 9496 41708
rect 9552 41652 9620 41708
rect 9676 41652 9744 41708
rect 9800 41652 9810 41708
rect 7874 41642 9810 41652
rect 10244 42948 12180 42958
rect 10244 42892 10254 42948
rect 10310 42892 10378 42948
rect 10434 42892 10502 42948
rect 10558 42892 10626 42948
rect 10682 42892 10750 42948
rect 10806 42892 10874 42948
rect 10930 42892 10998 42948
rect 11054 42892 11122 42948
rect 11178 42892 11246 42948
rect 11302 42892 11370 42948
rect 11426 42892 11494 42948
rect 11550 42892 11618 42948
rect 11674 42892 11742 42948
rect 11798 42892 11866 42948
rect 11922 42892 11990 42948
rect 12046 42892 12114 42948
rect 12170 42892 12180 42948
rect 10244 42824 12180 42892
rect 10244 42768 10254 42824
rect 10310 42768 10378 42824
rect 10434 42768 10502 42824
rect 10558 42768 10626 42824
rect 10682 42768 10750 42824
rect 10806 42768 10874 42824
rect 10930 42768 10998 42824
rect 11054 42768 11122 42824
rect 11178 42768 11246 42824
rect 11302 42768 11370 42824
rect 11426 42768 11494 42824
rect 11550 42768 11618 42824
rect 11674 42768 11742 42824
rect 11798 42768 11866 42824
rect 11922 42768 11990 42824
rect 12046 42768 12114 42824
rect 12170 42768 12180 42824
rect 10244 42700 12180 42768
rect 10244 42644 10254 42700
rect 10310 42644 10378 42700
rect 10434 42644 10502 42700
rect 10558 42644 10626 42700
rect 10682 42644 10750 42700
rect 10806 42644 10874 42700
rect 10930 42644 10998 42700
rect 11054 42644 11122 42700
rect 11178 42644 11246 42700
rect 11302 42644 11370 42700
rect 11426 42644 11494 42700
rect 11550 42644 11618 42700
rect 11674 42644 11742 42700
rect 11798 42644 11866 42700
rect 11922 42644 11990 42700
rect 12046 42644 12114 42700
rect 12170 42644 12180 42700
rect 10244 42576 12180 42644
rect 10244 42520 10254 42576
rect 10310 42520 10378 42576
rect 10434 42520 10502 42576
rect 10558 42520 10626 42576
rect 10682 42520 10750 42576
rect 10806 42520 10874 42576
rect 10930 42520 10998 42576
rect 11054 42520 11122 42576
rect 11178 42520 11246 42576
rect 11302 42520 11370 42576
rect 11426 42520 11494 42576
rect 11550 42520 11618 42576
rect 11674 42520 11742 42576
rect 11798 42520 11866 42576
rect 11922 42520 11990 42576
rect 12046 42520 12114 42576
rect 12170 42520 12180 42576
rect 10244 42452 12180 42520
rect 10244 42396 10254 42452
rect 10310 42396 10378 42452
rect 10434 42396 10502 42452
rect 10558 42396 10626 42452
rect 10682 42396 10750 42452
rect 10806 42396 10874 42452
rect 10930 42396 10998 42452
rect 11054 42396 11122 42452
rect 11178 42396 11246 42452
rect 11302 42396 11370 42452
rect 11426 42396 11494 42452
rect 11550 42396 11618 42452
rect 11674 42396 11742 42452
rect 11798 42396 11866 42452
rect 11922 42396 11990 42452
rect 12046 42396 12114 42452
rect 12170 42396 12180 42452
rect 10244 42328 12180 42396
rect 10244 42272 10254 42328
rect 10310 42272 10378 42328
rect 10434 42272 10502 42328
rect 10558 42272 10626 42328
rect 10682 42272 10750 42328
rect 10806 42272 10874 42328
rect 10930 42272 10998 42328
rect 11054 42272 11122 42328
rect 11178 42272 11246 42328
rect 11302 42272 11370 42328
rect 11426 42272 11494 42328
rect 11550 42272 11618 42328
rect 11674 42272 11742 42328
rect 11798 42272 11866 42328
rect 11922 42272 11990 42328
rect 12046 42272 12114 42328
rect 12170 42272 12180 42328
rect 10244 42204 12180 42272
rect 10244 42148 10254 42204
rect 10310 42148 10378 42204
rect 10434 42148 10502 42204
rect 10558 42148 10626 42204
rect 10682 42148 10750 42204
rect 10806 42148 10874 42204
rect 10930 42148 10998 42204
rect 11054 42148 11122 42204
rect 11178 42148 11246 42204
rect 11302 42148 11370 42204
rect 11426 42148 11494 42204
rect 11550 42148 11618 42204
rect 11674 42148 11742 42204
rect 11798 42148 11866 42204
rect 11922 42148 11990 42204
rect 12046 42148 12114 42204
rect 12170 42148 12180 42204
rect 10244 42080 12180 42148
rect 10244 42024 10254 42080
rect 10310 42024 10378 42080
rect 10434 42024 10502 42080
rect 10558 42024 10626 42080
rect 10682 42024 10750 42080
rect 10806 42024 10874 42080
rect 10930 42024 10998 42080
rect 11054 42024 11122 42080
rect 11178 42024 11246 42080
rect 11302 42024 11370 42080
rect 11426 42024 11494 42080
rect 11550 42024 11618 42080
rect 11674 42024 11742 42080
rect 11798 42024 11866 42080
rect 11922 42024 11990 42080
rect 12046 42024 12114 42080
rect 12170 42024 12180 42080
rect 10244 41956 12180 42024
rect 10244 41900 10254 41956
rect 10310 41900 10378 41956
rect 10434 41900 10502 41956
rect 10558 41900 10626 41956
rect 10682 41900 10750 41956
rect 10806 41900 10874 41956
rect 10930 41900 10998 41956
rect 11054 41900 11122 41956
rect 11178 41900 11246 41956
rect 11302 41900 11370 41956
rect 11426 41900 11494 41956
rect 11550 41900 11618 41956
rect 11674 41900 11742 41956
rect 11798 41900 11866 41956
rect 11922 41900 11990 41956
rect 12046 41900 12114 41956
rect 12170 41900 12180 41956
rect 10244 41832 12180 41900
rect 10244 41776 10254 41832
rect 10310 41776 10378 41832
rect 10434 41776 10502 41832
rect 10558 41776 10626 41832
rect 10682 41776 10750 41832
rect 10806 41776 10874 41832
rect 10930 41776 10998 41832
rect 11054 41776 11122 41832
rect 11178 41776 11246 41832
rect 11302 41776 11370 41832
rect 11426 41776 11494 41832
rect 11550 41776 11618 41832
rect 11674 41776 11742 41832
rect 11798 41776 11866 41832
rect 11922 41776 11990 41832
rect 12046 41776 12114 41832
rect 12170 41776 12180 41832
rect 10244 41708 12180 41776
rect 10244 41652 10254 41708
rect 10310 41652 10378 41708
rect 10434 41652 10502 41708
rect 10558 41652 10626 41708
rect 10682 41652 10750 41708
rect 10806 41652 10874 41708
rect 10930 41652 10998 41708
rect 11054 41652 11122 41708
rect 11178 41652 11246 41708
rect 11302 41652 11370 41708
rect 11426 41652 11494 41708
rect 11550 41652 11618 41708
rect 11674 41652 11742 41708
rect 11798 41652 11866 41708
rect 11922 41652 11990 41708
rect 12046 41652 12114 41708
rect 12170 41652 12180 41708
rect 10244 41642 12180 41652
rect 12861 42948 14673 42958
rect 12861 42892 12871 42948
rect 12927 42892 12995 42948
rect 13051 42892 13119 42948
rect 13175 42892 13243 42948
rect 13299 42892 13367 42948
rect 13423 42892 13491 42948
rect 13547 42892 13615 42948
rect 13671 42892 13739 42948
rect 13795 42892 13863 42948
rect 13919 42892 13987 42948
rect 14043 42892 14111 42948
rect 14167 42892 14235 42948
rect 14291 42892 14359 42948
rect 14415 42892 14483 42948
rect 14539 42892 14607 42948
rect 14663 42892 14673 42948
rect 12861 42824 14673 42892
rect 12861 42768 12871 42824
rect 12927 42768 12995 42824
rect 13051 42768 13119 42824
rect 13175 42768 13243 42824
rect 13299 42768 13367 42824
rect 13423 42768 13491 42824
rect 13547 42768 13615 42824
rect 13671 42768 13739 42824
rect 13795 42768 13863 42824
rect 13919 42768 13987 42824
rect 14043 42768 14111 42824
rect 14167 42768 14235 42824
rect 14291 42768 14359 42824
rect 14415 42768 14483 42824
rect 14539 42768 14607 42824
rect 14663 42768 14673 42824
rect 12861 42700 14673 42768
rect 12861 42644 12871 42700
rect 12927 42644 12995 42700
rect 13051 42644 13119 42700
rect 13175 42644 13243 42700
rect 13299 42644 13367 42700
rect 13423 42644 13491 42700
rect 13547 42644 13615 42700
rect 13671 42644 13739 42700
rect 13795 42644 13863 42700
rect 13919 42644 13987 42700
rect 14043 42644 14111 42700
rect 14167 42644 14235 42700
rect 14291 42644 14359 42700
rect 14415 42644 14483 42700
rect 14539 42644 14607 42700
rect 14663 42644 14673 42700
rect 12861 42576 14673 42644
rect 12861 42520 12871 42576
rect 12927 42520 12995 42576
rect 13051 42520 13119 42576
rect 13175 42520 13243 42576
rect 13299 42520 13367 42576
rect 13423 42520 13491 42576
rect 13547 42520 13615 42576
rect 13671 42520 13739 42576
rect 13795 42520 13863 42576
rect 13919 42520 13987 42576
rect 14043 42520 14111 42576
rect 14167 42520 14235 42576
rect 14291 42520 14359 42576
rect 14415 42520 14483 42576
rect 14539 42520 14607 42576
rect 14663 42520 14673 42576
rect 12861 42452 14673 42520
rect 12861 42396 12871 42452
rect 12927 42396 12995 42452
rect 13051 42396 13119 42452
rect 13175 42396 13243 42452
rect 13299 42396 13367 42452
rect 13423 42396 13491 42452
rect 13547 42396 13615 42452
rect 13671 42396 13739 42452
rect 13795 42396 13863 42452
rect 13919 42396 13987 42452
rect 14043 42396 14111 42452
rect 14167 42396 14235 42452
rect 14291 42396 14359 42452
rect 14415 42396 14483 42452
rect 14539 42396 14607 42452
rect 14663 42396 14673 42452
rect 12861 42328 14673 42396
rect 12861 42272 12871 42328
rect 12927 42272 12995 42328
rect 13051 42272 13119 42328
rect 13175 42272 13243 42328
rect 13299 42272 13367 42328
rect 13423 42272 13491 42328
rect 13547 42272 13615 42328
rect 13671 42272 13739 42328
rect 13795 42272 13863 42328
rect 13919 42272 13987 42328
rect 14043 42272 14111 42328
rect 14167 42272 14235 42328
rect 14291 42272 14359 42328
rect 14415 42272 14483 42328
rect 14539 42272 14607 42328
rect 14663 42272 14673 42328
rect 12861 42204 14673 42272
rect 12861 42148 12871 42204
rect 12927 42148 12995 42204
rect 13051 42148 13119 42204
rect 13175 42148 13243 42204
rect 13299 42148 13367 42204
rect 13423 42148 13491 42204
rect 13547 42148 13615 42204
rect 13671 42148 13739 42204
rect 13795 42148 13863 42204
rect 13919 42148 13987 42204
rect 14043 42148 14111 42204
rect 14167 42148 14235 42204
rect 14291 42148 14359 42204
rect 14415 42148 14483 42204
rect 14539 42148 14607 42204
rect 14663 42148 14673 42204
rect 12861 42080 14673 42148
rect 12861 42024 12871 42080
rect 12927 42024 12995 42080
rect 13051 42024 13119 42080
rect 13175 42024 13243 42080
rect 13299 42024 13367 42080
rect 13423 42024 13491 42080
rect 13547 42024 13615 42080
rect 13671 42024 13739 42080
rect 13795 42024 13863 42080
rect 13919 42024 13987 42080
rect 14043 42024 14111 42080
rect 14167 42024 14235 42080
rect 14291 42024 14359 42080
rect 14415 42024 14483 42080
rect 14539 42024 14607 42080
rect 14663 42024 14673 42080
rect 12861 41956 14673 42024
rect 12861 41900 12871 41956
rect 12927 41900 12995 41956
rect 13051 41900 13119 41956
rect 13175 41900 13243 41956
rect 13299 41900 13367 41956
rect 13423 41900 13491 41956
rect 13547 41900 13615 41956
rect 13671 41900 13739 41956
rect 13795 41900 13863 41956
rect 13919 41900 13987 41956
rect 14043 41900 14111 41956
rect 14167 41900 14235 41956
rect 14291 41900 14359 41956
rect 14415 41900 14483 41956
rect 14539 41900 14607 41956
rect 14663 41900 14673 41956
rect 12861 41832 14673 41900
rect 12861 41776 12871 41832
rect 12927 41776 12995 41832
rect 13051 41776 13119 41832
rect 13175 41776 13243 41832
rect 13299 41776 13367 41832
rect 13423 41776 13491 41832
rect 13547 41776 13615 41832
rect 13671 41776 13739 41832
rect 13795 41776 13863 41832
rect 13919 41776 13987 41832
rect 14043 41776 14111 41832
rect 14167 41776 14235 41832
rect 14291 41776 14359 41832
rect 14415 41776 14483 41832
rect 14539 41776 14607 41832
rect 14663 41776 14673 41832
rect 12861 41708 14673 41776
rect 12861 41652 12871 41708
rect 12927 41652 12995 41708
rect 13051 41652 13119 41708
rect 13175 41652 13243 41708
rect 13299 41652 13367 41708
rect 13423 41652 13491 41708
rect 13547 41652 13615 41708
rect 13671 41652 13739 41708
rect 13795 41652 13863 41708
rect 13919 41652 13987 41708
rect 14043 41652 14111 41708
rect 14167 41652 14235 41708
rect 14291 41652 14359 41708
rect 14415 41652 14483 41708
rect 14539 41652 14607 41708
rect 14663 41652 14673 41708
rect 12861 41642 14673 41652
rect 2798 41348 4734 41358
rect 2798 41292 2808 41348
rect 2864 41292 2932 41348
rect 2988 41292 3056 41348
rect 3112 41292 3180 41348
rect 3236 41292 3304 41348
rect 3360 41292 3428 41348
rect 3484 41292 3552 41348
rect 3608 41292 3676 41348
rect 3732 41292 3800 41348
rect 3856 41292 3924 41348
rect 3980 41292 4048 41348
rect 4104 41292 4172 41348
rect 4228 41292 4296 41348
rect 4352 41292 4420 41348
rect 4476 41292 4544 41348
rect 4600 41292 4668 41348
rect 4724 41292 4734 41348
rect 2798 41224 4734 41292
rect 2798 41168 2808 41224
rect 2864 41168 2932 41224
rect 2988 41168 3056 41224
rect 3112 41168 3180 41224
rect 3236 41168 3304 41224
rect 3360 41168 3428 41224
rect 3484 41168 3552 41224
rect 3608 41168 3676 41224
rect 3732 41168 3800 41224
rect 3856 41168 3924 41224
rect 3980 41168 4048 41224
rect 4104 41168 4172 41224
rect 4228 41168 4296 41224
rect 4352 41168 4420 41224
rect 4476 41168 4544 41224
rect 4600 41168 4668 41224
rect 4724 41168 4734 41224
rect 2798 41100 4734 41168
rect 2798 41044 2808 41100
rect 2864 41044 2932 41100
rect 2988 41044 3056 41100
rect 3112 41044 3180 41100
rect 3236 41044 3304 41100
rect 3360 41044 3428 41100
rect 3484 41044 3552 41100
rect 3608 41044 3676 41100
rect 3732 41044 3800 41100
rect 3856 41044 3924 41100
rect 3980 41044 4048 41100
rect 4104 41044 4172 41100
rect 4228 41044 4296 41100
rect 4352 41044 4420 41100
rect 4476 41044 4544 41100
rect 4600 41044 4668 41100
rect 4724 41044 4734 41100
rect 2798 40976 4734 41044
rect 2798 40920 2808 40976
rect 2864 40920 2932 40976
rect 2988 40920 3056 40976
rect 3112 40920 3180 40976
rect 3236 40920 3304 40976
rect 3360 40920 3428 40976
rect 3484 40920 3552 40976
rect 3608 40920 3676 40976
rect 3732 40920 3800 40976
rect 3856 40920 3924 40976
rect 3980 40920 4048 40976
rect 4104 40920 4172 40976
rect 4228 40920 4296 40976
rect 4352 40920 4420 40976
rect 4476 40920 4544 40976
rect 4600 40920 4668 40976
rect 4724 40920 4734 40976
rect 2798 40852 4734 40920
rect 2798 40796 2808 40852
rect 2864 40796 2932 40852
rect 2988 40796 3056 40852
rect 3112 40796 3180 40852
rect 3236 40796 3304 40852
rect 3360 40796 3428 40852
rect 3484 40796 3552 40852
rect 3608 40796 3676 40852
rect 3732 40796 3800 40852
rect 3856 40796 3924 40852
rect 3980 40796 4048 40852
rect 4104 40796 4172 40852
rect 4228 40796 4296 40852
rect 4352 40796 4420 40852
rect 4476 40796 4544 40852
rect 4600 40796 4668 40852
rect 4724 40796 4734 40852
rect 2798 40728 4734 40796
rect 2798 40672 2808 40728
rect 2864 40672 2932 40728
rect 2988 40672 3056 40728
rect 3112 40672 3180 40728
rect 3236 40672 3304 40728
rect 3360 40672 3428 40728
rect 3484 40672 3552 40728
rect 3608 40672 3676 40728
rect 3732 40672 3800 40728
rect 3856 40672 3924 40728
rect 3980 40672 4048 40728
rect 4104 40672 4172 40728
rect 4228 40672 4296 40728
rect 4352 40672 4420 40728
rect 4476 40672 4544 40728
rect 4600 40672 4668 40728
rect 4724 40672 4734 40728
rect 2798 40604 4734 40672
rect 2798 40548 2808 40604
rect 2864 40548 2932 40604
rect 2988 40548 3056 40604
rect 3112 40548 3180 40604
rect 3236 40548 3304 40604
rect 3360 40548 3428 40604
rect 3484 40548 3552 40604
rect 3608 40548 3676 40604
rect 3732 40548 3800 40604
rect 3856 40548 3924 40604
rect 3980 40548 4048 40604
rect 4104 40548 4172 40604
rect 4228 40548 4296 40604
rect 4352 40548 4420 40604
rect 4476 40548 4544 40604
rect 4600 40548 4668 40604
rect 4724 40548 4734 40604
rect 2798 40480 4734 40548
rect 2798 40424 2808 40480
rect 2864 40424 2932 40480
rect 2988 40424 3056 40480
rect 3112 40424 3180 40480
rect 3236 40424 3304 40480
rect 3360 40424 3428 40480
rect 3484 40424 3552 40480
rect 3608 40424 3676 40480
rect 3732 40424 3800 40480
rect 3856 40424 3924 40480
rect 3980 40424 4048 40480
rect 4104 40424 4172 40480
rect 4228 40424 4296 40480
rect 4352 40424 4420 40480
rect 4476 40424 4544 40480
rect 4600 40424 4668 40480
rect 4724 40424 4734 40480
rect 2798 40356 4734 40424
rect 2798 40300 2808 40356
rect 2864 40300 2932 40356
rect 2988 40300 3056 40356
rect 3112 40300 3180 40356
rect 3236 40300 3304 40356
rect 3360 40300 3428 40356
rect 3484 40300 3552 40356
rect 3608 40300 3676 40356
rect 3732 40300 3800 40356
rect 3856 40300 3924 40356
rect 3980 40300 4048 40356
rect 4104 40300 4172 40356
rect 4228 40300 4296 40356
rect 4352 40300 4420 40356
rect 4476 40300 4544 40356
rect 4600 40300 4668 40356
rect 4724 40300 4734 40356
rect 2798 40232 4734 40300
rect 2798 40176 2808 40232
rect 2864 40176 2932 40232
rect 2988 40176 3056 40232
rect 3112 40176 3180 40232
rect 3236 40176 3304 40232
rect 3360 40176 3428 40232
rect 3484 40176 3552 40232
rect 3608 40176 3676 40232
rect 3732 40176 3800 40232
rect 3856 40176 3924 40232
rect 3980 40176 4048 40232
rect 4104 40176 4172 40232
rect 4228 40176 4296 40232
rect 4352 40176 4420 40232
rect 4476 40176 4544 40232
rect 4600 40176 4668 40232
rect 4724 40176 4734 40232
rect 2798 40108 4734 40176
rect 2798 40052 2808 40108
rect 2864 40052 2932 40108
rect 2988 40052 3056 40108
rect 3112 40052 3180 40108
rect 3236 40052 3304 40108
rect 3360 40052 3428 40108
rect 3484 40052 3552 40108
rect 3608 40052 3676 40108
rect 3732 40052 3800 40108
rect 3856 40052 3924 40108
rect 3980 40052 4048 40108
rect 4104 40052 4172 40108
rect 4228 40052 4296 40108
rect 4352 40052 4420 40108
rect 4476 40052 4544 40108
rect 4600 40052 4668 40108
rect 4724 40052 4734 40108
rect 2798 40042 4734 40052
rect 5168 41348 7104 41358
rect 5168 41292 5178 41348
rect 5234 41292 5302 41348
rect 5358 41292 5426 41348
rect 5482 41292 5550 41348
rect 5606 41292 5674 41348
rect 5730 41292 5798 41348
rect 5854 41292 5922 41348
rect 5978 41292 6046 41348
rect 6102 41292 6170 41348
rect 6226 41292 6294 41348
rect 6350 41292 6418 41348
rect 6474 41292 6542 41348
rect 6598 41292 6666 41348
rect 6722 41292 6790 41348
rect 6846 41292 6914 41348
rect 6970 41292 7038 41348
rect 7094 41292 7104 41348
rect 5168 41224 7104 41292
rect 5168 41168 5178 41224
rect 5234 41168 5302 41224
rect 5358 41168 5426 41224
rect 5482 41168 5550 41224
rect 5606 41168 5674 41224
rect 5730 41168 5798 41224
rect 5854 41168 5922 41224
rect 5978 41168 6046 41224
rect 6102 41168 6170 41224
rect 6226 41168 6294 41224
rect 6350 41168 6418 41224
rect 6474 41168 6542 41224
rect 6598 41168 6666 41224
rect 6722 41168 6790 41224
rect 6846 41168 6914 41224
rect 6970 41168 7038 41224
rect 7094 41168 7104 41224
rect 5168 41100 7104 41168
rect 5168 41044 5178 41100
rect 5234 41044 5302 41100
rect 5358 41044 5426 41100
rect 5482 41044 5550 41100
rect 5606 41044 5674 41100
rect 5730 41044 5798 41100
rect 5854 41044 5922 41100
rect 5978 41044 6046 41100
rect 6102 41044 6170 41100
rect 6226 41044 6294 41100
rect 6350 41044 6418 41100
rect 6474 41044 6542 41100
rect 6598 41044 6666 41100
rect 6722 41044 6790 41100
rect 6846 41044 6914 41100
rect 6970 41044 7038 41100
rect 7094 41044 7104 41100
rect 5168 40976 7104 41044
rect 5168 40920 5178 40976
rect 5234 40920 5302 40976
rect 5358 40920 5426 40976
rect 5482 40920 5550 40976
rect 5606 40920 5674 40976
rect 5730 40920 5798 40976
rect 5854 40920 5922 40976
rect 5978 40920 6046 40976
rect 6102 40920 6170 40976
rect 6226 40920 6294 40976
rect 6350 40920 6418 40976
rect 6474 40920 6542 40976
rect 6598 40920 6666 40976
rect 6722 40920 6790 40976
rect 6846 40920 6914 40976
rect 6970 40920 7038 40976
rect 7094 40920 7104 40976
rect 5168 40852 7104 40920
rect 5168 40796 5178 40852
rect 5234 40796 5302 40852
rect 5358 40796 5426 40852
rect 5482 40796 5550 40852
rect 5606 40796 5674 40852
rect 5730 40796 5798 40852
rect 5854 40796 5922 40852
rect 5978 40796 6046 40852
rect 6102 40796 6170 40852
rect 6226 40796 6294 40852
rect 6350 40796 6418 40852
rect 6474 40796 6542 40852
rect 6598 40796 6666 40852
rect 6722 40796 6790 40852
rect 6846 40796 6914 40852
rect 6970 40796 7038 40852
rect 7094 40796 7104 40852
rect 5168 40728 7104 40796
rect 5168 40672 5178 40728
rect 5234 40672 5302 40728
rect 5358 40672 5426 40728
rect 5482 40672 5550 40728
rect 5606 40672 5674 40728
rect 5730 40672 5798 40728
rect 5854 40672 5922 40728
rect 5978 40672 6046 40728
rect 6102 40672 6170 40728
rect 6226 40672 6294 40728
rect 6350 40672 6418 40728
rect 6474 40672 6542 40728
rect 6598 40672 6666 40728
rect 6722 40672 6790 40728
rect 6846 40672 6914 40728
rect 6970 40672 7038 40728
rect 7094 40672 7104 40728
rect 5168 40604 7104 40672
rect 5168 40548 5178 40604
rect 5234 40548 5302 40604
rect 5358 40548 5426 40604
rect 5482 40548 5550 40604
rect 5606 40548 5674 40604
rect 5730 40548 5798 40604
rect 5854 40548 5922 40604
rect 5978 40548 6046 40604
rect 6102 40548 6170 40604
rect 6226 40548 6294 40604
rect 6350 40548 6418 40604
rect 6474 40548 6542 40604
rect 6598 40548 6666 40604
rect 6722 40548 6790 40604
rect 6846 40548 6914 40604
rect 6970 40548 7038 40604
rect 7094 40548 7104 40604
rect 5168 40480 7104 40548
rect 5168 40424 5178 40480
rect 5234 40424 5302 40480
rect 5358 40424 5426 40480
rect 5482 40424 5550 40480
rect 5606 40424 5674 40480
rect 5730 40424 5798 40480
rect 5854 40424 5922 40480
rect 5978 40424 6046 40480
rect 6102 40424 6170 40480
rect 6226 40424 6294 40480
rect 6350 40424 6418 40480
rect 6474 40424 6542 40480
rect 6598 40424 6666 40480
rect 6722 40424 6790 40480
rect 6846 40424 6914 40480
rect 6970 40424 7038 40480
rect 7094 40424 7104 40480
rect 5168 40356 7104 40424
rect 5168 40300 5178 40356
rect 5234 40300 5302 40356
rect 5358 40300 5426 40356
rect 5482 40300 5550 40356
rect 5606 40300 5674 40356
rect 5730 40300 5798 40356
rect 5854 40300 5922 40356
rect 5978 40300 6046 40356
rect 6102 40300 6170 40356
rect 6226 40300 6294 40356
rect 6350 40300 6418 40356
rect 6474 40300 6542 40356
rect 6598 40300 6666 40356
rect 6722 40300 6790 40356
rect 6846 40300 6914 40356
rect 6970 40300 7038 40356
rect 7094 40300 7104 40356
rect 5168 40232 7104 40300
rect 5168 40176 5178 40232
rect 5234 40176 5302 40232
rect 5358 40176 5426 40232
rect 5482 40176 5550 40232
rect 5606 40176 5674 40232
rect 5730 40176 5798 40232
rect 5854 40176 5922 40232
rect 5978 40176 6046 40232
rect 6102 40176 6170 40232
rect 6226 40176 6294 40232
rect 6350 40176 6418 40232
rect 6474 40176 6542 40232
rect 6598 40176 6666 40232
rect 6722 40176 6790 40232
rect 6846 40176 6914 40232
rect 6970 40176 7038 40232
rect 7094 40176 7104 40232
rect 5168 40108 7104 40176
rect 5168 40052 5178 40108
rect 5234 40052 5302 40108
rect 5358 40052 5426 40108
rect 5482 40052 5550 40108
rect 5606 40052 5674 40108
rect 5730 40052 5798 40108
rect 5854 40052 5922 40108
rect 5978 40052 6046 40108
rect 6102 40052 6170 40108
rect 6226 40052 6294 40108
rect 6350 40052 6418 40108
rect 6474 40052 6542 40108
rect 6598 40052 6666 40108
rect 6722 40052 6790 40108
rect 6846 40052 6914 40108
rect 6970 40052 7038 40108
rect 7094 40052 7104 40108
rect 5168 40042 7104 40052
rect 7874 41348 9810 41358
rect 7874 41292 7884 41348
rect 7940 41292 8008 41348
rect 8064 41292 8132 41348
rect 8188 41292 8256 41348
rect 8312 41292 8380 41348
rect 8436 41292 8504 41348
rect 8560 41292 8628 41348
rect 8684 41292 8752 41348
rect 8808 41292 8876 41348
rect 8932 41292 9000 41348
rect 9056 41292 9124 41348
rect 9180 41292 9248 41348
rect 9304 41292 9372 41348
rect 9428 41292 9496 41348
rect 9552 41292 9620 41348
rect 9676 41292 9744 41348
rect 9800 41292 9810 41348
rect 7874 41224 9810 41292
rect 7874 41168 7884 41224
rect 7940 41168 8008 41224
rect 8064 41168 8132 41224
rect 8188 41168 8256 41224
rect 8312 41168 8380 41224
rect 8436 41168 8504 41224
rect 8560 41168 8628 41224
rect 8684 41168 8752 41224
rect 8808 41168 8876 41224
rect 8932 41168 9000 41224
rect 9056 41168 9124 41224
rect 9180 41168 9248 41224
rect 9304 41168 9372 41224
rect 9428 41168 9496 41224
rect 9552 41168 9620 41224
rect 9676 41168 9744 41224
rect 9800 41168 9810 41224
rect 7874 41100 9810 41168
rect 7874 41044 7884 41100
rect 7940 41044 8008 41100
rect 8064 41044 8132 41100
rect 8188 41044 8256 41100
rect 8312 41044 8380 41100
rect 8436 41044 8504 41100
rect 8560 41044 8628 41100
rect 8684 41044 8752 41100
rect 8808 41044 8876 41100
rect 8932 41044 9000 41100
rect 9056 41044 9124 41100
rect 9180 41044 9248 41100
rect 9304 41044 9372 41100
rect 9428 41044 9496 41100
rect 9552 41044 9620 41100
rect 9676 41044 9744 41100
rect 9800 41044 9810 41100
rect 7874 40976 9810 41044
rect 7874 40920 7884 40976
rect 7940 40920 8008 40976
rect 8064 40920 8132 40976
rect 8188 40920 8256 40976
rect 8312 40920 8380 40976
rect 8436 40920 8504 40976
rect 8560 40920 8628 40976
rect 8684 40920 8752 40976
rect 8808 40920 8876 40976
rect 8932 40920 9000 40976
rect 9056 40920 9124 40976
rect 9180 40920 9248 40976
rect 9304 40920 9372 40976
rect 9428 40920 9496 40976
rect 9552 40920 9620 40976
rect 9676 40920 9744 40976
rect 9800 40920 9810 40976
rect 7874 40852 9810 40920
rect 7874 40796 7884 40852
rect 7940 40796 8008 40852
rect 8064 40796 8132 40852
rect 8188 40796 8256 40852
rect 8312 40796 8380 40852
rect 8436 40796 8504 40852
rect 8560 40796 8628 40852
rect 8684 40796 8752 40852
rect 8808 40796 8876 40852
rect 8932 40796 9000 40852
rect 9056 40796 9124 40852
rect 9180 40796 9248 40852
rect 9304 40796 9372 40852
rect 9428 40796 9496 40852
rect 9552 40796 9620 40852
rect 9676 40796 9744 40852
rect 9800 40796 9810 40852
rect 7874 40728 9810 40796
rect 7874 40672 7884 40728
rect 7940 40672 8008 40728
rect 8064 40672 8132 40728
rect 8188 40672 8256 40728
rect 8312 40672 8380 40728
rect 8436 40672 8504 40728
rect 8560 40672 8628 40728
rect 8684 40672 8752 40728
rect 8808 40672 8876 40728
rect 8932 40672 9000 40728
rect 9056 40672 9124 40728
rect 9180 40672 9248 40728
rect 9304 40672 9372 40728
rect 9428 40672 9496 40728
rect 9552 40672 9620 40728
rect 9676 40672 9744 40728
rect 9800 40672 9810 40728
rect 7874 40604 9810 40672
rect 7874 40548 7884 40604
rect 7940 40548 8008 40604
rect 8064 40548 8132 40604
rect 8188 40548 8256 40604
rect 8312 40548 8380 40604
rect 8436 40548 8504 40604
rect 8560 40548 8628 40604
rect 8684 40548 8752 40604
rect 8808 40548 8876 40604
rect 8932 40548 9000 40604
rect 9056 40548 9124 40604
rect 9180 40548 9248 40604
rect 9304 40548 9372 40604
rect 9428 40548 9496 40604
rect 9552 40548 9620 40604
rect 9676 40548 9744 40604
rect 9800 40548 9810 40604
rect 7874 40480 9810 40548
rect 7874 40424 7884 40480
rect 7940 40424 8008 40480
rect 8064 40424 8132 40480
rect 8188 40424 8256 40480
rect 8312 40424 8380 40480
rect 8436 40424 8504 40480
rect 8560 40424 8628 40480
rect 8684 40424 8752 40480
rect 8808 40424 8876 40480
rect 8932 40424 9000 40480
rect 9056 40424 9124 40480
rect 9180 40424 9248 40480
rect 9304 40424 9372 40480
rect 9428 40424 9496 40480
rect 9552 40424 9620 40480
rect 9676 40424 9744 40480
rect 9800 40424 9810 40480
rect 7874 40356 9810 40424
rect 7874 40300 7884 40356
rect 7940 40300 8008 40356
rect 8064 40300 8132 40356
rect 8188 40300 8256 40356
rect 8312 40300 8380 40356
rect 8436 40300 8504 40356
rect 8560 40300 8628 40356
rect 8684 40300 8752 40356
rect 8808 40300 8876 40356
rect 8932 40300 9000 40356
rect 9056 40300 9124 40356
rect 9180 40300 9248 40356
rect 9304 40300 9372 40356
rect 9428 40300 9496 40356
rect 9552 40300 9620 40356
rect 9676 40300 9744 40356
rect 9800 40300 9810 40356
rect 7874 40232 9810 40300
rect 7874 40176 7884 40232
rect 7940 40176 8008 40232
rect 8064 40176 8132 40232
rect 8188 40176 8256 40232
rect 8312 40176 8380 40232
rect 8436 40176 8504 40232
rect 8560 40176 8628 40232
rect 8684 40176 8752 40232
rect 8808 40176 8876 40232
rect 8932 40176 9000 40232
rect 9056 40176 9124 40232
rect 9180 40176 9248 40232
rect 9304 40176 9372 40232
rect 9428 40176 9496 40232
rect 9552 40176 9620 40232
rect 9676 40176 9744 40232
rect 9800 40176 9810 40232
rect 7874 40108 9810 40176
rect 7874 40052 7884 40108
rect 7940 40052 8008 40108
rect 8064 40052 8132 40108
rect 8188 40052 8256 40108
rect 8312 40052 8380 40108
rect 8436 40052 8504 40108
rect 8560 40052 8628 40108
rect 8684 40052 8752 40108
rect 8808 40052 8876 40108
rect 8932 40052 9000 40108
rect 9056 40052 9124 40108
rect 9180 40052 9248 40108
rect 9304 40052 9372 40108
rect 9428 40052 9496 40108
rect 9552 40052 9620 40108
rect 9676 40052 9744 40108
rect 9800 40052 9810 40108
rect 7874 40042 9810 40052
rect 10244 41348 12180 41358
rect 10244 41292 10254 41348
rect 10310 41292 10378 41348
rect 10434 41292 10502 41348
rect 10558 41292 10626 41348
rect 10682 41292 10750 41348
rect 10806 41292 10874 41348
rect 10930 41292 10998 41348
rect 11054 41292 11122 41348
rect 11178 41292 11246 41348
rect 11302 41292 11370 41348
rect 11426 41292 11494 41348
rect 11550 41292 11618 41348
rect 11674 41292 11742 41348
rect 11798 41292 11866 41348
rect 11922 41292 11990 41348
rect 12046 41292 12114 41348
rect 12170 41292 12180 41348
rect 10244 41224 12180 41292
rect 10244 41168 10254 41224
rect 10310 41168 10378 41224
rect 10434 41168 10502 41224
rect 10558 41168 10626 41224
rect 10682 41168 10750 41224
rect 10806 41168 10874 41224
rect 10930 41168 10998 41224
rect 11054 41168 11122 41224
rect 11178 41168 11246 41224
rect 11302 41168 11370 41224
rect 11426 41168 11494 41224
rect 11550 41168 11618 41224
rect 11674 41168 11742 41224
rect 11798 41168 11866 41224
rect 11922 41168 11990 41224
rect 12046 41168 12114 41224
rect 12170 41168 12180 41224
rect 10244 41100 12180 41168
rect 10244 41044 10254 41100
rect 10310 41044 10378 41100
rect 10434 41044 10502 41100
rect 10558 41044 10626 41100
rect 10682 41044 10750 41100
rect 10806 41044 10874 41100
rect 10930 41044 10998 41100
rect 11054 41044 11122 41100
rect 11178 41044 11246 41100
rect 11302 41044 11370 41100
rect 11426 41044 11494 41100
rect 11550 41044 11618 41100
rect 11674 41044 11742 41100
rect 11798 41044 11866 41100
rect 11922 41044 11990 41100
rect 12046 41044 12114 41100
rect 12170 41044 12180 41100
rect 10244 40976 12180 41044
rect 10244 40920 10254 40976
rect 10310 40920 10378 40976
rect 10434 40920 10502 40976
rect 10558 40920 10626 40976
rect 10682 40920 10750 40976
rect 10806 40920 10874 40976
rect 10930 40920 10998 40976
rect 11054 40920 11122 40976
rect 11178 40920 11246 40976
rect 11302 40920 11370 40976
rect 11426 40920 11494 40976
rect 11550 40920 11618 40976
rect 11674 40920 11742 40976
rect 11798 40920 11866 40976
rect 11922 40920 11990 40976
rect 12046 40920 12114 40976
rect 12170 40920 12180 40976
rect 10244 40852 12180 40920
rect 10244 40796 10254 40852
rect 10310 40796 10378 40852
rect 10434 40796 10502 40852
rect 10558 40796 10626 40852
rect 10682 40796 10750 40852
rect 10806 40796 10874 40852
rect 10930 40796 10998 40852
rect 11054 40796 11122 40852
rect 11178 40796 11246 40852
rect 11302 40796 11370 40852
rect 11426 40796 11494 40852
rect 11550 40796 11618 40852
rect 11674 40796 11742 40852
rect 11798 40796 11866 40852
rect 11922 40796 11990 40852
rect 12046 40796 12114 40852
rect 12170 40796 12180 40852
rect 10244 40728 12180 40796
rect 10244 40672 10254 40728
rect 10310 40672 10378 40728
rect 10434 40672 10502 40728
rect 10558 40672 10626 40728
rect 10682 40672 10750 40728
rect 10806 40672 10874 40728
rect 10930 40672 10998 40728
rect 11054 40672 11122 40728
rect 11178 40672 11246 40728
rect 11302 40672 11370 40728
rect 11426 40672 11494 40728
rect 11550 40672 11618 40728
rect 11674 40672 11742 40728
rect 11798 40672 11866 40728
rect 11922 40672 11990 40728
rect 12046 40672 12114 40728
rect 12170 40672 12180 40728
rect 10244 40604 12180 40672
rect 10244 40548 10254 40604
rect 10310 40548 10378 40604
rect 10434 40548 10502 40604
rect 10558 40548 10626 40604
rect 10682 40548 10750 40604
rect 10806 40548 10874 40604
rect 10930 40548 10998 40604
rect 11054 40548 11122 40604
rect 11178 40548 11246 40604
rect 11302 40548 11370 40604
rect 11426 40548 11494 40604
rect 11550 40548 11618 40604
rect 11674 40548 11742 40604
rect 11798 40548 11866 40604
rect 11922 40548 11990 40604
rect 12046 40548 12114 40604
rect 12170 40548 12180 40604
rect 10244 40480 12180 40548
rect 10244 40424 10254 40480
rect 10310 40424 10378 40480
rect 10434 40424 10502 40480
rect 10558 40424 10626 40480
rect 10682 40424 10750 40480
rect 10806 40424 10874 40480
rect 10930 40424 10998 40480
rect 11054 40424 11122 40480
rect 11178 40424 11246 40480
rect 11302 40424 11370 40480
rect 11426 40424 11494 40480
rect 11550 40424 11618 40480
rect 11674 40424 11742 40480
rect 11798 40424 11866 40480
rect 11922 40424 11990 40480
rect 12046 40424 12114 40480
rect 12170 40424 12180 40480
rect 10244 40356 12180 40424
rect 10244 40300 10254 40356
rect 10310 40300 10378 40356
rect 10434 40300 10502 40356
rect 10558 40300 10626 40356
rect 10682 40300 10750 40356
rect 10806 40300 10874 40356
rect 10930 40300 10998 40356
rect 11054 40300 11122 40356
rect 11178 40300 11246 40356
rect 11302 40300 11370 40356
rect 11426 40300 11494 40356
rect 11550 40300 11618 40356
rect 11674 40300 11742 40356
rect 11798 40300 11866 40356
rect 11922 40300 11990 40356
rect 12046 40300 12114 40356
rect 12170 40300 12180 40356
rect 10244 40232 12180 40300
rect 10244 40176 10254 40232
rect 10310 40176 10378 40232
rect 10434 40176 10502 40232
rect 10558 40176 10626 40232
rect 10682 40176 10750 40232
rect 10806 40176 10874 40232
rect 10930 40176 10998 40232
rect 11054 40176 11122 40232
rect 11178 40176 11246 40232
rect 11302 40176 11370 40232
rect 11426 40176 11494 40232
rect 11550 40176 11618 40232
rect 11674 40176 11742 40232
rect 11798 40176 11866 40232
rect 11922 40176 11990 40232
rect 12046 40176 12114 40232
rect 12170 40176 12180 40232
rect 10244 40108 12180 40176
rect 10244 40052 10254 40108
rect 10310 40052 10378 40108
rect 10434 40052 10502 40108
rect 10558 40052 10626 40108
rect 10682 40052 10750 40108
rect 10806 40052 10874 40108
rect 10930 40052 10998 40108
rect 11054 40052 11122 40108
rect 11178 40052 11246 40108
rect 11302 40052 11370 40108
rect 11426 40052 11494 40108
rect 11550 40052 11618 40108
rect 11674 40052 11742 40108
rect 11798 40052 11866 40108
rect 11922 40052 11990 40108
rect 12046 40052 12114 40108
rect 12170 40052 12180 40108
rect 10244 40042 12180 40052
rect 12861 41348 14673 41358
rect 12861 41292 12871 41348
rect 12927 41292 12995 41348
rect 13051 41292 13119 41348
rect 13175 41292 13243 41348
rect 13299 41292 13367 41348
rect 13423 41292 13491 41348
rect 13547 41292 13615 41348
rect 13671 41292 13739 41348
rect 13795 41292 13863 41348
rect 13919 41292 13987 41348
rect 14043 41292 14111 41348
rect 14167 41292 14235 41348
rect 14291 41292 14359 41348
rect 14415 41292 14483 41348
rect 14539 41292 14607 41348
rect 14663 41292 14673 41348
rect 12861 41224 14673 41292
rect 12861 41168 12871 41224
rect 12927 41168 12995 41224
rect 13051 41168 13119 41224
rect 13175 41168 13243 41224
rect 13299 41168 13367 41224
rect 13423 41168 13491 41224
rect 13547 41168 13615 41224
rect 13671 41168 13739 41224
rect 13795 41168 13863 41224
rect 13919 41168 13987 41224
rect 14043 41168 14111 41224
rect 14167 41168 14235 41224
rect 14291 41168 14359 41224
rect 14415 41168 14483 41224
rect 14539 41168 14607 41224
rect 14663 41168 14673 41224
rect 12861 41100 14673 41168
rect 12861 41044 12871 41100
rect 12927 41044 12995 41100
rect 13051 41044 13119 41100
rect 13175 41044 13243 41100
rect 13299 41044 13367 41100
rect 13423 41044 13491 41100
rect 13547 41044 13615 41100
rect 13671 41044 13739 41100
rect 13795 41044 13863 41100
rect 13919 41044 13987 41100
rect 14043 41044 14111 41100
rect 14167 41044 14235 41100
rect 14291 41044 14359 41100
rect 14415 41044 14483 41100
rect 14539 41044 14607 41100
rect 14663 41044 14673 41100
rect 12861 40976 14673 41044
rect 12861 40920 12871 40976
rect 12927 40920 12995 40976
rect 13051 40920 13119 40976
rect 13175 40920 13243 40976
rect 13299 40920 13367 40976
rect 13423 40920 13491 40976
rect 13547 40920 13615 40976
rect 13671 40920 13739 40976
rect 13795 40920 13863 40976
rect 13919 40920 13987 40976
rect 14043 40920 14111 40976
rect 14167 40920 14235 40976
rect 14291 40920 14359 40976
rect 14415 40920 14483 40976
rect 14539 40920 14607 40976
rect 14663 40920 14673 40976
rect 12861 40852 14673 40920
rect 12861 40796 12871 40852
rect 12927 40796 12995 40852
rect 13051 40796 13119 40852
rect 13175 40796 13243 40852
rect 13299 40796 13367 40852
rect 13423 40796 13491 40852
rect 13547 40796 13615 40852
rect 13671 40796 13739 40852
rect 13795 40796 13863 40852
rect 13919 40796 13987 40852
rect 14043 40796 14111 40852
rect 14167 40796 14235 40852
rect 14291 40796 14359 40852
rect 14415 40796 14483 40852
rect 14539 40796 14607 40852
rect 14663 40796 14673 40852
rect 12861 40728 14673 40796
rect 12861 40672 12871 40728
rect 12927 40672 12995 40728
rect 13051 40672 13119 40728
rect 13175 40672 13243 40728
rect 13299 40672 13367 40728
rect 13423 40672 13491 40728
rect 13547 40672 13615 40728
rect 13671 40672 13739 40728
rect 13795 40672 13863 40728
rect 13919 40672 13987 40728
rect 14043 40672 14111 40728
rect 14167 40672 14235 40728
rect 14291 40672 14359 40728
rect 14415 40672 14483 40728
rect 14539 40672 14607 40728
rect 14663 40672 14673 40728
rect 12861 40604 14673 40672
rect 12861 40548 12871 40604
rect 12927 40548 12995 40604
rect 13051 40548 13119 40604
rect 13175 40548 13243 40604
rect 13299 40548 13367 40604
rect 13423 40548 13491 40604
rect 13547 40548 13615 40604
rect 13671 40548 13739 40604
rect 13795 40548 13863 40604
rect 13919 40548 13987 40604
rect 14043 40548 14111 40604
rect 14167 40548 14235 40604
rect 14291 40548 14359 40604
rect 14415 40548 14483 40604
rect 14539 40548 14607 40604
rect 14663 40548 14673 40604
rect 12861 40480 14673 40548
rect 12861 40424 12871 40480
rect 12927 40424 12995 40480
rect 13051 40424 13119 40480
rect 13175 40424 13243 40480
rect 13299 40424 13367 40480
rect 13423 40424 13491 40480
rect 13547 40424 13615 40480
rect 13671 40424 13739 40480
rect 13795 40424 13863 40480
rect 13919 40424 13987 40480
rect 14043 40424 14111 40480
rect 14167 40424 14235 40480
rect 14291 40424 14359 40480
rect 14415 40424 14483 40480
rect 14539 40424 14607 40480
rect 14663 40424 14673 40480
rect 12861 40356 14673 40424
rect 12861 40300 12871 40356
rect 12927 40300 12995 40356
rect 13051 40300 13119 40356
rect 13175 40300 13243 40356
rect 13299 40300 13367 40356
rect 13423 40300 13491 40356
rect 13547 40300 13615 40356
rect 13671 40300 13739 40356
rect 13795 40300 13863 40356
rect 13919 40300 13987 40356
rect 14043 40300 14111 40356
rect 14167 40300 14235 40356
rect 14291 40300 14359 40356
rect 14415 40300 14483 40356
rect 14539 40300 14607 40356
rect 14663 40300 14673 40356
rect 12861 40232 14673 40300
rect 12861 40176 12871 40232
rect 12927 40176 12995 40232
rect 13051 40176 13119 40232
rect 13175 40176 13243 40232
rect 13299 40176 13367 40232
rect 13423 40176 13491 40232
rect 13547 40176 13615 40232
rect 13671 40176 13739 40232
rect 13795 40176 13863 40232
rect 13919 40176 13987 40232
rect 14043 40176 14111 40232
rect 14167 40176 14235 40232
rect 14291 40176 14359 40232
rect 14415 40176 14483 40232
rect 14539 40176 14607 40232
rect 14663 40176 14673 40232
rect 12861 40108 14673 40176
rect 12861 40052 12871 40108
rect 12927 40052 12995 40108
rect 13051 40052 13119 40108
rect 13175 40052 13243 40108
rect 13299 40052 13367 40108
rect 13423 40052 13491 40108
rect 13547 40052 13615 40108
rect 13671 40052 13739 40108
rect 13795 40052 13863 40108
rect 13919 40052 13987 40108
rect 14043 40052 14111 40108
rect 14167 40052 14235 40108
rect 14291 40052 14359 40108
rect 14415 40052 14483 40108
rect 14539 40052 14607 40108
rect 14663 40052 14673 40108
rect 12861 40042 14673 40052
rect 2798 39748 4734 39758
rect 2798 39692 2808 39748
rect 2864 39692 2932 39748
rect 2988 39692 3056 39748
rect 3112 39692 3180 39748
rect 3236 39692 3304 39748
rect 3360 39692 3428 39748
rect 3484 39692 3552 39748
rect 3608 39692 3676 39748
rect 3732 39692 3800 39748
rect 3856 39692 3924 39748
rect 3980 39692 4048 39748
rect 4104 39692 4172 39748
rect 4228 39692 4296 39748
rect 4352 39692 4420 39748
rect 4476 39692 4544 39748
rect 4600 39692 4668 39748
rect 4724 39692 4734 39748
rect 2798 39624 4734 39692
rect 2798 39568 2808 39624
rect 2864 39568 2932 39624
rect 2988 39568 3056 39624
rect 3112 39568 3180 39624
rect 3236 39568 3304 39624
rect 3360 39568 3428 39624
rect 3484 39568 3552 39624
rect 3608 39568 3676 39624
rect 3732 39568 3800 39624
rect 3856 39568 3924 39624
rect 3980 39568 4048 39624
rect 4104 39568 4172 39624
rect 4228 39568 4296 39624
rect 4352 39568 4420 39624
rect 4476 39568 4544 39624
rect 4600 39568 4668 39624
rect 4724 39568 4734 39624
rect 2798 39500 4734 39568
rect 2798 39444 2808 39500
rect 2864 39444 2932 39500
rect 2988 39444 3056 39500
rect 3112 39444 3180 39500
rect 3236 39444 3304 39500
rect 3360 39444 3428 39500
rect 3484 39444 3552 39500
rect 3608 39444 3676 39500
rect 3732 39444 3800 39500
rect 3856 39444 3924 39500
rect 3980 39444 4048 39500
rect 4104 39444 4172 39500
rect 4228 39444 4296 39500
rect 4352 39444 4420 39500
rect 4476 39444 4544 39500
rect 4600 39444 4668 39500
rect 4724 39444 4734 39500
rect 2798 39376 4734 39444
rect 2798 39320 2808 39376
rect 2864 39320 2932 39376
rect 2988 39320 3056 39376
rect 3112 39320 3180 39376
rect 3236 39320 3304 39376
rect 3360 39320 3428 39376
rect 3484 39320 3552 39376
rect 3608 39320 3676 39376
rect 3732 39320 3800 39376
rect 3856 39320 3924 39376
rect 3980 39320 4048 39376
rect 4104 39320 4172 39376
rect 4228 39320 4296 39376
rect 4352 39320 4420 39376
rect 4476 39320 4544 39376
rect 4600 39320 4668 39376
rect 4724 39320 4734 39376
rect 2798 39252 4734 39320
rect 2798 39196 2808 39252
rect 2864 39196 2932 39252
rect 2988 39196 3056 39252
rect 3112 39196 3180 39252
rect 3236 39196 3304 39252
rect 3360 39196 3428 39252
rect 3484 39196 3552 39252
rect 3608 39196 3676 39252
rect 3732 39196 3800 39252
rect 3856 39196 3924 39252
rect 3980 39196 4048 39252
rect 4104 39196 4172 39252
rect 4228 39196 4296 39252
rect 4352 39196 4420 39252
rect 4476 39196 4544 39252
rect 4600 39196 4668 39252
rect 4724 39196 4734 39252
rect 2798 39128 4734 39196
rect 2798 39072 2808 39128
rect 2864 39072 2932 39128
rect 2988 39072 3056 39128
rect 3112 39072 3180 39128
rect 3236 39072 3304 39128
rect 3360 39072 3428 39128
rect 3484 39072 3552 39128
rect 3608 39072 3676 39128
rect 3732 39072 3800 39128
rect 3856 39072 3924 39128
rect 3980 39072 4048 39128
rect 4104 39072 4172 39128
rect 4228 39072 4296 39128
rect 4352 39072 4420 39128
rect 4476 39072 4544 39128
rect 4600 39072 4668 39128
rect 4724 39072 4734 39128
rect 2798 39004 4734 39072
rect 2798 38948 2808 39004
rect 2864 38948 2932 39004
rect 2988 38948 3056 39004
rect 3112 38948 3180 39004
rect 3236 38948 3304 39004
rect 3360 38948 3428 39004
rect 3484 38948 3552 39004
rect 3608 38948 3676 39004
rect 3732 38948 3800 39004
rect 3856 38948 3924 39004
rect 3980 38948 4048 39004
rect 4104 38948 4172 39004
rect 4228 38948 4296 39004
rect 4352 38948 4420 39004
rect 4476 38948 4544 39004
rect 4600 38948 4668 39004
rect 4724 38948 4734 39004
rect 2798 38880 4734 38948
rect 2798 38824 2808 38880
rect 2864 38824 2932 38880
rect 2988 38824 3056 38880
rect 3112 38824 3180 38880
rect 3236 38824 3304 38880
rect 3360 38824 3428 38880
rect 3484 38824 3552 38880
rect 3608 38824 3676 38880
rect 3732 38824 3800 38880
rect 3856 38824 3924 38880
rect 3980 38824 4048 38880
rect 4104 38824 4172 38880
rect 4228 38824 4296 38880
rect 4352 38824 4420 38880
rect 4476 38824 4544 38880
rect 4600 38824 4668 38880
rect 4724 38824 4734 38880
rect 2798 38756 4734 38824
rect 2798 38700 2808 38756
rect 2864 38700 2932 38756
rect 2988 38700 3056 38756
rect 3112 38700 3180 38756
rect 3236 38700 3304 38756
rect 3360 38700 3428 38756
rect 3484 38700 3552 38756
rect 3608 38700 3676 38756
rect 3732 38700 3800 38756
rect 3856 38700 3924 38756
rect 3980 38700 4048 38756
rect 4104 38700 4172 38756
rect 4228 38700 4296 38756
rect 4352 38700 4420 38756
rect 4476 38700 4544 38756
rect 4600 38700 4668 38756
rect 4724 38700 4734 38756
rect 2798 38632 4734 38700
rect 2798 38576 2808 38632
rect 2864 38576 2932 38632
rect 2988 38576 3056 38632
rect 3112 38576 3180 38632
rect 3236 38576 3304 38632
rect 3360 38576 3428 38632
rect 3484 38576 3552 38632
rect 3608 38576 3676 38632
rect 3732 38576 3800 38632
rect 3856 38576 3924 38632
rect 3980 38576 4048 38632
rect 4104 38576 4172 38632
rect 4228 38576 4296 38632
rect 4352 38576 4420 38632
rect 4476 38576 4544 38632
rect 4600 38576 4668 38632
rect 4724 38576 4734 38632
rect 2798 38508 4734 38576
rect 2798 38452 2808 38508
rect 2864 38452 2932 38508
rect 2988 38452 3056 38508
rect 3112 38452 3180 38508
rect 3236 38452 3304 38508
rect 3360 38452 3428 38508
rect 3484 38452 3552 38508
rect 3608 38452 3676 38508
rect 3732 38452 3800 38508
rect 3856 38452 3924 38508
rect 3980 38452 4048 38508
rect 4104 38452 4172 38508
rect 4228 38452 4296 38508
rect 4352 38452 4420 38508
rect 4476 38452 4544 38508
rect 4600 38452 4668 38508
rect 4724 38452 4734 38508
rect 2798 38442 4734 38452
rect 5168 39748 7104 39758
rect 5168 39692 5178 39748
rect 5234 39692 5302 39748
rect 5358 39692 5426 39748
rect 5482 39692 5550 39748
rect 5606 39692 5674 39748
rect 5730 39692 5798 39748
rect 5854 39692 5922 39748
rect 5978 39692 6046 39748
rect 6102 39692 6170 39748
rect 6226 39692 6294 39748
rect 6350 39692 6418 39748
rect 6474 39692 6542 39748
rect 6598 39692 6666 39748
rect 6722 39692 6790 39748
rect 6846 39692 6914 39748
rect 6970 39692 7038 39748
rect 7094 39692 7104 39748
rect 5168 39624 7104 39692
rect 5168 39568 5178 39624
rect 5234 39568 5302 39624
rect 5358 39568 5426 39624
rect 5482 39568 5550 39624
rect 5606 39568 5674 39624
rect 5730 39568 5798 39624
rect 5854 39568 5922 39624
rect 5978 39568 6046 39624
rect 6102 39568 6170 39624
rect 6226 39568 6294 39624
rect 6350 39568 6418 39624
rect 6474 39568 6542 39624
rect 6598 39568 6666 39624
rect 6722 39568 6790 39624
rect 6846 39568 6914 39624
rect 6970 39568 7038 39624
rect 7094 39568 7104 39624
rect 5168 39500 7104 39568
rect 5168 39444 5178 39500
rect 5234 39444 5302 39500
rect 5358 39444 5426 39500
rect 5482 39444 5550 39500
rect 5606 39444 5674 39500
rect 5730 39444 5798 39500
rect 5854 39444 5922 39500
rect 5978 39444 6046 39500
rect 6102 39444 6170 39500
rect 6226 39444 6294 39500
rect 6350 39444 6418 39500
rect 6474 39444 6542 39500
rect 6598 39444 6666 39500
rect 6722 39444 6790 39500
rect 6846 39444 6914 39500
rect 6970 39444 7038 39500
rect 7094 39444 7104 39500
rect 5168 39376 7104 39444
rect 5168 39320 5178 39376
rect 5234 39320 5302 39376
rect 5358 39320 5426 39376
rect 5482 39320 5550 39376
rect 5606 39320 5674 39376
rect 5730 39320 5798 39376
rect 5854 39320 5922 39376
rect 5978 39320 6046 39376
rect 6102 39320 6170 39376
rect 6226 39320 6294 39376
rect 6350 39320 6418 39376
rect 6474 39320 6542 39376
rect 6598 39320 6666 39376
rect 6722 39320 6790 39376
rect 6846 39320 6914 39376
rect 6970 39320 7038 39376
rect 7094 39320 7104 39376
rect 5168 39252 7104 39320
rect 5168 39196 5178 39252
rect 5234 39196 5302 39252
rect 5358 39196 5426 39252
rect 5482 39196 5550 39252
rect 5606 39196 5674 39252
rect 5730 39196 5798 39252
rect 5854 39196 5922 39252
rect 5978 39196 6046 39252
rect 6102 39196 6170 39252
rect 6226 39196 6294 39252
rect 6350 39196 6418 39252
rect 6474 39196 6542 39252
rect 6598 39196 6666 39252
rect 6722 39196 6790 39252
rect 6846 39196 6914 39252
rect 6970 39196 7038 39252
rect 7094 39196 7104 39252
rect 5168 39128 7104 39196
rect 5168 39072 5178 39128
rect 5234 39072 5302 39128
rect 5358 39072 5426 39128
rect 5482 39072 5550 39128
rect 5606 39072 5674 39128
rect 5730 39072 5798 39128
rect 5854 39072 5922 39128
rect 5978 39072 6046 39128
rect 6102 39072 6170 39128
rect 6226 39072 6294 39128
rect 6350 39072 6418 39128
rect 6474 39072 6542 39128
rect 6598 39072 6666 39128
rect 6722 39072 6790 39128
rect 6846 39072 6914 39128
rect 6970 39072 7038 39128
rect 7094 39072 7104 39128
rect 5168 39004 7104 39072
rect 5168 38948 5178 39004
rect 5234 38948 5302 39004
rect 5358 38948 5426 39004
rect 5482 38948 5550 39004
rect 5606 38948 5674 39004
rect 5730 38948 5798 39004
rect 5854 38948 5922 39004
rect 5978 38948 6046 39004
rect 6102 38948 6170 39004
rect 6226 38948 6294 39004
rect 6350 38948 6418 39004
rect 6474 38948 6542 39004
rect 6598 38948 6666 39004
rect 6722 38948 6790 39004
rect 6846 38948 6914 39004
rect 6970 38948 7038 39004
rect 7094 38948 7104 39004
rect 5168 38880 7104 38948
rect 5168 38824 5178 38880
rect 5234 38824 5302 38880
rect 5358 38824 5426 38880
rect 5482 38824 5550 38880
rect 5606 38824 5674 38880
rect 5730 38824 5798 38880
rect 5854 38824 5922 38880
rect 5978 38824 6046 38880
rect 6102 38824 6170 38880
rect 6226 38824 6294 38880
rect 6350 38824 6418 38880
rect 6474 38824 6542 38880
rect 6598 38824 6666 38880
rect 6722 38824 6790 38880
rect 6846 38824 6914 38880
rect 6970 38824 7038 38880
rect 7094 38824 7104 38880
rect 5168 38756 7104 38824
rect 5168 38700 5178 38756
rect 5234 38700 5302 38756
rect 5358 38700 5426 38756
rect 5482 38700 5550 38756
rect 5606 38700 5674 38756
rect 5730 38700 5798 38756
rect 5854 38700 5922 38756
rect 5978 38700 6046 38756
rect 6102 38700 6170 38756
rect 6226 38700 6294 38756
rect 6350 38700 6418 38756
rect 6474 38700 6542 38756
rect 6598 38700 6666 38756
rect 6722 38700 6790 38756
rect 6846 38700 6914 38756
rect 6970 38700 7038 38756
rect 7094 38700 7104 38756
rect 5168 38632 7104 38700
rect 5168 38576 5178 38632
rect 5234 38576 5302 38632
rect 5358 38576 5426 38632
rect 5482 38576 5550 38632
rect 5606 38576 5674 38632
rect 5730 38576 5798 38632
rect 5854 38576 5922 38632
rect 5978 38576 6046 38632
rect 6102 38576 6170 38632
rect 6226 38576 6294 38632
rect 6350 38576 6418 38632
rect 6474 38576 6542 38632
rect 6598 38576 6666 38632
rect 6722 38576 6790 38632
rect 6846 38576 6914 38632
rect 6970 38576 7038 38632
rect 7094 38576 7104 38632
rect 5168 38508 7104 38576
rect 5168 38452 5178 38508
rect 5234 38452 5302 38508
rect 5358 38452 5426 38508
rect 5482 38452 5550 38508
rect 5606 38452 5674 38508
rect 5730 38452 5798 38508
rect 5854 38452 5922 38508
rect 5978 38452 6046 38508
rect 6102 38452 6170 38508
rect 6226 38452 6294 38508
rect 6350 38452 6418 38508
rect 6474 38452 6542 38508
rect 6598 38452 6666 38508
rect 6722 38452 6790 38508
rect 6846 38452 6914 38508
rect 6970 38452 7038 38508
rect 7094 38452 7104 38508
rect 5168 38442 7104 38452
rect 7874 39748 9810 39758
rect 7874 39692 7884 39748
rect 7940 39692 8008 39748
rect 8064 39692 8132 39748
rect 8188 39692 8256 39748
rect 8312 39692 8380 39748
rect 8436 39692 8504 39748
rect 8560 39692 8628 39748
rect 8684 39692 8752 39748
rect 8808 39692 8876 39748
rect 8932 39692 9000 39748
rect 9056 39692 9124 39748
rect 9180 39692 9248 39748
rect 9304 39692 9372 39748
rect 9428 39692 9496 39748
rect 9552 39692 9620 39748
rect 9676 39692 9744 39748
rect 9800 39692 9810 39748
rect 7874 39624 9810 39692
rect 7874 39568 7884 39624
rect 7940 39568 8008 39624
rect 8064 39568 8132 39624
rect 8188 39568 8256 39624
rect 8312 39568 8380 39624
rect 8436 39568 8504 39624
rect 8560 39568 8628 39624
rect 8684 39568 8752 39624
rect 8808 39568 8876 39624
rect 8932 39568 9000 39624
rect 9056 39568 9124 39624
rect 9180 39568 9248 39624
rect 9304 39568 9372 39624
rect 9428 39568 9496 39624
rect 9552 39568 9620 39624
rect 9676 39568 9744 39624
rect 9800 39568 9810 39624
rect 7874 39500 9810 39568
rect 7874 39444 7884 39500
rect 7940 39444 8008 39500
rect 8064 39444 8132 39500
rect 8188 39444 8256 39500
rect 8312 39444 8380 39500
rect 8436 39444 8504 39500
rect 8560 39444 8628 39500
rect 8684 39444 8752 39500
rect 8808 39444 8876 39500
rect 8932 39444 9000 39500
rect 9056 39444 9124 39500
rect 9180 39444 9248 39500
rect 9304 39444 9372 39500
rect 9428 39444 9496 39500
rect 9552 39444 9620 39500
rect 9676 39444 9744 39500
rect 9800 39444 9810 39500
rect 7874 39376 9810 39444
rect 7874 39320 7884 39376
rect 7940 39320 8008 39376
rect 8064 39320 8132 39376
rect 8188 39320 8256 39376
rect 8312 39320 8380 39376
rect 8436 39320 8504 39376
rect 8560 39320 8628 39376
rect 8684 39320 8752 39376
rect 8808 39320 8876 39376
rect 8932 39320 9000 39376
rect 9056 39320 9124 39376
rect 9180 39320 9248 39376
rect 9304 39320 9372 39376
rect 9428 39320 9496 39376
rect 9552 39320 9620 39376
rect 9676 39320 9744 39376
rect 9800 39320 9810 39376
rect 7874 39252 9810 39320
rect 7874 39196 7884 39252
rect 7940 39196 8008 39252
rect 8064 39196 8132 39252
rect 8188 39196 8256 39252
rect 8312 39196 8380 39252
rect 8436 39196 8504 39252
rect 8560 39196 8628 39252
rect 8684 39196 8752 39252
rect 8808 39196 8876 39252
rect 8932 39196 9000 39252
rect 9056 39196 9124 39252
rect 9180 39196 9248 39252
rect 9304 39196 9372 39252
rect 9428 39196 9496 39252
rect 9552 39196 9620 39252
rect 9676 39196 9744 39252
rect 9800 39196 9810 39252
rect 7874 39128 9810 39196
rect 7874 39072 7884 39128
rect 7940 39072 8008 39128
rect 8064 39072 8132 39128
rect 8188 39072 8256 39128
rect 8312 39072 8380 39128
rect 8436 39072 8504 39128
rect 8560 39072 8628 39128
rect 8684 39072 8752 39128
rect 8808 39072 8876 39128
rect 8932 39072 9000 39128
rect 9056 39072 9124 39128
rect 9180 39072 9248 39128
rect 9304 39072 9372 39128
rect 9428 39072 9496 39128
rect 9552 39072 9620 39128
rect 9676 39072 9744 39128
rect 9800 39072 9810 39128
rect 7874 39004 9810 39072
rect 7874 38948 7884 39004
rect 7940 38948 8008 39004
rect 8064 38948 8132 39004
rect 8188 38948 8256 39004
rect 8312 38948 8380 39004
rect 8436 38948 8504 39004
rect 8560 38948 8628 39004
rect 8684 38948 8752 39004
rect 8808 38948 8876 39004
rect 8932 38948 9000 39004
rect 9056 38948 9124 39004
rect 9180 38948 9248 39004
rect 9304 38948 9372 39004
rect 9428 38948 9496 39004
rect 9552 38948 9620 39004
rect 9676 38948 9744 39004
rect 9800 38948 9810 39004
rect 7874 38880 9810 38948
rect 7874 38824 7884 38880
rect 7940 38824 8008 38880
rect 8064 38824 8132 38880
rect 8188 38824 8256 38880
rect 8312 38824 8380 38880
rect 8436 38824 8504 38880
rect 8560 38824 8628 38880
rect 8684 38824 8752 38880
rect 8808 38824 8876 38880
rect 8932 38824 9000 38880
rect 9056 38824 9124 38880
rect 9180 38824 9248 38880
rect 9304 38824 9372 38880
rect 9428 38824 9496 38880
rect 9552 38824 9620 38880
rect 9676 38824 9744 38880
rect 9800 38824 9810 38880
rect 7874 38756 9810 38824
rect 7874 38700 7884 38756
rect 7940 38700 8008 38756
rect 8064 38700 8132 38756
rect 8188 38700 8256 38756
rect 8312 38700 8380 38756
rect 8436 38700 8504 38756
rect 8560 38700 8628 38756
rect 8684 38700 8752 38756
rect 8808 38700 8876 38756
rect 8932 38700 9000 38756
rect 9056 38700 9124 38756
rect 9180 38700 9248 38756
rect 9304 38700 9372 38756
rect 9428 38700 9496 38756
rect 9552 38700 9620 38756
rect 9676 38700 9744 38756
rect 9800 38700 9810 38756
rect 7874 38632 9810 38700
rect 7874 38576 7884 38632
rect 7940 38576 8008 38632
rect 8064 38576 8132 38632
rect 8188 38576 8256 38632
rect 8312 38576 8380 38632
rect 8436 38576 8504 38632
rect 8560 38576 8628 38632
rect 8684 38576 8752 38632
rect 8808 38576 8876 38632
rect 8932 38576 9000 38632
rect 9056 38576 9124 38632
rect 9180 38576 9248 38632
rect 9304 38576 9372 38632
rect 9428 38576 9496 38632
rect 9552 38576 9620 38632
rect 9676 38576 9744 38632
rect 9800 38576 9810 38632
rect 7874 38508 9810 38576
rect 7874 38452 7884 38508
rect 7940 38452 8008 38508
rect 8064 38452 8132 38508
rect 8188 38452 8256 38508
rect 8312 38452 8380 38508
rect 8436 38452 8504 38508
rect 8560 38452 8628 38508
rect 8684 38452 8752 38508
rect 8808 38452 8876 38508
rect 8932 38452 9000 38508
rect 9056 38452 9124 38508
rect 9180 38452 9248 38508
rect 9304 38452 9372 38508
rect 9428 38452 9496 38508
rect 9552 38452 9620 38508
rect 9676 38452 9744 38508
rect 9800 38452 9810 38508
rect 7874 38442 9810 38452
rect 10244 39748 12180 39758
rect 10244 39692 10254 39748
rect 10310 39692 10378 39748
rect 10434 39692 10502 39748
rect 10558 39692 10626 39748
rect 10682 39692 10750 39748
rect 10806 39692 10874 39748
rect 10930 39692 10998 39748
rect 11054 39692 11122 39748
rect 11178 39692 11246 39748
rect 11302 39692 11370 39748
rect 11426 39692 11494 39748
rect 11550 39692 11618 39748
rect 11674 39692 11742 39748
rect 11798 39692 11866 39748
rect 11922 39692 11990 39748
rect 12046 39692 12114 39748
rect 12170 39692 12180 39748
rect 10244 39624 12180 39692
rect 10244 39568 10254 39624
rect 10310 39568 10378 39624
rect 10434 39568 10502 39624
rect 10558 39568 10626 39624
rect 10682 39568 10750 39624
rect 10806 39568 10874 39624
rect 10930 39568 10998 39624
rect 11054 39568 11122 39624
rect 11178 39568 11246 39624
rect 11302 39568 11370 39624
rect 11426 39568 11494 39624
rect 11550 39568 11618 39624
rect 11674 39568 11742 39624
rect 11798 39568 11866 39624
rect 11922 39568 11990 39624
rect 12046 39568 12114 39624
rect 12170 39568 12180 39624
rect 10244 39500 12180 39568
rect 10244 39444 10254 39500
rect 10310 39444 10378 39500
rect 10434 39444 10502 39500
rect 10558 39444 10626 39500
rect 10682 39444 10750 39500
rect 10806 39444 10874 39500
rect 10930 39444 10998 39500
rect 11054 39444 11122 39500
rect 11178 39444 11246 39500
rect 11302 39444 11370 39500
rect 11426 39444 11494 39500
rect 11550 39444 11618 39500
rect 11674 39444 11742 39500
rect 11798 39444 11866 39500
rect 11922 39444 11990 39500
rect 12046 39444 12114 39500
rect 12170 39444 12180 39500
rect 10244 39376 12180 39444
rect 10244 39320 10254 39376
rect 10310 39320 10378 39376
rect 10434 39320 10502 39376
rect 10558 39320 10626 39376
rect 10682 39320 10750 39376
rect 10806 39320 10874 39376
rect 10930 39320 10998 39376
rect 11054 39320 11122 39376
rect 11178 39320 11246 39376
rect 11302 39320 11370 39376
rect 11426 39320 11494 39376
rect 11550 39320 11618 39376
rect 11674 39320 11742 39376
rect 11798 39320 11866 39376
rect 11922 39320 11990 39376
rect 12046 39320 12114 39376
rect 12170 39320 12180 39376
rect 10244 39252 12180 39320
rect 10244 39196 10254 39252
rect 10310 39196 10378 39252
rect 10434 39196 10502 39252
rect 10558 39196 10626 39252
rect 10682 39196 10750 39252
rect 10806 39196 10874 39252
rect 10930 39196 10998 39252
rect 11054 39196 11122 39252
rect 11178 39196 11246 39252
rect 11302 39196 11370 39252
rect 11426 39196 11494 39252
rect 11550 39196 11618 39252
rect 11674 39196 11742 39252
rect 11798 39196 11866 39252
rect 11922 39196 11990 39252
rect 12046 39196 12114 39252
rect 12170 39196 12180 39252
rect 10244 39128 12180 39196
rect 10244 39072 10254 39128
rect 10310 39072 10378 39128
rect 10434 39072 10502 39128
rect 10558 39072 10626 39128
rect 10682 39072 10750 39128
rect 10806 39072 10874 39128
rect 10930 39072 10998 39128
rect 11054 39072 11122 39128
rect 11178 39072 11246 39128
rect 11302 39072 11370 39128
rect 11426 39072 11494 39128
rect 11550 39072 11618 39128
rect 11674 39072 11742 39128
rect 11798 39072 11866 39128
rect 11922 39072 11990 39128
rect 12046 39072 12114 39128
rect 12170 39072 12180 39128
rect 10244 39004 12180 39072
rect 10244 38948 10254 39004
rect 10310 38948 10378 39004
rect 10434 38948 10502 39004
rect 10558 38948 10626 39004
rect 10682 38948 10750 39004
rect 10806 38948 10874 39004
rect 10930 38948 10998 39004
rect 11054 38948 11122 39004
rect 11178 38948 11246 39004
rect 11302 38948 11370 39004
rect 11426 38948 11494 39004
rect 11550 38948 11618 39004
rect 11674 38948 11742 39004
rect 11798 38948 11866 39004
rect 11922 38948 11990 39004
rect 12046 38948 12114 39004
rect 12170 38948 12180 39004
rect 10244 38880 12180 38948
rect 10244 38824 10254 38880
rect 10310 38824 10378 38880
rect 10434 38824 10502 38880
rect 10558 38824 10626 38880
rect 10682 38824 10750 38880
rect 10806 38824 10874 38880
rect 10930 38824 10998 38880
rect 11054 38824 11122 38880
rect 11178 38824 11246 38880
rect 11302 38824 11370 38880
rect 11426 38824 11494 38880
rect 11550 38824 11618 38880
rect 11674 38824 11742 38880
rect 11798 38824 11866 38880
rect 11922 38824 11990 38880
rect 12046 38824 12114 38880
rect 12170 38824 12180 38880
rect 10244 38756 12180 38824
rect 10244 38700 10254 38756
rect 10310 38700 10378 38756
rect 10434 38700 10502 38756
rect 10558 38700 10626 38756
rect 10682 38700 10750 38756
rect 10806 38700 10874 38756
rect 10930 38700 10998 38756
rect 11054 38700 11122 38756
rect 11178 38700 11246 38756
rect 11302 38700 11370 38756
rect 11426 38700 11494 38756
rect 11550 38700 11618 38756
rect 11674 38700 11742 38756
rect 11798 38700 11866 38756
rect 11922 38700 11990 38756
rect 12046 38700 12114 38756
rect 12170 38700 12180 38756
rect 10244 38632 12180 38700
rect 10244 38576 10254 38632
rect 10310 38576 10378 38632
rect 10434 38576 10502 38632
rect 10558 38576 10626 38632
rect 10682 38576 10750 38632
rect 10806 38576 10874 38632
rect 10930 38576 10998 38632
rect 11054 38576 11122 38632
rect 11178 38576 11246 38632
rect 11302 38576 11370 38632
rect 11426 38576 11494 38632
rect 11550 38576 11618 38632
rect 11674 38576 11742 38632
rect 11798 38576 11866 38632
rect 11922 38576 11990 38632
rect 12046 38576 12114 38632
rect 12170 38576 12180 38632
rect 10244 38508 12180 38576
rect 10244 38452 10254 38508
rect 10310 38452 10378 38508
rect 10434 38452 10502 38508
rect 10558 38452 10626 38508
rect 10682 38452 10750 38508
rect 10806 38452 10874 38508
rect 10930 38452 10998 38508
rect 11054 38452 11122 38508
rect 11178 38452 11246 38508
rect 11302 38452 11370 38508
rect 11426 38452 11494 38508
rect 11550 38452 11618 38508
rect 11674 38452 11742 38508
rect 11798 38452 11866 38508
rect 11922 38452 11990 38508
rect 12046 38452 12114 38508
rect 12170 38452 12180 38508
rect 10244 38442 12180 38452
rect 12861 39748 14673 39758
rect 12861 39692 12871 39748
rect 12927 39692 12995 39748
rect 13051 39692 13119 39748
rect 13175 39692 13243 39748
rect 13299 39692 13367 39748
rect 13423 39692 13491 39748
rect 13547 39692 13615 39748
rect 13671 39692 13739 39748
rect 13795 39692 13863 39748
rect 13919 39692 13987 39748
rect 14043 39692 14111 39748
rect 14167 39692 14235 39748
rect 14291 39692 14359 39748
rect 14415 39692 14483 39748
rect 14539 39692 14607 39748
rect 14663 39692 14673 39748
rect 12861 39624 14673 39692
rect 12861 39568 12871 39624
rect 12927 39568 12995 39624
rect 13051 39568 13119 39624
rect 13175 39568 13243 39624
rect 13299 39568 13367 39624
rect 13423 39568 13491 39624
rect 13547 39568 13615 39624
rect 13671 39568 13739 39624
rect 13795 39568 13863 39624
rect 13919 39568 13987 39624
rect 14043 39568 14111 39624
rect 14167 39568 14235 39624
rect 14291 39568 14359 39624
rect 14415 39568 14483 39624
rect 14539 39568 14607 39624
rect 14663 39568 14673 39624
rect 12861 39500 14673 39568
rect 12861 39444 12871 39500
rect 12927 39444 12995 39500
rect 13051 39444 13119 39500
rect 13175 39444 13243 39500
rect 13299 39444 13367 39500
rect 13423 39444 13491 39500
rect 13547 39444 13615 39500
rect 13671 39444 13739 39500
rect 13795 39444 13863 39500
rect 13919 39444 13987 39500
rect 14043 39444 14111 39500
rect 14167 39444 14235 39500
rect 14291 39444 14359 39500
rect 14415 39444 14483 39500
rect 14539 39444 14607 39500
rect 14663 39444 14673 39500
rect 12861 39376 14673 39444
rect 12861 39320 12871 39376
rect 12927 39320 12995 39376
rect 13051 39320 13119 39376
rect 13175 39320 13243 39376
rect 13299 39320 13367 39376
rect 13423 39320 13491 39376
rect 13547 39320 13615 39376
rect 13671 39320 13739 39376
rect 13795 39320 13863 39376
rect 13919 39320 13987 39376
rect 14043 39320 14111 39376
rect 14167 39320 14235 39376
rect 14291 39320 14359 39376
rect 14415 39320 14483 39376
rect 14539 39320 14607 39376
rect 14663 39320 14673 39376
rect 12861 39252 14673 39320
rect 12861 39196 12871 39252
rect 12927 39196 12995 39252
rect 13051 39196 13119 39252
rect 13175 39196 13243 39252
rect 13299 39196 13367 39252
rect 13423 39196 13491 39252
rect 13547 39196 13615 39252
rect 13671 39196 13739 39252
rect 13795 39196 13863 39252
rect 13919 39196 13987 39252
rect 14043 39196 14111 39252
rect 14167 39196 14235 39252
rect 14291 39196 14359 39252
rect 14415 39196 14483 39252
rect 14539 39196 14607 39252
rect 14663 39196 14673 39252
rect 12861 39128 14673 39196
rect 12861 39072 12871 39128
rect 12927 39072 12995 39128
rect 13051 39072 13119 39128
rect 13175 39072 13243 39128
rect 13299 39072 13367 39128
rect 13423 39072 13491 39128
rect 13547 39072 13615 39128
rect 13671 39072 13739 39128
rect 13795 39072 13863 39128
rect 13919 39072 13987 39128
rect 14043 39072 14111 39128
rect 14167 39072 14235 39128
rect 14291 39072 14359 39128
rect 14415 39072 14483 39128
rect 14539 39072 14607 39128
rect 14663 39072 14673 39128
rect 12861 39004 14673 39072
rect 12861 38948 12871 39004
rect 12927 38948 12995 39004
rect 13051 38948 13119 39004
rect 13175 38948 13243 39004
rect 13299 38948 13367 39004
rect 13423 38948 13491 39004
rect 13547 38948 13615 39004
rect 13671 38948 13739 39004
rect 13795 38948 13863 39004
rect 13919 38948 13987 39004
rect 14043 38948 14111 39004
rect 14167 38948 14235 39004
rect 14291 38948 14359 39004
rect 14415 38948 14483 39004
rect 14539 38948 14607 39004
rect 14663 38948 14673 39004
rect 12861 38880 14673 38948
rect 12861 38824 12871 38880
rect 12927 38824 12995 38880
rect 13051 38824 13119 38880
rect 13175 38824 13243 38880
rect 13299 38824 13367 38880
rect 13423 38824 13491 38880
rect 13547 38824 13615 38880
rect 13671 38824 13739 38880
rect 13795 38824 13863 38880
rect 13919 38824 13987 38880
rect 14043 38824 14111 38880
rect 14167 38824 14235 38880
rect 14291 38824 14359 38880
rect 14415 38824 14483 38880
rect 14539 38824 14607 38880
rect 14663 38824 14673 38880
rect 12861 38756 14673 38824
rect 12861 38700 12871 38756
rect 12927 38700 12995 38756
rect 13051 38700 13119 38756
rect 13175 38700 13243 38756
rect 13299 38700 13367 38756
rect 13423 38700 13491 38756
rect 13547 38700 13615 38756
rect 13671 38700 13739 38756
rect 13795 38700 13863 38756
rect 13919 38700 13987 38756
rect 14043 38700 14111 38756
rect 14167 38700 14235 38756
rect 14291 38700 14359 38756
rect 14415 38700 14483 38756
rect 14539 38700 14607 38756
rect 14663 38700 14673 38756
rect 12861 38632 14673 38700
rect 12861 38576 12871 38632
rect 12927 38576 12995 38632
rect 13051 38576 13119 38632
rect 13175 38576 13243 38632
rect 13299 38576 13367 38632
rect 13423 38576 13491 38632
rect 13547 38576 13615 38632
rect 13671 38576 13739 38632
rect 13795 38576 13863 38632
rect 13919 38576 13987 38632
rect 14043 38576 14111 38632
rect 14167 38576 14235 38632
rect 14291 38576 14359 38632
rect 14415 38576 14483 38632
rect 14539 38576 14607 38632
rect 14663 38576 14673 38632
rect 12861 38508 14673 38576
rect 12861 38452 12871 38508
rect 12927 38452 12995 38508
rect 13051 38452 13119 38508
rect 13175 38452 13243 38508
rect 13299 38452 13367 38508
rect 13423 38452 13491 38508
rect 13547 38452 13615 38508
rect 13671 38452 13739 38508
rect 13795 38452 13863 38508
rect 13919 38452 13987 38508
rect 14043 38452 14111 38508
rect 14167 38452 14235 38508
rect 14291 38452 14359 38508
rect 14415 38452 14483 38508
rect 14539 38452 14607 38508
rect 14663 38452 14673 38508
rect 12861 38442 14673 38452
rect 2279 38079 2289 38135
rect 2345 38079 2355 38135
rect 2279 38003 2355 38079
rect 2279 37947 2289 38003
rect 2345 37947 2355 38003
rect 2279 37871 2355 37947
rect 2279 37815 2289 37871
rect 2345 37815 2355 37871
rect 2279 37739 2355 37815
rect 2279 37683 2289 37739
rect 2345 37683 2355 37739
rect 2279 37607 2355 37683
rect 2279 37551 2289 37607
rect 2345 37551 2355 37607
rect 2279 37475 2355 37551
rect 2279 37419 2289 37475
rect 2345 37419 2355 37475
rect 2279 37343 2355 37419
rect 2279 37287 2289 37343
rect 2345 37287 2355 37343
rect 2279 37211 2355 37287
rect 2279 37155 2289 37211
rect 2345 37155 2355 37211
rect 2279 37079 2355 37155
rect 2279 37023 2289 37079
rect 2345 37023 2355 37079
rect 2279 36947 2355 37023
rect 2279 36891 2289 36947
rect 2345 36891 2355 36947
rect 2279 36800 2355 36891
rect 14892 38176 14989 38200
rect 14892 36824 14902 38176
rect 14958 36824 14989 38176
rect 14892 36800 14989 36824
rect 2481 36554 2681 36564
rect 2481 36498 2491 36554
rect 2547 36498 2615 36554
rect 2671 36498 2681 36554
rect 2481 36430 2681 36498
rect 2481 36374 2491 36430
rect 2547 36374 2615 36430
rect 2671 36374 2681 36430
rect 2481 36306 2681 36374
rect 2481 36250 2491 36306
rect 2547 36250 2615 36306
rect 2671 36250 2681 36306
rect 2481 36182 2681 36250
rect 2481 36126 2491 36182
rect 2547 36126 2615 36182
rect 2671 36126 2681 36182
rect 2481 36058 2681 36126
rect 2481 36002 2491 36058
rect 2547 36002 2615 36058
rect 2671 36002 2681 36058
rect 2481 35934 2681 36002
rect 2481 35878 2491 35934
rect 2547 35878 2615 35934
rect 2671 35878 2681 35934
rect 2481 35810 2681 35878
rect 2481 35754 2491 35810
rect 2547 35754 2615 35810
rect 2671 35754 2681 35810
rect 2481 35686 2681 35754
rect 2481 35630 2491 35686
rect 2547 35630 2615 35686
rect 2671 35630 2681 35686
rect 2481 35562 2681 35630
rect 2481 35506 2491 35562
rect 2547 35506 2615 35562
rect 2671 35506 2681 35562
rect 2481 35438 2681 35506
rect 2481 35382 2491 35438
rect 2547 35382 2615 35438
rect 2671 35382 2681 35438
rect 2481 35314 2681 35382
rect 2481 35258 2491 35314
rect 2547 35258 2615 35314
rect 2671 35258 2681 35314
rect 2481 35190 2681 35258
rect 2481 35134 2491 35190
rect 2547 35134 2615 35190
rect 2671 35134 2681 35190
rect 2481 35066 2681 35134
rect 2481 35010 2491 35066
rect 2547 35010 2615 35066
rect 2671 35010 2681 35066
rect 2481 34942 2681 35010
rect 2481 34886 2491 34942
rect 2547 34886 2615 34942
rect 2671 34886 2681 34942
rect 2481 34818 2681 34886
rect 2481 34762 2491 34818
rect 2547 34762 2615 34818
rect 2671 34762 2681 34818
rect 2481 34694 2681 34762
rect 2481 34638 2491 34694
rect 2547 34638 2615 34694
rect 2671 34638 2681 34694
rect 2481 34570 2681 34638
rect 2481 34514 2491 34570
rect 2547 34514 2615 34570
rect 2671 34514 2681 34570
rect 2481 34446 2681 34514
rect 2481 34390 2491 34446
rect 2547 34390 2615 34446
rect 2671 34390 2681 34446
rect 2481 34322 2681 34390
rect 2481 34266 2491 34322
rect 2547 34266 2615 34322
rect 2671 34266 2681 34322
rect 2481 34198 2681 34266
rect 2481 34142 2491 34198
rect 2547 34142 2615 34198
rect 2671 34142 2681 34198
rect 2481 34074 2681 34142
rect 2481 34018 2491 34074
rect 2547 34018 2615 34074
rect 2671 34018 2681 34074
rect 2481 33950 2681 34018
rect 2481 33894 2491 33950
rect 2547 33894 2615 33950
rect 2671 33894 2681 33950
rect 2481 33826 2681 33894
rect 2481 33770 2491 33826
rect 2547 33770 2615 33826
rect 2671 33770 2681 33826
rect 2481 33702 2681 33770
rect 2481 33646 2491 33702
rect 2547 33646 2615 33702
rect 2671 33646 2681 33702
rect 2481 33636 2681 33646
rect 4851 36554 5051 36564
rect 4851 36498 4861 36554
rect 4917 36498 4985 36554
rect 5041 36498 5051 36554
rect 4851 36430 5051 36498
rect 4851 36374 4861 36430
rect 4917 36374 4985 36430
rect 5041 36374 5051 36430
rect 4851 36306 5051 36374
rect 4851 36250 4861 36306
rect 4917 36250 4985 36306
rect 5041 36250 5051 36306
rect 4851 36182 5051 36250
rect 4851 36126 4861 36182
rect 4917 36126 4985 36182
rect 5041 36126 5051 36182
rect 4851 36058 5051 36126
rect 4851 36002 4861 36058
rect 4917 36002 4985 36058
rect 5041 36002 5051 36058
rect 4851 35934 5051 36002
rect 4851 35878 4861 35934
rect 4917 35878 4985 35934
rect 5041 35878 5051 35934
rect 4851 35810 5051 35878
rect 4851 35754 4861 35810
rect 4917 35754 4985 35810
rect 5041 35754 5051 35810
rect 4851 35686 5051 35754
rect 4851 35630 4861 35686
rect 4917 35630 4985 35686
rect 5041 35630 5051 35686
rect 4851 35562 5051 35630
rect 4851 35506 4861 35562
rect 4917 35506 4985 35562
rect 5041 35506 5051 35562
rect 4851 35438 5051 35506
rect 4851 35382 4861 35438
rect 4917 35382 4985 35438
rect 5041 35382 5051 35438
rect 4851 35314 5051 35382
rect 4851 35258 4861 35314
rect 4917 35258 4985 35314
rect 5041 35258 5051 35314
rect 4851 35190 5051 35258
rect 4851 35134 4861 35190
rect 4917 35134 4985 35190
rect 5041 35134 5051 35190
rect 4851 35066 5051 35134
rect 4851 35010 4861 35066
rect 4917 35010 4985 35066
rect 5041 35010 5051 35066
rect 4851 34942 5051 35010
rect 4851 34886 4861 34942
rect 4917 34886 4985 34942
rect 5041 34886 5051 34942
rect 4851 34818 5051 34886
rect 4851 34762 4861 34818
rect 4917 34762 4985 34818
rect 5041 34762 5051 34818
rect 4851 34694 5051 34762
rect 4851 34638 4861 34694
rect 4917 34638 4985 34694
rect 5041 34638 5051 34694
rect 4851 34570 5051 34638
rect 4851 34514 4861 34570
rect 4917 34514 4985 34570
rect 5041 34514 5051 34570
rect 4851 34446 5051 34514
rect 4851 34390 4861 34446
rect 4917 34390 4985 34446
rect 5041 34390 5051 34446
rect 4851 34322 5051 34390
rect 4851 34266 4861 34322
rect 4917 34266 4985 34322
rect 5041 34266 5051 34322
rect 4851 34198 5051 34266
rect 4851 34142 4861 34198
rect 4917 34142 4985 34198
rect 5041 34142 5051 34198
rect 4851 34074 5051 34142
rect 4851 34018 4861 34074
rect 4917 34018 4985 34074
rect 5041 34018 5051 34074
rect 4851 33950 5051 34018
rect 4851 33894 4861 33950
rect 4917 33894 4985 33950
rect 5041 33894 5051 33950
rect 4851 33826 5051 33894
rect 4851 33770 4861 33826
rect 4917 33770 4985 33826
rect 5041 33770 5051 33826
rect 4851 33702 5051 33770
rect 4851 33646 4861 33702
rect 4917 33646 4985 33702
rect 5041 33646 5051 33702
rect 4851 33636 5051 33646
rect 7265 36554 7713 36564
rect 7265 36498 7275 36554
rect 7331 36498 7399 36554
rect 7455 36498 7523 36554
rect 7579 36498 7647 36554
rect 7703 36498 7713 36554
rect 7265 36430 7713 36498
rect 7265 36374 7275 36430
rect 7331 36374 7399 36430
rect 7455 36374 7523 36430
rect 7579 36374 7647 36430
rect 7703 36374 7713 36430
rect 7265 36306 7713 36374
rect 7265 36250 7275 36306
rect 7331 36250 7399 36306
rect 7455 36250 7523 36306
rect 7579 36250 7647 36306
rect 7703 36250 7713 36306
rect 7265 36182 7713 36250
rect 7265 36126 7275 36182
rect 7331 36126 7399 36182
rect 7455 36126 7523 36182
rect 7579 36126 7647 36182
rect 7703 36126 7713 36182
rect 7265 36058 7713 36126
rect 7265 36002 7275 36058
rect 7331 36002 7399 36058
rect 7455 36002 7523 36058
rect 7579 36002 7647 36058
rect 7703 36002 7713 36058
rect 7265 35934 7713 36002
rect 7265 35878 7275 35934
rect 7331 35878 7399 35934
rect 7455 35878 7523 35934
rect 7579 35878 7647 35934
rect 7703 35878 7713 35934
rect 7265 35810 7713 35878
rect 7265 35754 7275 35810
rect 7331 35754 7399 35810
rect 7455 35754 7523 35810
rect 7579 35754 7647 35810
rect 7703 35754 7713 35810
rect 7265 35686 7713 35754
rect 7265 35630 7275 35686
rect 7331 35630 7399 35686
rect 7455 35630 7523 35686
rect 7579 35630 7647 35686
rect 7703 35630 7713 35686
rect 7265 35562 7713 35630
rect 7265 35506 7275 35562
rect 7331 35506 7399 35562
rect 7455 35506 7523 35562
rect 7579 35506 7647 35562
rect 7703 35506 7713 35562
rect 7265 35438 7713 35506
rect 7265 35382 7275 35438
rect 7331 35382 7399 35438
rect 7455 35382 7523 35438
rect 7579 35382 7647 35438
rect 7703 35382 7713 35438
rect 7265 35314 7713 35382
rect 7265 35258 7275 35314
rect 7331 35258 7399 35314
rect 7455 35258 7523 35314
rect 7579 35258 7647 35314
rect 7703 35258 7713 35314
rect 7265 35190 7713 35258
rect 7265 35134 7275 35190
rect 7331 35134 7399 35190
rect 7455 35134 7523 35190
rect 7579 35134 7647 35190
rect 7703 35134 7713 35190
rect 7265 35066 7713 35134
rect 7265 35010 7275 35066
rect 7331 35010 7399 35066
rect 7455 35010 7523 35066
rect 7579 35010 7647 35066
rect 7703 35010 7713 35066
rect 7265 34942 7713 35010
rect 7265 34886 7275 34942
rect 7331 34886 7399 34942
rect 7455 34886 7523 34942
rect 7579 34886 7647 34942
rect 7703 34886 7713 34942
rect 7265 34818 7713 34886
rect 7265 34762 7275 34818
rect 7331 34762 7399 34818
rect 7455 34762 7523 34818
rect 7579 34762 7647 34818
rect 7703 34762 7713 34818
rect 7265 34694 7713 34762
rect 7265 34638 7275 34694
rect 7331 34638 7399 34694
rect 7455 34638 7523 34694
rect 7579 34638 7647 34694
rect 7703 34638 7713 34694
rect 7265 34570 7713 34638
rect 7265 34514 7275 34570
rect 7331 34514 7399 34570
rect 7455 34514 7523 34570
rect 7579 34514 7647 34570
rect 7703 34514 7713 34570
rect 7265 34446 7713 34514
rect 7265 34390 7275 34446
rect 7331 34390 7399 34446
rect 7455 34390 7523 34446
rect 7579 34390 7647 34446
rect 7703 34390 7713 34446
rect 7265 34322 7713 34390
rect 7265 34266 7275 34322
rect 7331 34266 7399 34322
rect 7455 34266 7523 34322
rect 7579 34266 7647 34322
rect 7703 34266 7713 34322
rect 7265 34198 7713 34266
rect 7265 34142 7275 34198
rect 7331 34142 7399 34198
rect 7455 34142 7523 34198
rect 7579 34142 7647 34198
rect 7703 34142 7713 34198
rect 7265 34074 7713 34142
rect 7265 34018 7275 34074
rect 7331 34018 7399 34074
rect 7455 34018 7523 34074
rect 7579 34018 7647 34074
rect 7703 34018 7713 34074
rect 7265 33950 7713 34018
rect 7265 33894 7275 33950
rect 7331 33894 7399 33950
rect 7455 33894 7523 33950
rect 7579 33894 7647 33950
rect 7703 33894 7713 33950
rect 7265 33826 7713 33894
rect 7265 33770 7275 33826
rect 7331 33770 7399 33826
rect 7455 33770 7523 33826
rect 7579 33770 7647 33826
rect 7703 33770 7713 33826
rect 7265 33702 7713 33770
rect 7265 33646 7275 33702
rect 7331 33646 7399 33702
rect 7455 33646 7523 33702
rect 7579 33646 7647 33702
rect 7703 33646 7713 33702
rect 7265 33636 7713 33646
rect 9927 36554 10127 36564
rect 9927 36498 9937 36554
rect 9993 36498 10061 36554
rect 10117 36498 10127 36554
rect 9927 36430 10127 36498
rect 9927 36374 9937 36430
rect 9993 36374 10061 36430
rect 10117 36374 10127 36430
rect 9927 36306 10127 36374
rect 9927 36250 9937 36306
rect 9993 36250 10061 36306
rect 10117 36250 10127 36306
rect 9927 36182 10127 36250
rect 9927 36126 9937 36182
rect 9993 36126 10061 36182
rect 10117 36126 10127 36182
rect 9927 36058 10127 36126
rect 9927 36002 9937 36058
rect 9993 36002 10061 36058
rect 10117 36002 10127 36058
rect 9927 35934 10127 36002
rect 9927 35878 9937 35934
rect 9993 35878 10061 35934
rect 10117 35878 10127 35934
rect 9927 35810 10127 35878
rect 9927 35754 9937 35810
rect 9993 35754 10061 35810
rect 10117 35754 10127 35810
rect 9927 35686 10127 35754
rect 9927 35630 9937 35686
rect 9993 35630 10061 35686
rect 10117 35630 10127 35686
rect 9927 35562 10127 35630
rect 9927 35506 9937 35562
rect 9993 35506 10061 35562
rect 10117 35506 10127 35562
rect 9927 35438 10127 35506
rect 9927 35382 9937 35438
rect 9993 35382 10061 35438
rect 10117 35382 10127 35438
rect 9927 35314 10127 35382
rect 9927 35258 9937 35314
rect 9993 35258 10061 35314
rect 10117 35258 10127 35314
rect 9927 35190 10127 35258
rect 9927 35134 9937 35190
rect 9993 35134 10061 35190
rect 10117 35134 10127 35190
rect 9927 35066 10127 35134
rect 9927 35010 9937 35066
rect 9993 35010 10061 35066
rect 10117 35010 10127 35066
rect 9927 34942 10127 35010
rect 9927 34886 9937 34942
rect 9993 34886 10061 34942
rect 10117 34886 10127 34942
rect 9927 34818 10127 34886
rect 9927 34762 9937 34818
rect 9993 34762 10061 34818
rect 10117 34762 10127 34818
rect 9927 34694 10127 34762
rect 9927 34638 9937 34694
rect 9993 34638 10061 34694
rect 10117 34638 10127 34694
rect 9927 34570 10127 34638
rect 9927 34514 9937 34570
rect 9993 34514 10061 34570
rect 10117 34514 10127 34570
rect 9927 34446 10127 34514
rect 9927 34390 9937 34446
rect 9993 34390 10061 34446
rect 10117 34390 10127 34446
rect 9927 34322 10127 34390
rect 9927 34266 9937 34322
rect 9993 34266 10061 34322
rect 10117 34266 10127 34322
rect 9927 34198 10127 34266
rect 9927 34142 9937 34198
rect 9993 34142 10061 34198
rect 10117 34142 10127 34198
rect 9927 34074 10127 34142
rect 9927 34018 9937 34074
rect 9993 34018 10061 34074
rect 10117 34018 10127 34074
rect 9927 33950 10127 34018
rect 9927 33894 9937 33950
rect 9993 33894 10061 33950
rect 10117 33894 10127 33950
rect 9927 33826 10127 33894
rect 9927 33770 9937 33826
rect 9993 33770 10061 33826
rect 10117 33770 10127 33826
rect 9927 33702 10127 33770
rect 9927 33646 9937 33702
rect 9993 33646 10061 33702
rect 10117 33646 10127 33702
rect 9927 33636 10127 33646
rect 12297 36554 12497 36564
rect 12297 36498 12307 36554
rect 12363 36498 12431 36554
rect 12487 36498 12497 36554
rect 12297 36430 12497 36498
rect 12297 36374 12307 36430
rect 12363 36374 12431 36430
rect 12487 36374 12497 36430
rect 12297 36306 12497 36374
rect 12297 36250 12307 36306
rect 12363 36250 12431 36306
rect 12487 36250 12497 36306
rect 12297 36182 12497 36250
rect 12297 36126 12307 36182
rect 12363 36126 12431 36182
rect 12487 36126 12497 36182
rect 12297 36058 12497 36126
rect 12297 36002 12307 36058
rect 12363 36002 12431 36058
rect 12487 36002 12497 36058
rect 12297 35934 12497 36002
rect 12297 35878 12307 35934
rect 12363 35878 12431 35934
rect 12487 35878 12497 35934
rect 12297 35810 12497 35878
rect 12297 35754 12307 35810
rect 12363 35754 12431 35810
rect 12487 35754 12497 35810
rect 12297 35686 12497 35754
rect 12297 35630 12307 35686
rect 12363 35630 12431 35686
rect 12487 35630 12497 35686
rect 12297 35562 12497 35630
rect 12297 35506 12307 35562
rect 12363 35506 12431 35562
rect 12487 35506 12497 35562
rect 12297 35438 12497 35506
rect 12297 35382 12307 35438
rect 12363 35382 12431 35438
rect 12487 35382 12497 35438
rect 12297 35314 12497 35382
rect 12297 35258 12307 35314
rect 12363 35258 12431 35314
rect 12487 35258 12497 35314
rect 12297 35190 12497 35258
rect 12297 35134 12307 35190
rect 12363 35134 12431 35190
rect 12487 35134 12497 35190
rect 12297 35066 12497 35134
rect 12297 35010 12307 35066
rect 12363 35010 12431 35066
rect 12487 35010 12497 35066
rect 12297 34942 12497 35010
rect 12297 34886 12307 34942
rect 12363 34886 12431 34942
rect 12487 34886 12497 34942
rect 12297 34818 12497 34886
rect 12297 34762 12307 34818
rect 12363 34762 12431 34818
rect 12487 34762 12497 34818
rect 12297 34694 12497 34762
rect 12297 34638 12307 34694
rect 12363 34638 12431 34694
rect 12487 34638 12497 34694
rect 12297 34570 12497 34638
rect 12297 34514 12307 34570
rect 12363 34514 12431 34570
rect 12487 34514 12497 34570
rect 12297 34446 12497 34514
rect 12297 34390 12307 34446
rect 12363 34390 12431 34446
rect 12487 34390 12497 34446
rect 12297 34322 12497 34390
rect 12297 34266 12307 34322
rect 12363 34266 12431 34322
rect 12487 34266 12497 34322
rect 12297 34198 12497 34266
rect 12297 34142 12307 34198
rect 12363 34142 12431 34198
rect 12487 34142 12497 34198
rect 12297 34074 12497 34142
rect 12297 34018 12307 34074
rect 12363 34018 12431 34074
rect 12487 34018 12497 34074
rect 12297 33950 12497 34018
rect 12297 33894 12307 33950
rect 12363 33894 12431 33950
rect 12487 33894 12497 33950
rect 12297 33826 12497 33894
rect 12297 33770 12307 33826
rect 12363 33770 12431 33826
rect 12487 33770 12497 33826
rect 12297 33702 12497 33770
rect 12297 33646 12307 33702
rect 12363 33646 12431 33702
rect 12487 33646 12497 33702
rect 12297 33636 12497 33646
rect 305 33354 2117 33364
rect 305 33298 315 33354
rect 371 33298 439 33354
rect 495 33298 563 33354
rect 619 33298 687 33354
rect 743 33298 811 33354
rect 867 33298 935 33354
rect 991 33298 1059 33354
rect 1115 33298 1183 33354
rect 1239 33298 1307 33354
rect 1363 33298 1431 33354
rect 1487 33298 1555 33354
rect 1611 33298 1679 33354
rect 1735 33298 1803 33354
rect 1859 33298 1927 33354
rect 1983 33298 2051 33354
rect 2107 33298 2117 33354
rect 305 33230 2117 33298
rect 305 33174 315 33230
rect 371 33174 439 33230
rect 495 33174 563 33230
rect 619 33174 687 33230
rect 743 33174 811 33230
rect 867 33174 935 33230
rect 991 33174 1059 33230
rect 1115 33174 1183 33230
rect 1239 33174 1307 33230
rect 1363 33174 1431 33230
rect 1487 33174 1555 33230
rect 1611 33174 1679 33230
rect 1735 33174 1803 33230
rect 1859 33174 1927 33230
rect 1983 33174 2051 33230
rect 2107 33174 2117 33230
rect 305 33106 2117 33174
rect 305 33050 315 33106
rect 371 33050 439 33106
rect 495 33050 563 33106
rect 619 33050 687 33106
rect 743 33050 811 33106
rect 867 33050 935 33106
rect 991 33050 1059 33106
rect 1115 33050 1183 33106
rect 1239 33050 1307 33106
rect 1363 33050 1431 33106
rect 1487 33050 1555 33106
rect 1611 33050 1679 33106
rect 1735 33050 1803 33106
rect 1859 33050 1927 33106
rect 1983 33050 2051 33106
rect 2107 33050 2117 33106
rect 305 32982 2117 33050
rect 305 32926 315 32982
rect 371 32926 439 32982
rect 495 32926 563 32982
rect 619 32926 687 32982
rect 743 32926 811 32982
rect 867 32926 935 32982
rect 991 32926 1059 32982
rect 1115 32926 1183 32982
rect 1239 32926 1307 32982
rect 1363 32926 1431 32982
rect 1487 32926 1555 32982
rect 1611 32926 1679 32982
rect 1735 32926 1803 32982
rect 1859 32926 1927 32982
rect 1983 32926 2051 32982
rect 2107 32926 2117 32982
rect 305 32858 2117 32926
rect 305 32802 315 32858
rect 371 32802 439 32858
rect 495 32802 563 32858
rect 619 32802 687 32858
rect 743 32802 811 32858
rect 867 32802 935 32858
rect 991 32802 1059 32858
rect 1115 32802 1183 32858
rect 1239 32802 1307 32858
rect 1363 32802 1431 32858
rect 1487 32802 1555 32858
rect 1611 32802 1679 32858
rect 1735 32802 1803 32858
rect 1859 32802 1927 32858
rect 1983 32802 2051 32858
rect 2107 32802 2117 32858
rect 305 32734 2117 32802
rect 305 32678 315 32734
rect 371 32678 439 32734
rect 495 32678 563 32734
rect 619 32678 687 32734
rect 743 32678 811 32734
rect 867 32678 935 32734
rect 991 32678 1059 32734
rect 1115 32678 1183 32734
rect 1239 32678 1307 32734
rect 1363 32678 1431 32734
rect 1487 32678 1555 32734
rect 1611 32678 1679 32734
rect 1735 32678 1803 32734
rect 1859 32678 1927 32734
rect 1983 32678 2051 32734
rect 2107 32678 2117 32734
rect 305 32610 2117 32678
rect 305 32554 315 32610
rect 371 32554 439 32610
rect 495 32554 563 32610
rect 619 32554 687 32610
rect 743 32554 811 32610
rect 867 32554 935 32610
rect 991 32554 1059 32610
rect 1115 32554 1183 32610
rect 1239 32554 1307 32610
rect 1363 32554 1431 32610
rect 1487 32554 1555 32610
rect 1611 32554 1679 32610
rect 1735 32554 1803 32610
rect 1859 32554 1927 32610
rect 1983 32554 2051 32610
rect 2107 32554 2117 32610
rect 305 32486 2117 32554
rect 305 32430 315 32486
rect 371 32430 439 32486
rect 495 32430 563 32486
rect 619 32430 687 32486
rect 743 32430 811 32486
rect 867 32430 935 32486
rect 991 32430 1059 32486
rect 1115 32430 1183 32486
rect 1239 32430 1307 32486
rect 1363 32430 1431 32486
rect 1487 32430 1555 32486
rect 1611 32430 1679 32486
rect 1735 32430 1803 32486
rect 1859 32430 1927 32486
rect 1983 32430 2051 32486
rect 2107 32430 2117 32486
rect 305 32362 2117 32430
rect 305 32306 315 32362
rect 371 32306 439 32362
rect 495 32306 563 32362
rect 619 32306 687 32362
rect 743 32306 811 32362
rect 867 32306 935 32362
rect 991 32306 1059 32362
rect 1115 32306 1183 32362
rect 1239 32306 1307 32362
rect 1363 32306 1431 32362
rect 1487 32306 1555 32362
rect 1611 32306 1679 32362
rect 1735 32306 1803 32362
rect 1859 32306 1927 32362
rect 1983 32306 2051 32362
rect 2107 32306 2117 32362
rect 305 32238 2117 32306
rect 305 32182 315 32238
rect 371 32182 439 32238
rect 495 32182 563 32238
rect 619 32182 687 32238
rect 743 32182 811 32238
rect 867 32182 935 32238
rect 991 32182 1059 32238
rect 1115 32182 1183 32238
rect 1239 32182 1307 32238
rect 1363 32182 1431 32238
rect 1487 32182 1555 32238
rect 1611 32182 1679 32238
rect 1735 32182 1803 32238
rect 1859 32182 1927 32238
rect 1983 32182 2051 32238
rect 2107 32182 2117 32238
rect 305 32114 2117 32182
rect 305 32058 315 32114
rect 371 32058 439 32114
rect 495 32058 563 32114
rect 619 32058 687 32114
rect 743 32058 811 32114
rect 867 32058 935 32114
rect 991 32058 1059 32114
rect 1115 32058 1183 32114
rect 1239 32058 1307 32114
rect 1363 32058 1431 32114
rect 1487 32058 1555 32114
rect 1611 32058 1679 32114
rect 1735 32058 1803 32114
rect 1859 32058 1927 32114
rect 1983 32058 2051 32114
rect 2107 32058 2117 32114
rect 305 31990 2117 32058
rect 305 31934 315 31990
rect 371 31934 439 31990
rect 495 31934 563 31990
rect 619 31934 687 31990
rect 743 31934 811 31990
rect 867 31934 935 31990
rect 991 31934 1059 31990
rect 1115 31934 1183 31990
rect 1239 31934 1307 31990
rect 1363 31934 1431 31990
rect 1487 31934 1555 31990
rect 1611 31934 1679 31990
rect 1735 31934 1803 31990
rect 1859 31934 1927 31990
rect 1983 31934 2051 31990
rect 2107 31934 2117 31990
rect 305 31866 2117 31934
rect 305 31810 315 31866
rect 371 31810 439 31866
rect 495 31810 563 31866
rect 619 31810 687 31866
rect 743 31810 811 31866
rect 867 31810 935 31866
rect 991 31810 1059 31866
rect 1115 31810 1183 31866
rect 1239 31810 1307 31866
rect 1363 31810 1431 31866
rect 1487 31810 1555 31866
rect 1611 31810 1679 31866
rect 1735 31810 1803 31866
rect 1859 31810 1927 31866
rect 1983 31810 2051 31866
rect 2107 31810 2117 31866
rect 305 31742 2117 31810
rect 305 31686 315 31742
rect 371 31686 439 31742
rect 495 31686 563 31742
rect 619 31686 687 31742
rect 743 31686 811 31742
rect 867 31686 935 31742
rect 991 31686 1059 31742
rect 1115 31686 1183 31742
rect 1239 31686 1307 31742
rect 1363 31686 1431 31742
rect 1487 31686 1555 31742
rect 1611 31686 1679 31742
rect 1735 31686 1803 31742
rect 1859 31686 1927 31742
rect 1983 31686 2051 31742
rect 2107 31686 2117 31742
rect 305 31618 2117 31686
rect 305 31562 315 31618
rect 371 31562 439 31618
rect 495 31562 563 31618
rect 619 31562 687 31618
rect 743 31562 811 31618
rect 867 31562 935 31618
rect 991 31562 1059 31618
rect 1115 31562 1183 31618
rect 1239 31562 1307 31618
rect 1363 31562 1431 31618
rect 1487 31562 1555 31618
rect 1611 31562 1679 31618
rect 1735 31562 1803 31618
rect 1859 31562 1927 31618
rect 1983 31562 2051 31618
rect 2107 31562 2117 31618
rect 305 31494 2117 31562
rect 305 31438 315 31494
rect 371 31438 439 31494
rect 495 31438 563 31494
rect 619 31438 687 31494
rect 743 31438 811 31494
rect 867 31438 935 31494
rect 991 31438 1059 31494
rect 1115 31438 1183 31494
rect 1239 31438 1307 31494
rect 1363 31438 1431 31494
rect 1487 31438 1555 31494
rect 1611 31438 1679 31494
rect 1735 31438 1803 31494
rect 1859 31438 1927 31494
rect 1983 31438 2051 31494
rect 2107 31438 2117 31494
rect 305 31370 2117 31438
rect 305 31314 315 31370
rect 371 31314 439 31370
rect 495 31314 563 31370
rect 619 31314 687 31370
rect 743 31314 811 31370
rect 867 31314 935 31370
rect 991 31314 1059 31370
rect 1115 31314 1183 31370
rect 1239 31314 1307 31370
rect 1363 31314 1431 31370
rect 1487 31314 1555 31370
rect 1611 31314 1679 31370
rect 1735 31314 1803 31370
rect 1859 31314 1927 31370
rect 1983 31314 2051 31370
rect 2107 31314 2117 31370
rect 305 31246 2117 31314
rect 305 31190 315 31246
rect 371 31190 439 31246
rect 495 31190 563 31246
rect 619 31190 687 31246
rect 743 31190 811 31246
rect 867 31190 935 31246
rect 991 31190 1059 31246
rect 1115 31190 1183 31246
rect 1239 31190 1307 31246
rect 1363 31190 1431 31246
rect 1487 31190 1555 31246
rect 1611 31190 1679 31246
rect 1735 31190 1803 31246
rect 1859 31190 1927 31246
rect 1983 31190 2051 31246
rect 2107 31190 2117 31246
rect 305 31122 2117 31190
rect 305 31066 315 31122
rect 371 31066 439 31122
rect 495 31066 563 31122
rect 619 31066 687 31122
rect 743 31066 811 31122
rect 867 31066 935 31122
rect 991 31066 1059 31122
rect 1115 31066 1183 31122
rect 1239 31066 1307 31122
rect 1363 31066 1431 31122
rect 1487 31066 1555 31122
rect 1611 31066 1679 31122
rect 1735 31066 1803 31122
rect 1859 31066 1927 31122
rect 1983 31066 2051 31122
rect 2107 31066 2117 31122
rect 305 30998 2117 31066
rect 305 30942 315 30998
rect 371 30942 439 30998
rect 495 30942 563 30998
rect 619 30942 687 30998
rect 743 30942 811 30998
rect 867 30942 935 30998
rect 991 30942 1059 30998
rect 1115 30942 1183 30998
rect 1239 30942 1307 30998
rect 1363 30942 1431 30998
rect 1487 30942 1555 30998
rect 1611 30942 1679 30998
rect 1735 30942 1803 30998
rect 1859 30942 1927 30998
rect 1983 30942 2051 30998
rect 2107 30942 2117 30998
rect 305 30874 2117 30942
rect 305 30818 315 30874
rect 371 30818 439 30874
rect 495 30818 563 30874
rect 619 30818 687 30874
rect 743 30818 811 30874
rect 867 30818 935 30874
rect 991 30818 1059 30874
rect 1115 30818 1183 30874
rect 1239 30818 1307 30874
rect 1363 30818 1431 30874
rect 1487 30818 1555 30874
rect 1611 30818 1679 30874
rect 1735 30818 1803 30874
rect 1859 30818 1927 30874
rect 1983 30818 2051 30874
rect 2107 30818 2117 30874
rect 305 30750 2117 30818
rect 305 30694 315 30750
rect 371 30694 439 30750
rect 495 30694 563 30750
rect 619 30694 687 30750
rect 743 30694 811 30750
rect 867 30694 935 30750
rect 991 30694 1059 30750
rect 1115 30694 1183 30750
rect 1239 30694 1307 30750
rect 1363 30694 1431 30750
rect 1487 30694 1555 30750
rect 1611 30694 1679 30750
rect 1735 30694 1803 30750
rect 1859 30694 1927 30750
rect 1983 30694 2051 30750
rect 2107 30694 2117 30750
rect 305 30626 2117 30694
rect 305 30570 315 30626
rect 371 30570 439 30626
rect 495 30570 563 30626
rect 619 30570 687 30626
rect 743 30570 811 30626
rect 867 30570 935 30626
rect 991 30570 1059 30626
rect 1115 30570 1183 30626
rect 1239 30570 1307 30626
rect 1363 30570 1431 30626
rect 1487 30570 1555 30626
rect 1611 30570 1679 30626
rect 1735 30570 1803 30626
rect 1859 30570 1927 30626
rect 1983 30570 2051 30626
rect 2107 30570 2117 30626
rect 305 30502 2117 30570
rect 305 30446 315 30502
rect 371 30446 439 30502
rect 495 30446 563 30502
rect 619 30446 687 30502
rect 743 30446 811 30502
rect 867 30446 935 30502
rect 991 30446 1059 30502
rect 1115 30446 1183 30502
rect 1239 30446 1307 30502
rect 1363 30446 1431 30502
rect 1487 30446 1555 30502
rect 1611 30446 1679 30502
rect 1735 30446 1803 30502
rect 1859 30446 1927 30502
rect 1983 30446 2051 30502
rect 2107 30446 2117 30502
rect 305 30436 2117 30446
rect 2798 33354 4734 33364
rect 2798 33298 2808 33354
rect 2864 33298 2932 33354
rect 2988 33298 3056 33354
rect 3112 33298 3180 33354
rect 3236 33298 3304 33354
rect 3360 33298 3428 33354
rect 3484 33298 3552 33354
rect 3608 33298 3676 33354
rect 3732 33298 3800 33354
rect 3856 33298 3924 33354
rect 3980 33298 4048 33354
rect 4104 33298 4172 33354
rect 4228 33298 4296 33354
rect 4352 33298 4420 33354
rect 4476 33298 4544 33354
rect 4600 33298 4668 33354
rect 4724 33298 4734 33354
rect 2798 33230 4734 33298
rect 2798 33174 2808 33230
rect 2864 33174 2932 33230
rect 2988 33174 3056 33230
rect 3112 33174 3180 33230
rect 3236 33174 3304 33230
rect 3360 33174 3428 33230
rect 3484 33174 3552 33230
rect 3608 33174 3676 33230
rect 3732 33174 3800 33230
rect 3856 33174 3924 33230
rect 3980 33174 4048 33230
rect 4104 33174 4172 33230
rect 4228 33174 4296 33230
rect 4352 33174 4420 33230
rect 4476 33174 4544 33230
rect 4600 33174 4668 33230
rect 4724 33174 4734 33230
rect 2798 33106 4734 33174
rect 2798 33050 2808 33106
rect 2864 33050 2932 33106
rect 2988 33050 3056 33106
rect 3112 33050 3180 33106
rect 3236 33050 3304 33106
rect 3360 33050 3428 33106
rect 3484 33050 3552 33106
rect 3608 33050 3676 33106
rect 3732 33050 3800 33106
rect 3856 33050 3924 33106
rect 3980 33050 4048 33106
rect 4104 33050 4172 33106
rect 4228 33050 4296 33106
rect 4352 33050 4420 33106
rect 4476 33050 4544 33106
rect 4600 33050 4668 33106
rect 4724 33050 4734 33106
rect 2798 32982 4734 33050
rect 2798 32926 2808 32982
rect 2864 32926 2932 32982
rect 2988 32926 3056 32982
rect 3112 32926 3180 32982
rect 3236 32926 3304 32982
rect 3360 32926 3428 32982
rect 3484 32926 3552 32982
rect 3608 32926 3676 32982
rect 3732 32926 3800 32982
rect 3856 32926 3924 32982
rect 3980 32926 4048 32982
rect 4104 32926 4172 32982
rect 4228 32926 4296 32982
rect 4352 32926 4420 32982
rect 4476 32926 4544 32982
rect 4600 32926 4668 32982
rect 4724 32926 4734 32982
rect 2798 32858 4734 32926
rect 2798 32802 2808 32858
rect 2864 32802 2932 32858
rect 2988 32802 3056 32858
rect 3112 32802 3180 32858
rect 3236 32802 3304 32858
rect 3360 32802 3428 32858
rect 3484 32802 3552 32858
rect 3608 32802 3676 32858
rect 3732 32802 3800 32858
rect 3856 32802 3924 32858
rect 3980 32802 4048 32858
rect 4104 32802 4172 32858
rect 4228 32802 4296 32858
rect 4352 32802 4420 32858
rect 4476 32802 4544 32858
rect 4600 32802 4668 32858
rect 4724 32802 4734 32858
rect 2798 32734 4734 32802
rect 2798 32678 2808 32734
rect 2864 32678 2932 32734
rect 2988 32678 3056 32734
rect 3112 32678 3180 32734
rect 3236 32678 3304 32734
rect 3360 32678 3428 32734
rect 3484 32678 3552 32734
rect 3608 32678 3676 32734
rect 3732 32678 3800 32734
rect 3856 32678 3924 32734
rect 3980 32678 4048 32734
rect 4104 32678 4172 32734
rect 4228 32678 4296 32734
rect 4352 32678 4420 32734
rect 4476 32678 4544 32734
rect 4600 32678 4668 32734
rect 4724 32678 4734 32734
rect 2798 32610 4734 32678
rect 2798 32554 2808 32610
rect 2864 32554 2932 32610
rect 2988 32554 3056 32610
rect 3112 32554 3180 32610
rect 3236 32554 3304 32610
rect 3360 32554 3428 32610
rect 3484 32554 3552 32610
rect 3608 32554 3676 32610
rect 3732 32554 3800 32610
rect 3856 32554 3924 32610
rect 3980 32554 4048 32610
rect 4104 32554 4172 32610
rect 4228 32554 4296 32610
rect 4352 32554 4420 32610
rect 4476 32554 4544 32610
rect 4600 32554 4668 32610
rect 4724 32554 4734 32610
rect 2798 32486 4734 32554
rect 2798 32430 2808 32486
rect 2864 32430 2932 32486
rect 2988 32430 3056 32486
rect 3112 32430 3180 32486
rect 3236 32430 3304 32486
rect 3360 32430 3428 32486
rect 3484 32430 3552 32486
rect 3608 32430 3676 32486
rect 3732 32430 3800 32486
rect 3856 32430 3924 32486
rect 3980 32430 4048 32486
rect 4104 32430 4172 32486
rect 4228 32430 4296 32486
rect 4352 32430 4420 32486
rect 4476 32430 4544 32486
rect 4600 32430 4668 32486
rect 4724 32430 4734 32486
rect 2798 32362 4734 32430
rect 2798 32306 2808 32362
rect 2864 32306 2932 32362
rect 2988 32306 3056 32362
rect 3112 32306 3180 32362
rect 3236 32306 3304 32362
rect 3360 32306 3428 32362
rect 3484 32306 3552 32362
rect 3608 32306 3676 32362
rect 3732 32306 3800 32362
rect 3856 32306 3924 32362
rect 3980 32306 4048 32362
rect 4104 32306 4172 32362
rect 4228 32306 4296 32362
rect 4352 32306 4420 32362
rect 4476 32306 4544 32362
rect 4600 32306 4668 32362
rect 4724 32306 4734 32362
rect 2798 32238 4734 32306
rect 2798 32182 2808 32238
rect 2864 32182 2932 32238
rect 2988 32182 3056 32238
rect 3112 32182 3180 32238
rect 3236 32182 3304 32238
rect 3360 32182 3428 32238
rect 3484 32182 3552 32238
rect 3608 32182 3676 32238
rect 3732 32182 3800 32238
rect 3856 32182 3924 32238
rect 3980 32182 4048 32238
rect 4104 32182 4172 32238
rect 4228 32182 4296 32238
rect 4352 32182 4420 32238
rect 4476 32182 4544 32238
rect 4600 32182 4668 32238
rect 4724 32182 4734 32238
rect 2798 32114 4734 32182
rect 2798 32058 2808 32114
rect 2864 32058 2932 32114
rect 2988 32058 3056 32114
rect 3112 32058 3180 32114
rect 3236 32058 3304 32114
rect 3360 32058 3428 32114
rect 3484 32058 3552 32114
rect 3608 32058 3676 32114
rect 3732 32058 3800 32114
rect 3856 32058 3924 32114
rect 3980 32058 4048 32114
rect 4104 32058 4172 32114
rect 4228 32058 4296 32114
rect 4352 32058 4420 32114
rect 4476 32058 4544 32114
rect 4600 32058 4668 32114
rect 4724 32058 4734 32114
rect 2798 31990 4734 32058
rect 2798 31934 2808 31990
rect 2864 31934 2932 31990
rect 2988 31934 3056 31990
rect 3112 31934 3180 31990
rect 3236 31934 3304 31990
rect 3360 31934 3428 31990
rect 3484 31934 3552 31990
rect 3608 31934 3676 31990
rect 3732 31934 3800 31990
rect 3856 31934 3924 31990
rect 3980 31934 4048 31990
rect 4104 31934 4172 31990
rect 4228 31934 4296 31990
rect 4352 31934 4420 31990
rect 4476 31934 4544 31990
rect 4600 31934 4668 31990
rect 4724 31934 4734 31990
rect 2798 31866 4734 31934
rect 2798 31810 2808 31866
rect 2864 31810 2932 31866
rect 2988 31810 3056 31866
rect 3112 31810 3180 31866
rect 3236 31810 3304 31866
rect 3360 31810 3428 31866
rect 3484 31810 3552 31866
rect 3608 31810 3676 31866
rect 3732 31810 3800 31866
rect 3856 31810 3924 31866
rect 3980 31810 4048 31866
rect 4104 31810 4172 31866
rect 4228 31810 4296 31866
rect 4352 31810 4420 31866
rect 4476 31810 4544 31866
rect 4600 31810 4668 31866
rect 4724 31810 4734 31866
rect 2798 31742 4734 31810
rect 2798 31686 2808 31742
rect 2864 31686 2932 31742
rect 2988 31686 3056 31742
rect 3112 31686 3180 31742
rect 3236 31686 3304 31742
rect 3360 31686 3428 31742
rect 3484 31686 3552 31742
rect 3608 31686 3676 31742
rect 3732 31686 3800 31742
rect 3856 31686 3924 31742
rect 3980 31686 4048 31742
rect 4104 31686 4172 31742
rect 4228 31686 4296 31742
rect 4352 31686 4420 31742
rect 4476 31686 4544 31742
rect 4600 31686 4668 31742
rect 4724 31686 4734 31742
rect 2798 31618 4734 31686
rect 2798 31562 2808 31618
rect 2864 31562 2932 31618
rect 2988 31562 3056 31618
rect 3112 31562 3180 31618
rect 3236 31562 3304 31618
rect 3360 31562 3428 31618
rect 3484 31562 3552 31618
rect 3608 31562 3676 31618
rect 3732 31562 3800 31618
rect 3856 31562 3924 31618
rect 3980 31562 4048 31618
rect 4104 31562 4172 31618
rect 4228 31562 4296 31618
rect 4352 31562 4420 31618
rect 4476 31562 4544 31618
rect 4600 31562 4668 31618
rect 4724 31562 4734 31618
rect 2798 31494 4734 31562
rect 2798 31438 2808 31494
rect 2864 31438 2932 31494
rect 2988 31438 3056 31494
rect 3112 31438 3180 31494
rect 3236 31438 3304 31494
rect 3360 31438 3428 31494
rect 3484 31438 3552 31494
rect 3608 31438 3676 31494
rect 3732 31438 3800 31494
rect 3856 31438 3924 31494
rect 3980 31438 4048 31494
rect 4104 31438 4172 31494
rect 4228 31438 4296 31494
rect 4352 31438 4420 31494
rect 4476 31438 4544 31494
rect 4600 31438 4668 31494
rect 4724 31438 4734 31494
rect 2798 31370 4734 31438
rect 2798 31314 2808 31370
rect 2864 31314 2932 31370
rect 2988 31314 3056 31370
rect 3112 31314 3180 31370
rect 3236 31314 3304 31370
rect 3360 31314 3428 31370
rect 3484 31314 3552 31370
rect 3608 31314 3676 31370
rect 3732 31314 3800 31370
rect 3856 31314 3924 31370
rect 3980 31314 4048 31370
rect 4104 31314 4172 31370
rect 4228 31314 4296 31370
rect 4352 31314 4420 31370
rect 4476 31314 4544 31370
rect 4600 31314 4668 31370
rect 4724 31314 4734 31370
rect 2798 31246 4734 31314
rect 2798 31190 2808 31246
rect 2864 31190 2932 31246
rect 2988 31190 3056 31246
rect 3112 31190 3180 31246
rect 3236 31190 3304 31246
rect 3360 31190 3428 31246
rect 3484 31190 3552 31246
rect 3608 31190 3676 31246
rect 3732 31190 3800 31246
rect 3856 31190 3924 31246
rect 3980 31190 4048 31246
rect 4104 31190 4172 31246
rect 4228 31190 4296 31246
rect 4352 31190 4420 31246
rect 4476 31190 4544 31246
rect 4600 31190 4668 31246
rect 4724 31190 4734 31246
rect 2798 31122 4734 31190
rect 2798 31066 2808 31122
rect 2864 31066 2932 31122
rect 2988 31066 3056 31122
rect 3112 31066 3180 31122
rect 3236 31066 3304 31122
rect 3360 31066 3428 31122
rect 3484 31066 3552 31122
rect 3608 31066 3676 31122
rect 3732 31066 3800 31122
rect 3856 31066 3924 31122
rect 3980 31066 4048 31122
rect 4104 31066 4172 31122
rect 4228 31066 4296 31122
rect 4352 31066 4420 31122
rect 4476 31066 4544 31122
rect 4600 31066 4668 31122
rect 4724 31066 4734 31122
rect 2798 30998 4734 31066
rect 2798 30942 2808 30998
rect 2864 30942 2932 30998
rect 2988 30942 3056 30998
rect 3112 30942 3180 30998
rect 3236 30942 3304 30998
rect 3360 30942 3428 30998
rect 3484 30942 3552 30998
rect 3608 30942 3676 30998
rect 3732 30942 3800 30998
rect 3856 30942 3924 30998
rect 3980 30942 4048 30998
rect 4104 30942 4172 30998
rect 4228 30942 4296 30998
rect 4352 30942 4420 30998
rect 4476 30942 4544 30998
rect 4600 30942 4668 30998
rect 4724 30942 4734 30998
rect 2798 30874 4734 30942
rect 2798 30818 2808 30874
rect 2864 30818 2932 30874
rect 2988 30818 3056 30874
rect 3112 30818 3180 30874
rect 3236 30818 3304 30874
rect 3360 30818 3428 30874
rect 3484 30818 3552 30874
rect 3608 30818 3676 30874
rect 3732 30818 3800 30874
rect 3856 30818 3924 30874
rect 3980 30818 4048 30874
rect 4104 30818 4172 30874
rect 4228 30818 4296 30874
rect 4352 30818 4420 30874
rect 4476 30818 4544 30874
rect 4600 30818 4668 30874
rect 4724 30818 4734 30874
rect 2798 30750 4734 30818
rect 2798 30694 2808 30750
rect 2864 30694 2932 30750
rect 2988 30694 3056 30750
rect 3112 30694 3180 30750
rect 3236 30694 3304 30750
rect 3360 30694 3428 30750
rect 3484 30694 3552 30750
rect 3608 30694 3676 30750
rect 3732 30694 3800 30750
rect 3856 30694 3924 30750
rect 3980 30694 4048 30750
rect 4104 30694 4172 30750
rect 4228 30694 4296 30750
rect 4352 30694 4420 30750
rect 4476 30694 4544 30750
rect 4600 30694 4668 30750
rect 4724 30694 4734 30750
rect 2798 30626 4734 30694
rect 2798 30570 2808 30626
rect 2864 30570 2932 30626
rect 2988 30570 3056 30626
rect 3112 30570 3180 30626
rect 3236 30570 3304 30626
rect 3360 30570 3428 30626
rect 3484 30570 3552 30626
rect 3608 30570 3676 30626
rect 3732 30570 3800 30626
rect 3856 30570 3924 30626
rect 3980 30570 4048 30626
rect 4104 30570 4172 30626
rect 4228 30570 4296 30626
rect 4352 30570 4420 30626
rect 4476 30570 4544 30626
rect 4600 30570 4668 30626
rect 4724 30570 4734 30626
rect 2798 30502 4734 30570
rect 2798 30446 2808 30502
rect 2864 30446 2932 30502
rect 2988 30446 3056 30502
rect 3112 30446 3180 30502
rect 3236 30446 3304 30502
rect 3360 30446 3428 30502
rect 3484 30446 3552 30502
rect 3608 30446 3676 30502
rect 3732 30446 3800 30502
rect 3856 30446 3924 30502
rect 3980 30446 4048 30502
rect 4104 30446 4172 30502
rect 4228 30446 4296 30502
rect 4352 30446 4420 30502
rect 4476 30446 4544 30502
rect 4600 30446 4668 30502
rect 4724 30446 4734 30502
rect 2798 30436 4734 30446
rect 5168 33354 7104 33364
rect 5168 33298 5178 33354
rect 5234 33298 5302 33354
rect 5358 33298 5426 33354
rect 5482 33298 5550 33354
rect 5606 33298 5674 33354
rect 5730 33298 5798 33354
rect 5854 33298 5922 33354
rect 5978 33298 6046 33354
rect 6102 33298 6170 33354
rect 6226 33298 6294 33354
rect 6350 33298 6418 33354
rect 6474 33298 6542 33354
rect 6598 33298 6666 33354
rect 6722 33298 6790 33354
rect 6846 33298 6914 33354
rect 6970 33298 7038 33354
rect 7094 33298 7104 33354
rect 5168 33230 7104 33298
rect 5168 33174 5178 33230
rect 5234 33174 5302 33230
rect 5358 33174 5426 33230
rect 5482 33174 5550 33230
rect 5606 33174 5674 33230
rect 5730 33174 5798 33230
rect 5854 33174 5922 33230
rect 5978 33174 6046 33230
rect 6102 33174 6170 33230
rect 6226 33174 6294 33230
rect 6350 33174 6418 33230
rect 6474 33174 6542 33230
rect 6598 33174 6666 33230
rect 6722 33174 6790 33230
rect 6846 33174 6914 33230
rect 6970 33174 7038 33230
rect 7094 33174 7104 33230
rect 5168 33106 7104 33174
rect 5168 33050 5178 33106
rect 5234 33050 5302 33106
rect 5358 33050 5426 33106
rect 5482 33050 5550 33106
rect 5606 33050 5674 33106
rect 5730 33050 5798 33106
rect 5854 33050 5922 33106
rect 5978 33050 6046 33106
rect 6102 33050 6170 33106
rect 6226 33050 6294 33106
rect 6350 33050 6418 33106
rect 6474 33050 6542 33106
rect 6598 33050 6666 33106
rect 6722 33050 6790 33106
rect 6846 33050 6914 33106
rect 6970 33050 7038 33106
rect 7094 33050 7104 33106
rect 5168 32982 7104 33050
rect 5168 32926 5178 32982
rect 5234 32926 5302 32982
rect 5358 32926 5426 32982
rect 5482 32926 5550 32982
rect 5606 32926 5674 32982
rect 5730 32926 5798 32982
rect 5854 32926 5922 32982
rect 5978 32926 6046 32982
rect 6102 32926 6170 32982
rect 6226 32926 6294 32982
rect 6350 32926 6418 32982
rect 6474 32926 6542 32982
rect 6598 32926 6666 32982
rect 6722 32926 6790 32982
rect 6846 32926 6914 32982
rect 6970 32926 7038 32982
rect 7094 32926 7104 32982
rect 5168 32858 7104 32926
rect 5168 32802 5178 32858
rect 5234 32802 5302 32858
rect 5358 32802 5426 32858
rect 5482 32802 5550 32858
rect 5606 32802 5674 32858
rect 5730 32802 5798 32858
rect 5854 32802 5922 32858
rect 5978 32802 6046 32858
rect 6102 32802 6170 32858
rect 6226 32802 6294 32858
rect 6350 32802 6418 32858
rect 6474 32802 6542 32858
rect 6598 32802 6666 32858
rect 6722 32802 6790 32858
rect 6846 32802 6914 32858
rect 6970 32802 7038 32858
rect 7094 32802 7104 32858
rect 5168 32734 7104 32802
rect 5168 32678 5178 32734
rect 5234 32678 5302 32734
rect 5358 32678 5426 32734
rect 5482 32678 5550 32734
rect 5606 32678 5674 32734
rect 5730 32678 5798 32734
rect 5854 32678 5922 32734
rect 5978 32678 6046 32734
rect 6102 32678 6170 32734
rect 6226 32678 6294 32734
rect 6350 32678 6418 32734
rect 6474 32678 6542 32734
rect 6598 32678 6666 32734
rect 6722 32678 6790 32734
rect 6846 32678 6914 32734
rect 6970 32678 7038 32734
rect 7094 32678 7104 32734
rect 5168 32610 7104 32678
rect 5168 32554 5178 32610
rect 5234 32554 5302 32610
rect 5358 32554 5426 32610
rect 5482 32554 5550 32610
rect 5606 32554 5674 32610
rect 5730 32554 5798 32610
rect 5854 32554 5922 32610
rect 5978 32554 6046 32610
rect 6102 32554 6170 32610
rect 6226 32554 6294 32610
rect 6350 32554 6418 32610
rect 6474 32554 6542 32610
rect 6598 32554 6666 32610
rect 6722 32554 6790 32610
rect 6846 32554 6914 32610
rect 6970 32554 7038 32610
rect 7094 32554 7104 32610
rect 5168 32486 7104 32554
rect 5168 32430 5178 32486
rect 5234 32430 5302 32486
rect 5358 32430 5426 32486
rect 5482 32430 5550 32486
rect 5606 32430 5674 32486
rect 5730 32430 5798 32486
rect 5854 32430 5922 32486
rect 5978 32430 6046 32486
rect 6102 32430 6170 32486
rect 6226 32430 6294 32486
rect 6350 32430 6418 32486
rect 6474 32430 6542 32486
rect 6598 32430 6666 32486
rect 6722 32430 6790 32486
rect 6846 32430 6914 32486
rect 6970 32430 7038 32486
rect 7094 32430 7104 32486
rect 5168 32362 7104 32430
rect 5168 32306 5178 32362
rect 5234 32306 5302 32362
rect 5358 32306 5426 32362
rect 5482 32306 5550 32362
rect 5606 32306 5674 32362
rect 5730 32306 5798 32362
rect 5854 32306 5922 32362
rect 5978 32306 6046 32362
rect 6102 32306 6170 32362
rect 6226 32306 6294 32362
rect 6350 32306 6418 32362
rect 6474 32306 6542 32362
rect 6598 32306 6666 32362
rect 6722 32306 6790 32362
rect 6846 32306 6914 32362
rect 6970 32306 7038 32362
rect 7094 32306 7104 32362
rect 5168 32238 7104 32306
rect 5168 32182 5178 32238
rect 5234 32182 5302 32238
rect 5358 32182 5426 32238
rect 5482 32182 5550 32238
rect 5606 32182 5674 32238
rect 5730 32182 5798 32238
rect 5854 32182 5922 32238
rect 5978 32182 6046 32238
rect 6102 32182 6170 32238
rect 6226 32182 6294 32238
rect 6350 32182 6418 32238
rect 6474 32182 6542 32238
rect 6598 32182 6666 32238
rect 6722 32182 6790 32238
rect 6846 32182 6914 32238
rect 6970 32182 7038 32238
rect 7094 32182 7104 32238
rect 5168 32114 7104 32182
rect 5168 32058 5178 32114
rect 5234 32058 5302 32114
rect 5358 32058 5426 32114
rect 5482 32058 5550 32114
rect 5606 32058 5674 32114
rect 5730 32058 5798 32114
rect 5854 32058 5922 32114
rect 5978 32058 6046 32114
rect 6102 32058 6170 32114
rect 6226 32058 6294 32114
rect 6350 32058 6418 32114
rect 6474 32058 6542 32114
rect 6598 32058 6666 32114
rect 6722 32058 6790 32114
rect 6846 32058 6914 32114
rect 6970 32058 7038 32114
rect 7094 32058 7104 32114
rect 5168 31990 7104 32058
rect 5168 31934 5178 31990
rect 5234 31934 5302 31990
rect 5358 31934 5426 31990
rect 5482 31934 5550 31990
rect 5606 31934 5674 31990
rect 5730 31934 5798 31990
rect 5854 31934 5922 31990
rect 5978 31934 6046 31990
rect 6102 31934 6170 31990
rect 6226 31934 6294 31990
rect 6350 31934 6418 31990
rect 6474 31934 6542 31990
rect 6598 31934 6666 31990
rect 6722 31934 6790 31990
rect 6846 31934 6914 31990
rect 6970 31934 7038 31990
rect 7094 31934 7104 31990
rect 5168 31866 7104 31934
rect 5168 31810 5178 31866
rect 5234 31810 5302 31866
rect 5358 31810 5426 31866
rect 5482 31810 5550 31866
rect 5606 31810 5674 31866
rect 5730 31810 5798 31866
rect 5854 31810 5922 31866
rect 5978 31810 6046 31866
rect 6102 31810 6170 31866
rect 6226 31810 6294 31866
rect 6350 31810 6418 31866
rect 6474 31810 6542 31866
rect 6598 31810 6666 31866
rect 6722 31810 6790 31866
rect 6846 31810 6914 31866
rect 6970 31810 7038 31866
rect 7094 31810 7104 31866
rect 5168 31742 7104 31810
rect 5168 31686 5178 31742
rect 5234 31686 5302 31742
rect 5358 31686 5426 31742
rect 5482 31686 5550 31742
rect 5606 31686 5674 31742
rect 5730 31686 5798 31742
rect 5854 31686 5922 31742
rect 5978 31686 6046 31742
rect 6102 31686 6170 31742
rect 6226 31686 6294 31742
rect 6350 31686 6418 31742
rect 6474 31686 6542 31742
rect 6598 31686 6666 31742
rect 6722 31686 6790 31742
rect 6846 31686 6914 31742
rect 6970 31686 7038 31742
rect 7094 31686 7104 31742
rect 5168 31618 7104 31686
rect 5168 31562 5178 31618
rect 5234 31562 5302 31618
rect 5358 31562 5426 31618
rect 5482 31562 5550 31618
rect 5606 31562 5674 31618
rect 5730 31562 5798 31618
rect 5854 31562 5922 31618
rect 5978 31562 6046 31618
rect 6102 31562 6170 31618
rect 6226 31562 6294 31618
rect 6350 31562 6418 31618
rect 6474 31562 6542 31618
rect 6598 31562 6666 31618
rect 6722 31562 6790 31618
rect 6846 31562 6914 31618
rect 6970 31562 7038 31618
rect 7094 31562 7104 31618
rect 5168 31494 7104 31562
rect 5168 31438 5178 31494
rect 5234 31438 5302 31494
rect 5358 31438 5426 31494
rect 5482 31438 5550 31494
rect 5606 31438 5674 31494
rect 5730 31438 5798 31494
rect 5854 31438 5922 31494
rect 5978 31438 6046 31494
rect 6102 31438 6170 31494
rect 6226 31438 6294 31494
rect 6350 31438 6418 31494
rect 6474 31438 6542 31494
rect 6598 31438 6666 31494
rect 6722 31438 6790 31494
rect 6846 31438 6914 31494
rect 6970 31438 7038 31494
rect 7094 31438 7104 31494
rect 5168 31370 7104 31438
rect 5168 31314 5178 31370
rect 5234 31314 5302 31370
rect 5358 31314 5426 31370
rect 5482 31314 5550 31370
rect 5606 31314 5674 31370
rect 5730 31314 5798 31370
rect 5854 31314 5922 31370
rect 5978 31314 6046 31370
rect 6102 31314 6170 31370
rect 6226 31314 6294 31370
rect 6350 31314 6418 31370
rect 6474 31314 6542 31370
rect 6598 31314 6666 31370
rect 6722 31314 6790 31370
rect 6846 31314 6914 31370
rect 6970 31314 7038 31370
rect 7094 31314 7104 31370
rect 5168 31246 7104 31314
rect 5168 31190 5178 31246
rect 5234 31190 5302 31246
rect 5358 31190 5426 31246
rect 5482 31190 5550 31246
rect 5606 31190 5674 31246
rect 5730 31190 5798 31246
rect 5854 31190 5922 31246
rect 5978 31190 6046 31246
rect 6102 31190 6170 31246
rect 6226 31190 6294 31246
rect 6350 31190 6418 31246
rect 6474 31190 6542 31246
rect 6598 31190 6666 31246
rect 6722 31190 6790 31246
rect 6846 31190 6914 31246
rect 6970 31190 7038 31246
rect 7094 31190 7104 31246
rect 5168 31122 7104 31190
rect 5168 31066 5178 31122
rect 5234 31066 5302 31122
rect 5358 31066 5426 31122
rect 5482 31066 5550 31122
rect 5606 31066 5674 31122
rect 5730 31066 5798 31122
rect 5854 31066 5922 31122
rect 5978 31066 6046 31122
rect 6102 31066 6170 31122
rect 6226 31066 6294 31122
rect 6350 31066 6418 31122
rect 6474 31066 6542 31122
rect 6598 31066 6666 31122
rect 6722 31066 6790 31122
rect 6846 31066 6914 31122
rect 6970 31066 7038 31122
rect 7094 31066 7104 31122
rect 5168 30998 7104 31066
rect 5168 30942 5178 30998
rect 5234 30942 5302 30998
rect 5358 30942 5426 30998
rect 5482 30942 5550 30998
rect 5606 30942 5674 30998
rect 5730 30942 5798 30998
rect 5854 30942 5922 30998
rect 5978 30942 6046 30998
rect 6102 30942 6170 30998
rect 6226 30942 6294 30998
rect 6350 30942 6418 30998
rect 6474 30942 6542 30998
rect 6598 30942 6666 30998
rect 6722 30942 6790 30998
rect 6846 30942 6914 30998
rect 6970 30942 7038 30998
rect 7094 30942 7104 30998
rect 5168 30874 7104 30942
rect 5168 30818 5178 30874
rect 5234 30818 5302 30874
rect 5358 30818 5426 30874
rect 5482 30818 5550 30874
rect 5606 30818 5674 30874
rect 5730 30818 5798 30874
rect 5854 30818 5922 30874
rect 5978 30818 6046 30874
rect 6102 30818 6170 30874
rect 6226 30818 6294 30874
rect 6350 30818 6418 30874
rect 6474 30818 6542 30874
rect 6598 30818 6666 30874
rect 6722 30818 6790 30874
rect 6846 30818 6914 30874
rect 6970 30818 7038 30874
rect 7094 30818 7104 30874
rect 5168 30750 7104 30818
rect 5168 30694 5178 30750
rect 5234 30694 5302 30750
rect 5358 30694 5426 30750
rect 5482 30694 5550 30750
rect 5606 30694 5674 30750
rect 5730 30694 5798 30750
rect 5854 30694 5922 30750
rect 5978 30694 6046 30750
rect 6102 30694 6170 30750
rect 6226 30694 6294 30750
rect 6350 30694 6418 30750
rect 6474 30694 6542 30750
rect 6598 30694 6666 30750
rect 6722 30694 6790 30750
rect 6846 30694 6914 30750
rect 6970 30694 7038 30750
rect 7094 30694 7104 30750
rect 5168 30626 7104 30694
rect 5168 30570 5178 30626
rect 5234 30570 5302 30626
rect 5358 30570 5426 30626
rect 5482 30570 5550 30626
rect 5606 30570 5674 30626
rect 5730 30570 5798 30626
rect 5854 30570 5922 30626
rect 5978 30570 6046 30626
rect 6102 30570 6170 30626
rect 6226 30570 6294 30626
rect 6350 30570 6418 30626
rect 6474 30570 6542 30626
rect 6598 30570 6666 30626
rect 6722 30570 6790 30626
rect 6846 30570 6914 30626
rect 6970 30570 7038 30626
rect 7094 30570 7104 30626
rect 5168 30502 7104 30570
rect 5168 30446 5178 30502
rect 5234 30446 5302 30502
rect 5358 30446 5426 30502
rect 5482 30446 5550 30502
rect 5606 30446 5674 30502
rect 5730 30446 5798 30502
rect 5854 30446 5922 30502
rect 5978 30446 6046 30502
rect 6102 30446 6170 30502
rect 6226 30446 6294 30502
rect 6350 30446 6418 30502
rect 6474 30446 6542 30502
rect 6598 30446 6666 30502
rect 6722 30446 6790 30502
rect 6846 30446 6914 30502
rect 6970 30446 7038 30502
rect 7094 30446 7104 30502
rect 5168 30436 7104 30446
rect 7874 33354 9810 33364
rect 7874 33298 7884 33354
rect 7940 33298 8008 33354
rect 8064 33298 8132 33354
rect 8188 33298 8256 33354
rect 8312 33298 8380 33354
rect 8436 33298 8504 33354
rect 8560 33298 8628 33354
rect 8684 33298 8752 33354
rect 8808 33298 8876 33354
rect 8932 33298 9000 33354
rect 9056 33298 9124 33354
rect 9180 33298 9248 33354
rect 9304 33298 9372 33354
rect 9428 33298 9496 33354
rect 9552 33298 9620 33354
rect 9676 33298 9744 33354
rect 9800 33298 9810 33354
rect 7874 33230 9810 33298
rect 7874 33174 7884 33230
rect 7940 33174 8008 33230
rect 8064 33174 8132 33230
rect 8188 33174 8256 33230
rect 8312 33174 8380 33230
rect 8436 33174 8504 33230
rect 8560 33174 8628 33230
rect 8684 33174 8752 33230
rect 8808 33174 8876 33230
rect 8932 33174 9000 33230
rect 9056 33174 9124 33230
rect 9180 33174 9248 33230
rect 9304 33174 9372 33230
rect 9428 33174 9496 33230
rect 9552 33174 9620 33230
rect 9676 33174 9744 33230
rect 9800 33174 9810 33230
rect 7874 33106 9810 33174
rect 7874 33050 7884 33106
rect 7940 33050 8008 33106
rect 8064 33050 8132 33106
rect 8188 33050 8256 33106
rect 8312 33050 8380 33106
rect 8436 33050 8504 33106
rect 8560 33050 8628 33106
rect 8684 33050 8752 33106
rect 8808 33050 8876 33106
rect 8932 33050 9000 33106
rect 9056 33050 9124 33106
rect 9180 33050 9248 33106
rect 9304 33050 9372 33106
rect 9428 33050 9496 33106
rect 9552 33050 9620 33106
rect 9676 33050 9744 33106
rect 9800 33050 9810 33106
rect 7874 32982 9810 33050
rect 7874 32926 7884 32982
rect 7940 32926 8008 32982
rect 8064 32926 8132 32982
rect 8188 32926 8256 32982
rect 8312 32926 8380 32982
rect 8436 32926 8504 32982
rect 8560 32926 8628 32982
rect 8684 32926 8752 32982
rect 8808 32926 8876 32982
rect 8932 32926 9000 32982
rect 9056 32926 9124 32982
rect 9180 32926 9248 32982
rect 9304 32926 9372 32982
rect 9428 32926 9496 32982
rect 9552 32926 9620 32982
rect 9676 32926 9744 32982
rect 9800 32926 9810 32982
rect 7874 32858 9810 32926
rect 7874 32802 7884 32858
rect 7940 32802 8008 32858
rect 8064 32802 8132 32858
rect 8188 32802 8256 32858
rect 8312 32802 8380 32858
rect 8436 32802 8504 32858
rect 8560 32802 8628 32858
rect 8684 32802 8752 32858
rect 8808 32802 8876 32858
rect 8932 32802 9000 32858
rect 9056 32802 9124 32858
rect 9180 32802 9248 32858
rect 9304 32802 9372 32858
rect 9428 32802 9496 32858
rect 9552 32802 9620 32858
rect 9676 32802 9744 32858
rect 9800 32802 9810 32858
rect 7874 32734 9810 32802
rect 7874 32678 7884 32734
rect 7940 32678 8008 32734
rect 8064 32678 8132 32734
rect 8188 32678 8256 32734
rect 8312 32678 8380 32734
rect 8436 32678 8504 32734
rect 8560 32678 8628 32734
rect 8684 32678 8752 32734
rect 8808 32678 8876 32734
rect 8932 32678 9000 32734
rect 9056 32678 9124 32734
rect 9180 32678 9248 32734
rect 9304 32678 9372 32734
rect 9428 32678 9496 32734
rect 9552 32678 9620 32734
rect 9676 32678 9744 32734
rect 9800 32678 9810 32734
rect 7874 32610 9810 32678
rect 7874 32554 7884 32610
rect 7940 32554 8008 32610
rect 8064 32554 8132 32610
rect 8188 32554 8256 32610
rect 8312 32554 8380 32610
rect 8436 32554 8504 32610
rect 8560 32554 8628 32610
rect 8684 32554 8752 32610
rect 8808 32554 8876 32610
rect 8932 32554 9000 32610
rect 9056 32554 9124 32610
rect 9180 32554 9248 32610
rect 9304 32554 9372 32610
rect 9428 32554 9496 32610
rect 9552 32554 9620 32610
rect 9676 32554 9744 32610
rect 9800 32554 9810 32610
rect 7874 32486 9810 32554
rect 7874 32430 7884 32486
rect 7940 32430 8008 32486
rect 8064 32430 8132 32486
rect 8188 32430 8256 32486
rect 8312 32430 8380 32486
rect 8436 32430 8504 32486
rect 8560 32430 8628 32486
rect 8684 32430 8752 32486
rect 8808 32430 8876 32486
rect 8932 32430 9000 32486
rect 9056 32430 9124 32486
rect 9180 32430 9248 32486
rect 9304 32430 9372 32486
rect 9428 32430 9496 32486
rect 9552 32430 9620 32486
rect 9676 32430 9744 32486
rect 9800 32430 9810 32486
rect 7874 32362 9810 32430
rect 7874 32306 7884 32362
rect 7940 32306 8008 32362
rect 8064 32306 8132 32362
rect 8188 32306 8256 32362
rect 8312 32306 8380 32362
rect 8436 32306 8504 32362
rect 8560 32306 8628 32362
rect 8684 32306 8752 32362
rect 8808 32306 8876 32362
rect 8932 32306 9000 32362
rect 9056 32306 9124 32362
rect 9180 32306 9248 32362
rect 9304 32306 9372 32362
rect 9428 32306 9496 32362
rect 9552 32306 9620 32362
rect 9676 32306 9744 32362
rect 9800 32306 9810 32362
rect 7874 32238 9810 32306
rect 7874 32182 7884 32238
rect 7940 32182 8008 32238
rect 8064 32182 8132 32238
rect 8188 32182 8256 32238
rect 8312 32182 8380 32238
rect 8436 32182 8504 32238
rect 8560 32182 8628 32238
rect 8684 32182 8752 32238
rect 8808 32182 8876 32238
rect 8932 32182 9000 32238
rect 9056 32182 9124 32238
rect 9180 32182 9248 32238
rect 9304 32182 9372 32238
rect 9428 32182 9496 32238
rect 9552 32182 9620 32238
rect 9676 32182 9744 32238
rect 9800 32182 9810 32238
rect 7874 32114 9810 32182
rect 7874 32058 7884 32114
rect 7940 32058 8008 32114
rect 8064 32058 8132 32114
rect 8188 32058 8256 32114
rect 8312 32058 8380 32114
rect 8436 32058 8504 32114
rect 8560 32058 8628 32114
rect 8684 32058 8752 32114
rect 8808 32058 8876 32114
rect 8932 32058 9000 32114
rect 9056 32058 9124 32114
rect 9180 32058 9248 32114
rect 9304 32058 9372 32114
rect 9428 32058 9496 32114
rect 9552 32058 9620 32114
rect 9676 32058 9744 32114
rect 9800 32058 9810 32114
rect 7874 31990 9810 32058
rect 7874 31934 7884 31990
rect 7940 31934 8008 31990
rect 8064 31934 8132 31990
rect 8188 31934 8256 31990
rect 8312 31934 8380 31990
rect 8436 31934 8504 31990
rect 8560 31934 8628 31990
rect 8684 31934 8752 31990
rect 8808 31934 8876 31990
rect 8932 31934 9000 31990
rect 9056 31934 9124 31990
rect 9180 31934 9248 31990
rect 9304 31934 9372 31990
rect 9428 31934 9496 31990
rect 9552 31934 9620 31990
rect 9676 31934 9744 31990
rect 9800 31934 9810 31990
rect 7874 31866 9810 31934
rect 7874 31810 7884 31866
rect 7940 31810 8008 31866
rect 8064 31810 8132 31866
rect 8188 31810 8256 31866
rect 8312 31810 8380 31866
rect 8436 31810 8504 31866
rect 8560 31810 8628 31866
rect 8684 31810 8752 31866
rect 8808 31810 8876 31866
rect 8932 31810 9000 31866
rect 9056 31810 9124 31866
rect 9180 31810 9248 31866
rect 9304 31810 9372 31866
rect 9428 31810 9496 31866
rect 9552 31810 9620 31866
rect 9676 31810 9744 31866
rect 9800 31810 9810 31866
rect 7874 31742 9810 31810
rect 7874 31686 7884 31742
rect 7940 31686 8008 31742
rect 8064 31686 8132 31742
rect 8188 31686 8256 31742
rect 8312 31686 8380 31742
rect 8436 31686 8504 31742
rect 8560 31686 8628 31742
rect 8684 31686 8752 31742
rect 8808 31686 8876 31742
rect 8932 31686 9000 31742
rect 9056 31686 9124 31742
rect 9180 31686 9248 31742
rect 9304 31686 9372 31742
rect 9428 31686 9496 31742
rect 9552 31686 9620 31742
rect 9676 31686 9744 31742
rect 9800 31686 9810 31742
rect 7874 31618 9810 31686
rect 7874 31562 7884 31618
rect 7940 31562 8008 31618
rect 8064 31562 8132 31618
rect 8188 31562 8256 31618
rect 8312 31562 8380 31618
rect 8436 31562 8504 31618
rect 8560 31562 8628 31618
rect 8684 31562 8752 31618
rect 8808 31562 8876 31618
rect 8932 31562 9000 31618
rect 9056 31562 9124 31618
rect 9180 31562 9248 31618
rect 9304 31562 9372 31618
rect 9428 31562 9496 31618
rect 9552 31562 9620 31618
rect 9676 31562 9744 31618
rect 9800 31562 9810 31618
rect 7874 31494 9810 31562
rect 7874 31438 7884 31494
rect 7940 31438 8008 31494
rect 8064 31438 8132 31494
rect 8188 31438 8256 31494
rect 8312 31438 8380 31494
rect 8436 31438 8504 31494
rect 8560 31438 8628 31494
rect 8684 31438 8752 31494
rect 8808 31438 8876 31494
rect 8932 31438 9000 31494
rect 9056 31438 9124 31494
rect 9180 31438 9248 31494
rect 9304 31438 9372 31494
rect 9428 31438 9496 31494
rect 9552 31438 9620 31494
rect 9676 31438 9744 31494
rect 9800 31438 9810 31494
rect 7874 31370 9810 31438
rect 7874 31314 7884 31370
rect 7940 31314 8008 31370
rect 8064 31314 8132 31370
rect 8188 31314 8256 31370
rect 8312 31314 8380 31370
rect 8436 31314 8504 31370
rect 8560 31314 8628 31370
rect 8684 31314 8752 31370
rect 8808 31314 8876 31370
rect 8932 31314 9000 31370
rect 9056 31314 9124 31370
rect 9180 31314 9248 31370
rect 9304 31314 9372 31370
rect 9428 31314 9496 31370
rect 9552 31314 9620 31370
rect 9676 31314 9744 31370
rect 9800 31314 9810 31370
rect 7874 31246 9810 31314
rect 7874 31190 7884 31246
rect 7940 31190 8008 31246
rect 8064 31190 8132 31246
rect 8188 31190 8256 31246
rect 8312 31190 8380 31246
rect 8436 31190 8504 31246
rect 8560 31190 8628 31246
rect 8684 31190 8752 31246
rect 8808 31190 8876 31246
rect 8932 31190 9000 31246
rect 9056 31190 9124 31246
rect 9180 31190 9248 31246
rect 9304 31190 9372 31246
rect 9428 31190 9496 31246
rect 9552 31190 9620 31246
rect 9676 31190 9744 31246
rect 9800 31190 9810 31246
rect 7874 31122 9810 31190
rect 7874 31066 7884 31122
rect 7940 31066 8008 31122
rect 8064 31066 8132 31122
rect 8188 31066 8256 31122
rect 8312 31066 8380 31122
rect 8436 31066 8504 31122
rect 8560 31066 8628 31122
rect 8684 31066 8752 31122
rect 8808 31066 8876 31122
rect 8932 31066 9000 31122
rect 9056 31066 9124 31122
rect 9180 31066 9248 31122
rect 9304 31066 9372 31122
rect 9428 31066 9496 31122
rect 9552 31066 9620 31122
rect 9676 31066 9744 31122
rect 9800 31066 9810 31122
rect 7874 30998 9810 31066
rect 7874 30942 7884 30998
rect 7940 30942 8008 30998
rect 8064 30942 8132 30998
rect 8188 30942 8256 30998
rect 8312 30942 8380 30998
rect 8436 30942 8504 30998
rect 8560 30942 8628 30998
rect 8684 30942 8752 30998
rect 8808 30942 8876 30998
rect 8932 30942 9000 30998
rect 9056 30942 9124 30998
rect 9180 30942 9248 30998
rect 9304 30942 9372 30998
rect 9428 30942 9496 30998
rect 9552 30942 9620 30998
rect 9676 30942 9744 30998
rect 9800 30942 9810 30998
rect 7874 30874 9810 30942
rect 7874 30818 7884 30874
rect 7940 30818 8008 30874
rect 8064 30818 8132 30874
rect 8188 30818 8256 30874
rect 8312 30818 8380 30874
rect 8436 30818 8504 30874
rect 8560 30818 8628 30874
rect 8684 30818 8752 30874
rect 8808 30818 8876 30874
rect 8932 30818 9000 30874
rect 9056 30818 9124 30874
rect 9180 30818 9248 30874
rect 9304 30818 9372 30874
rect 9428 30818 9496 30874
rect 9552 30818 9620 30874
rect 9676 30818 9744 30874
rect 9800 30818 9810 30874
rect 7874 30750 9810 30818
rect 7874 30694 7884 30750
rect 7940 30694 8008 30750
rect 8064 30694 8132 30750
rect 8188 30694 8256 30750
rect 8312 30694 8380 30750
rect 8436 30694 8504 30750
rect 8560 30694 8628 30750
rect 8684 30694 8752 30750
rect 8808 30694 8876 30750
rect 8932 30694 9000 30750
rect 9056 30694 9124 30750
rect 9180 30694 9248 30750
rect 9304 30694 9372 30750
rect 9428 30694 9496 30750
rect 9552 30694 9620 30750
rect 9676 30694 9744 30750
rect 9800 30694 9810 30750
rect 7874 30626 9810 30694
rect 7874 30570 7884 30626
rect 7940 30570 8008 30626
rect 8064 30570 8132 30626
rect 8188 30570 8256 30626
rect 8312 30570 8380 30626
rect 8436 30570 8504 30626
rect 8560 30570 8628 30626
rect 8684 30570 8752 30626
rect 8808 30570 8876 30626
rect 8932 30570 9000 30626
rect 9056 30570 9124 30626
rect 9180 30570 9248 30626
rect 9304 30570 9372 30626
rect 9428 30570 9496 30626
rect 9552 30570 9620 30626
rect 9676 30570 9744 30626
rect 9800 30570 9810 30626
rect 7874 30502 9810 30570
rect 7874 30446 7884 30502
rect 7940 30446 8008 30502
rect 8064 30446 8132 30502
rect 8188 30446 8256 30502
rect 8312 30446 8380 30502
rect 8436 30446 8504 30502
rect 8560 30446 8628 30502
rect 8684 30446 8752 30502
rect 8808 30446 8876 30502
rect 8932 30446 9000 30502
rect 9056 30446 9124 30502
rect 9180 30446 9248 30502
rect 9304 30446 9372 30502
rect 9428 30446 9496 30502
rect 9552 30446 9620 30502
rect 9676 30446 9744 30502
rect 9800 30446 9810 30502
rect 7874 30436 9810 30446
rect 10244 33354 12180 33364
rect 10244 33298 10254 33354
rect 10310 33298 10378 33354
rect 10434 33298 10502 33354
rect 10558 33298 10626 33354
rect 10682 33298 10750 33354
rect 10806 33298 10874 33354
rect 10930 33298 10998 33354
rect 11054 33298 11122 33354
rect 11178 33298 11246 33354
rect 11302 33298 11370 33354
rect 11426 33298 11494 33354
rect 11550 33298 11618 33354
rect 11674 33298 11742 33354
rect 11798 33298 11866 33354
rect 11922 33298 11990 33354
rect 12046 33298 12114 33354
rect 12170 33298 12180 33354
rect 10244 33230 12180 33298
rect 10244 33174 10254 33230
rect 10310 33174 10378 33230
rect 10434 33174 10502 33230
rect 10558 33174 10626 33230
rect 10682 33174 10750 33230
rect 10806 33174 10874 33230
rect 10930 33174 10998 33230
rect 11054 33174 11122 33230
rect 11178 33174 11246 33230
rect 11302 33174 11370 33230
rect 11426 33174 11494 33230
rect 11550 33174 11618 33230
rect 11674 33174 11742 33230
rect 11798 33174 11866 33230
rect 11922 33174 11990 33230
rect 12046 33174 12114 33230
rect 12170 33174 12180 33230
rect 10244 33106 12180 33174
rect 10244 33050 10254 33106
rect 10310 33050 10378 33106
rect 10434 33050 10502 33106
rect 10558 33050 10626 33106
rect 10682 33050 10750 33106
rect 10806 33050 10874 33106
rect 10930 33050 10998 33106
rect 11054 33050 11122 33106
rect 11178 33050 11246 33106
rect 11302 33050 11370 33106
rect 11426 33050 11494 33106
rect 11550 33050 11618 33106
rect 11674 33050 11742 33106
rect 11798 33050 11866 33106
rect 11922 33050 11990 33106
rect 12046 33050 12114 33106
rect 12170 33050 12180 33106
rect 10244 32982 12180 33050
rect 10244 32926 10254 32982
rect 10310 32926 10378 32982
rect 10434 32926 10502 32982
rect 10558 32926 10626 32982
rect 10682 32926 10750 32982
rect 10806 32926 10874 32982
rect 10930 32926 10998 32982
rect 11054 32926 11122 32982
rect 11178 32926 11246 32982
rect 11302 32926 11370 32982
rect 11426 32926 11494 32982
rect 11550 32926 11618 32982
rect 11674 32926 11742 32982
rect 11798 32926 11866 32982
rect 11922 32926 11990 32982
rect 12046 32926 12114 32982
rect 12170 32926 12180 32982
rect 10244 32858 12180 32926
rect 10244 32802 10254 32858
rect 10310 32802 10378 32858
rect 10434 32802 10502 32858
rect 10558 32802 10626 32858
rect 10682 32802 10750 32858
rect 10806 32802 10874 32858
rect 10930 32802 10998 32858
rect 11054 32802 11122 32858
rect 11178 32802 11246 32858
rect 11302 32802 11370 32858
rect 11426 32802 11494 32858
rect 11550 32802 11618 32858
rect 11674 32802 11742 32858
rect 11798 32802 11866 32858
rect 11922 32802 11990 32858
rect 12046 32802 12114 32858
rect 12170 32802 12180 32858
rect 10244 32734 12180 32802
rect 10244 32678 10254 32734
rect 10310 32678 10378 32734
rect 10434 32678 10502 32734
rect 10558 32678 10626 32734
rect 10682 32678 10750 32734
rect 10806 32678 10874 32734
rect 10930 32678 10998 32734
rect 11054 32678 11122 32734
rect 11178 32678 11246 32734
rect 11302 32678 11370 32734
rect 11426 32678 11494 32734
rect 11550 32678 11618 32734
rect 11674 32678 11742 32734
rect 11798 32678 11866 32734
rect 11922 32678 11990 32734
rect 12046 32678 12114 32734
rect 12170 32678 12180 32734
rect 10244 32610 12180 32678
rect 10244 32554 10254 32610
rect 10310 32554 10378 32610
rect 10434 32554 10502 32610
rect 10558 32554 10626 32610
rect 10682 32554 10750 32610
rect 10806 32554 10874 32610
rect 10930 32554 10998 32610
rect 11054 32554 11122 32610
rect 11178 32554 11246 32610
rect 11302 32554 11370 32610
rect 11426 32554 11494 32610
rect 11550 32554 11618 32610
rect 11674 32554 11742 32610
rect 11798 32554 11866 32610
rect 11922 32554 11990 32610
rect 12046 32554 12114 32610
rect 12170 32554 12180 32610
rect 10244 32486 12180 32554
rect 10244 32430 10254 32486
rect 10310 32430 10378 32486
rect 10434 32430 10502 32486
rect 10558 32430 10626 32486
rect 10682 32430 10750 32486
rect 10806 32430 10874 32486
rect 10930 32430 10998 32486
rect 11054 32430 11122 32486
rect 11178 32430 11246 32486
rect 11302 32430 11370 32486
rect 11426 32430 11494 32486
rect 11550 32430 11618 32486
rect 11674 32430 11742 32486
rect 11798 32430 11866 32486
rect 11922 32430 11990 32486
rect 12046 32430 12114 32486
rect 12170 32430 12180 32486
rect 10244 32362 12180 32430
rect 10244 32306 10254 32362
rect 10310 32306 10378 32362
rect 10434 32306 10502 32362
rect 10558 32306 10626 32362
rect 10682 32306 10750 32362
rect 10806 32306 10874 32362
rect 10930 32306 10998 32362
rect 11054 32306 11122 32362
rect 11178 32306 11246 32362
rect 11302 32306 11370 32362
rect 11426 32306 11494 32362
rect 11550 32306 11618 32362
rect 11674 32306 11742 32362
rect 11798 32306 11866 32362
rect 11922 32306 11990 32362
rect 12046 32306 12114 32362
rect 12170 32306 12180 32362
rect 10244 32238 12180 32306
rect 10244 32182 10254 32238
rect 10310 32182 10378 32238
rect 10434 32182 10502 32238
rect 10558 32182 10626 32238
rect 10682 32182 10750 32238
rect 10806 32182 10874 32238
rect 10930 32182 10998 32238
rect 11054 32182 11122 32238
rect 11178 32182 11246 32238
rect 11302 32182 11370 32238
rect 11426 32182 11494 32238
rect 11550 32182 11618 32238
rect 11674 32182 11742 32238
rect 11798 32182 11866 32238
rect 11922 32182 11990 32238
rect 12046 32182 12114 32238
rect 12170 32182 12180 32238
rect 10244 32114 12180 32182
rect 10244 32058 10254 32114
rect 10310 32058 10378 32114
rect 10434 32058 10502 32114
rect 10558 32058 10626 32114
rect 10682 32058 10750 32114
rect 10806 32058 10874 32114
rect 10930 32058 10998 32114
rect 11054 32058 11122 32114
rect 11178 32058 11246 32114
rect 11302 32058 11370 32114
rect 11426 32058 11494 32114
rect 11550 32058 11618 32114
rect 11674 32058 11742 32114
rect 11798 32058 11866 32114
rect 11922 32058 11990 32114
rect 12046 32058 12114 32114
rect 12170 32058 12180 32114
rect 10244 31990 12180 32058
rect 10244 31934 10254 31990
rect 10310 31934 10378 31990
rect 10434 31934 10502 31990
rect 10558 31934 10626 31990
rect 10682 31934 10750 31990
rect 10806 31934 10874 31990
rect 10930 31934 10998 31990
rect 11054 31934 11122 31990
rect 11178 31934 11246 31990
rect 11302 31934 11370 31990
rect 11426 31934 11494 31990
rect 11550 31934 11618 31990
rect 11674 31934 11742 31990
rect 11798 31934 11866 31990
rect 11922 31934 11990 31990
rect 12046 31934 12114 31990
rect 12170 31934 12180 31990
rect 10244 31866 12180 31934
rect 10244 31810 10254 31866
rect 10310 31810 10378 31866
rect 10434 31810 10502 31866
rect 10558 31810 10626 31866
rect 10682 31810 10750 31866
rect 10806 31810 10874 31866
rect 10930 31810 10998 31866
rect 11054 31810 11122 31866
rect 11178 31810 11246 31866
rect 11302 31810 11370 31866
rect 11426 31810 11494 31866
rect 11550 31810 11618 31866
rect 11674 31810 11742 31866
rect 11798 31810 11866 31866
rect 11922 31810 11990 31866
rect 12046 31810 12114 31866
rect 12170 31810 12180 31866
rect 10244 31742 12180 31810
rect 10244 31686 10254 31742
rect 10310 31686 10378 31742
rect 10434 31686 10502 31742
rect 10558 31686 10626 31742
rect 10682 31686 10750 31742
rect 10806 31686 10874 31742
rect 10930 31686 10998 31742
rect 11054 31686 11122 31742
rect 11178 31686 11246 31742
rect 11302 31686 11370 31742
rect 11426 31686 11494 31742
rect 11550 31686 11618 31742
rect 11674 31686 11742 31742
rect 11798 31686 11866 31742
rect 11922 31686 11990 31742
rect 12046 31686 12114 31742
rect 12170 31686 12180 31742
rect 10244 31618 12180 31686
rect 10244 31562 10254 31618
rect 10310 31562 10378 31618
rect 10434 31562 10502 31618
rect 10558 31562 10626 31618
rect 10682 31562 10750 31618
rect 10806 31562 10874 31618
rect 10930 31562 10998 31618
rect 11054 31562 11122 31618
rect 11178 31562 11246 31618
rect 11302 31562 11370 31618
rect 11426 31562 11494 31618
rect 11550 31562 11618 31618
rect 11674 31562 11742 31618
rect 11798 31562 11866 31618
rect 11922 31562 11990 31618
rect 12046 31562 12114 31618
rect 12170 31562 12180 31618
rect 10244 31494 12180 31562
rect 10244 31438 10254 31494
rect 10310 31438 10378 31494
rect 10434 31438 10502 31494
rect 10558 31438 10626 31494
rect 10682 31438 10750 31494
rect 10806 31438 10874 31494
rect 10930 31438 10998 31494
rect 11054 31438 11122 31494
rect 11178 31438 11246 31494
rect 11302 31438 11370 31494
rect 11426 31438 11494 31494
rect 11550 31438 11618 31494
rect 11674 31438 11742 31494
rect 11798 31438 11866 31494
rect 11922 31438 11990 31494
rect 12046 31438 12114 31494
rect 12170 31438 12180 31494
rect 10244 31370 12180 31438
rect 10244 31314 10254 31370
rect 10310 31314 10378 31370
rect 10434 31314 10502 31370
rect 10558 31314 10626 31370
rect 10682 31314 10750 31370
rect 10806 31314 10874 31370
rect 10930 31314 10998 31370
rect 11054 31314 11122 31370
rect 11178 31314 11246 31370
rect 11302 31314 11370 31370
rect 11426 31314 11494 31370
rect 11550 31314 11618 31370
rect 11674 31314 11742 31370
rect 11798 31314 11866 31370
rect 11922 31314 11990 31370
rect 12046 31314 12114 31370
rect 12170 31314 12180 31370
rect 10244 31246 12180 31314
rect 10244 31190 10254 31246
rect 10310 31190 10378 31246
rect 10434 31190 10502 31246
rect 10558 31190 10626 31246
rect 10682 31190 10750 31246
rect 10806 31190 10874 31246
rect 10930 31190 10998 31246
rect 11054 31190 11122 31246
rect 11178 31190 11246 31246
rect 11302 31190 11370 31246
rect 11426 31190 11494 31246
rect 11550 31190 11618 31246
rect 11674 31190 11742 31246
rect 11798 31190 11866 31246
rect 11922 31190 11990 31246
rect 12046 31190 12114 31246
rect 12170 31190 12180 31246
rect 10244 31122 12180 31190
rect 10244 31066 10254 31122
rect 10310 31066 10378 31122
rect 10434 31066 10502 31122
rect 10558 31066 10626 31122
rect 10682 31066 10750 31122
rect 10806 31066 10874 31122
rect 10930 31066 10998 31122
rect 11054 31066 11122 31122
rect 11178 31066 11246 31122
rect 11302 31066 11370 31122
rect 11426 31066 11494 31122
rect 11550 31066 11618 31122
rect 11674 31066 11742 31122
rect 11798 31066 11866 31122
rect 11922 31066 11990 31122
rect 12046 31066 12114 31122
rect 12170 31066 12180 31122
rect 10244 30998 12180 31066
rect 10244 30942 10254 30998
rect 10310 30942 10378 30998
rect 10434 30942 10502 30998
rect 10558 30942 10626 30998
rect 10682 30942 10750 30998
rect 10806 30942 10874 30998
rect 10930 30942 10998 30998
rect 11054 30942 11122 30998
rect 11178 30942 11246 30998
rect 11302 30942 11370 30998
rect 11426 30942 11494 30998
rect 11550 30942 11618 30998
rect 11674 30942 11742 30998
rect 11798 30942 11866 30998
rect 11922 30942 11990 30998
rect 12046 30942 12114 30998
rect 12170 30942 12180 30998
rect 10244 30874 12180 30942
rect 10244 30818 10254 30874
rect 10310 30818 10378 30874
rect 10434 30818 10502 30874
rect 10558 30818 10626 30874
rect 10682 30818 10750 30874
rect 10806 30818 10874 30874
rect 10930 30818 10998 30874
rect 11054 30818 11122 30874
rect 11178 30818 11246 30874
rect 11302 30818 11370 30874
rect 11426 30818 11494 30874
rect 11550 30818 11618 30874
rect 11674 30818 11742 30874
rect 11798 30818 11866 30874
rect 11922 30818 11990 30874
rect 12046 30818 12114 30874
rect 12170 30818 12180 30874
rect 10244 30750 12180 30818
rect 10244 30694 10254 30750
rect 10310 30694 10378 30750
rect 10434 30694 10502 30750
rect 10558 30694 10626 30750
rect 10682 30694 10750 30750
rect 10806 30694 10874 30750
rect 10930 30694 10998 30750
rect 11054 30694 11122 30750
rect 11178 30694 11246 30750
rect 11302 30694 11370 30750
rect 11426 30694 11494 30750
rect 11550 30694 11618 30750
rect 11674 30694 11742 30750
rect 11798 30694 11866 30750
rect 11922 30694 11990 30750
rect 12046 30694 12114 30750
rect 12170 30694 12180 30750
rect 10244 30626 12180 30694
rect 10244 30570 10254 30626
rect 10310 30570 10378 30626
rect 10434 30570 10502 30626
rect 10558 30570 10626 30626
rect 10682 30570 10750 30626
rect 10806 30570 10874 30626
rect 10930 30570 10998 30626
rect 11054 30570 11122 30626
rect 11178 30570 11246 30626
rect 11302 30570 11370 30626
rect 11426 30570 11494 30626
rect 11550 30570 11618 30626
rect 11674 30570 11742 30626
rect 11798 30570 11866 30626
rect 11922 30570 11990 30626
rect 12046 30570 12114 30626
rect 12170 30570 12180 30626
rect 10244 30502 12180 30570
rect 10244 30446 10254 30502
rect 10310 30446 10378 30502
rect 10434 30446 10502 30502
rect 10558 30446 10626 30502
rect 10682 30446 10750 30502
rect 10806 30446 10874 30502
rect 10930 30446 10998 30502
rect 11054 30446 11122 30502
rect 11178 30446 11246 30502
rect 11302 30446 11370 30502
rect 11426 30446 11494 30502
rect 11550 30446 11618 30502
rect 11674 30446 11742 30502
rect 11798 30446 11866 30502
rect 11922 30446 11990 30502
rect 12046 30446 12114 30502
rect 12170 30446 12180 30502
rect 10244 30436 12180 30446
rect 12861 33354 14673 33364
rect 12861 33298 12871 33354
rect 12927 33298 12995 33354
rect 13051 33298 13119 33354
rect 13175 33298 13243 33354
rect 13299 33298 13367 33354
rect 13423 33298 13491 33354
rect 13547 33298 13615 33354
rect 13671 33298 13739 33354
rect 13795 33298 13863 33354
rect 13919 33298 13987 33354
rect 14043 33298 14111 33354
rect 14167 33298 14235 33354
rect 14291 33298 14359 33354
rect 14415 33298 14483 33354
rect 14539 33298 14607 33354
rect 14663 33298 14673 33354
rect 12861 33230 14673 33298
rect 12861 33174 12871 33230
rect 12927 33174 12995 33230
rect 13051 33174 13119 33230
rect 13175 33174 13243 33230
rect 13299 33174 13367 33230
rect 13423 33174 13491 33230
rect 13547 33174 13615 33230
rect 13671 33174 13739 33230
rect 13795 33174 13863 33230
rect 13919 33174 13987 33230
rect 14043 33174 14111 33230
rect 14167 33174 14235 33230
rect 14291 33174 14359 33230
rect 14415 33174 14483 33230
rect 14539 33174 14607 33230
rect 14663 33174 14673 33230
rect 12861 33106 14673 33174
rect 12861 33050 12871 33106
rect 12927 33050 12995 33106
rect 13051 33050 13119 33106
rect 13175 33050 13243 33106
rect 13299 33050 13367 33106
rect 13423 33050 13491 33106
rect 13547 33050 13615 33106
rect 13671 33050 13739 33106
rect 13795 33050 13863 33106
rect 13919 33050 13987 33106
rect 14043 33050 14111 33106
rect 14167 33050 14235 33106
rect 14291 33050 14359 33106
rect 14415 33050 14483 33106
rect 14539 33050 14607 33106
rect 14663 33050 14673 33106
rect 12861 32982 14673 33050
rect 12861 32926 12871 32982
rect 12927 32926 12995 32982
rect 13051 32926 13119 32982
rect 13175 32926 13243 32982
rect 13299 32926 13367 32982
rect 13423 32926 13491 32982
rect 13547 32926 13615 32982
rect 13671 32926 13739 32982
rect 13795 32926 13863 32982
rect 13919 32926 13987 32982
rect 14043 32926 14111 32982
rect 14167 32926 14235 32982
rect 14291 32926 14359 32982
rect 14415 32926 14483 32982
rect 14539 32926 14607 32982
rect 14663 32926 14673 32982
rect 12861 32858 14673 32926
rect 12861 32802 12871 32858
rect 12927 32802 12995 32858
rect 13051 32802 13119 32858
rect 13175 32802 13243 32858
rect 13299 32802 13367 32858
rect 13423 32802 13491 32858
rect 13547 32802 13615 32858
rect 13671 32802 13739 32858
rect 13795 32802 13863 32858
rect 13919 32802 13987 32858
rect 14043 32802 14111 32858
rect 14167 32802 14235 32858
rect 14291 32802 14359 32858
rect 14415 32802 14483 32858
rect 14539 32802 14607 32858
rect 14663 32802 14673 32858
rect 12861 32734 14673 32802
rect 12861 32678 12871 32734
rect 12927 32678 12995 32734
rect 13051 32678 13119 32734
rect 13175 32678 13243 32734
rect 13299 32678 13367 32734
rect 13423 32678 13491 32734
rect 13547 32678 13615 32734
rect 13671 32678 13739 32734
rect 13795 32678 13863 32734
rect 13919 32678 13987 32734
rect 14043 32678 14111 32734
rect 14167 32678 14235 32734
rect 14291 32678 14359 32734
rect 14415 32678 14483 32734
rect 14539 32678 14607 32734
rect 14663 32678 14673 32734
rect 12861 32610 14673 32678
rect 12861 32554 12871 32610
rect 12927 32554 12995 32610
rect 13051 32554 13119 32610
rect 13175 32554 13243 32610
rect 13299 32554 13367 32610
rect 13423 32554 13491 32610
rect 13547 32554 13615 32610
rect 13671 32554 13739 32610
rect 13795 32554 13863 32610
rect 13919 32554 13987 32610
rect 14043 32554 14111 32610
rect 14167 32554 14235 32610
rect 14291 32554 14359 32610
rect 14415 32554 14483 32610
rect 14539 32554 14607 32610
rect 14663 32554 14673 32610
rect 12861 32486 14673 32554
rect 12861 32430 12871 32486
rect 12927 32430 12995 32486
rect 13051 32430 13119 32486
rect 13175 32430 13243 32486
rect 13299 32430 13367 32486
rect 13423 32430 13491 32486
rect 13547 32430 13615 32486
rect 13671 32430 13739 32486
rect 13795 32430 13863 32486
rect 13919 32430 13987 32486
rect 14043 32430 14111 32486
rect 14167 32430 14235 32486
rect 14291 32430 14359 32486
rect 14415 32430 14483 32486
rect 14539 32430 14607 32486
rect 14663 32430 14673 32486
rect 12861 32362 14673 32430
rect 12861 32306 12871 32362
rect 12927 32306 12995 32362
rect 13051 32306 13119 32362
rect 13175 32306 13243 32362
rect 13299 32306 13367 32362
rect 13423 32306 13491 32362
rect 13547 32306 13615 32362
rect 13671 32306 13739 32362
rect 13795 32306 13863 32362
rect 13919 32306 13987 32362
rect 14043 32306 14111 32362
rect 14167 32306 14235 32362
rect 14291 32306 14359 32362
rect 14415 32306 14483 32362
rect 14539 32306 14607 32362
rect 14663 32306 14673 32362
rect 12861 32238 14673 32306
rect 12861 32182 12871 32238
rect 12927 32182 12995 32238
rect 13051 32182 13119 32238
rect 13175 32182 13243 32238
rect 13299 32182 13367 32238
rect 13423 32182 13491 32238
rect 13547 32182 13615 32238
rect 13671 32182 13739 32238
rect 13795 32182 13863 32238
rect 13919 32182 13987 32238
rect 14043 32182 14111 32238
rect 14167 32182 14235 32238
rect 14291 32182 14359 32238
rect 14415 32182 14483 32238
rect 14539 32182 14607 32238
rect 14663 32182 14673 32238
rect 12861 32114 14673 32182
rect 12861 32058 12871 32114
rect 12927 32058 12995 32114
rect 13051 32058 13119 32114
rect 13175 32058 13243 32114
rect 13299 32058 13367 32114
rect 13423 32058 13491 32114
rect 13547 32058 13615 32114
rect 13671 32058 13739 32114
rect 13795 32058 13863 32114
rect 13919 32058 13987 32114
rect 14043 32058 14111 32114
rect 14167 32058 14235 32114
rect 14291 32058 14359 32114
rect 14415 32058 14483 32114
rect 14539 32058 14607 32114
rect 14663 32058 14673 32114
rect 12861 31990 14673 32058
rect 12861 31934 12871 31990
rect 12927 31934 12995 31990
rect 13051 31934 13119 31990
rect 13175 31934 13243 31990
rect 13299 31934 13367 31990
rect 13423 31934 13491 31990
rect 13547 31934 13615 31990
rect 13671 31934 13739 31990
rect 13795 31934 13863 31990
rect 13919 31934 13987 31990
rect 14043 31934 14111 31990
rect 14167 31934 14235 31990
rect 14291 31934 14359 31990
rect 14415 31934 14483 31990
rect 14539 31934 14607 31990
rect 14663 31934 14673 31990
rect 12861 31866 14673 31934
rect 12861 31810 12871 31866
rect 12927 31810 12995 31866
rect 13051 31810 13119 31866
rect 13175 31810 13243 31866
rect 13299 31810 13367 31866
rect 13423 31810 13491 31866
rect 13547 31810 13615 31866
rect 13671 31810 13739 31866
rect 13795 31810 13863 31866
rect 13919 31810 13987 31866
rect 14043 31810 14111 31866
rect 14167 31810 14235 31866
rect 14291 31810 14359 31866
rect 14415 31810 14483 31866
rect 14539 31810 14607 31866
rect 14663 31810 14673 31866
rect 12861 31742 14673 31810
rect 12861 31686 12871 31742
rect 12927 31686 12995 31742
rect 13051 31686 13119 31742
rect 13175 31686 13243 31742
rect 13299 31686 13367 31742
rect 13423 31686 13491 31742
rect 13547 31686 13615 31742
rect 13671 31686 13739 31742
rect 13795 31686 13863 31742
rect 13919 31686 13987 31742
rect 14043 31686 14111 31742
rect 14167 31686 14235 31742
rect 14291 31686 14359 31742
rect 14415 31686 14483 31742
rect 14539 31686 14607 31742
rect 14663 31686 14673 31742
rect 12861 31618 14673 31686
rect 12861 31562 12871 31618
rect 12927 31562 12995 31618
rect 13051 31562 13119 31618
rect 13175 31562 13243 31618
rect 13299 31562 13367 31618
rect 13423 31562 13491 31618
rect 13547 31562 13615 31618
rect 13671 31562 13739 31618
rect 13795 31562 13863 31618
rect 13919 31562 13987 31618
rect 14043 31562 14111 31618
rect 14167 31562 14235 31618
rect 14291 31562 14359 31618
rect 14415 31562 14483 31618
rect 14539 31562 14607 31618
rect 14663 31562 14673 31618
rect 12861 31494 14673 31562
rect 12861 31438 12871 31494
rect 12927 31438 12995 31494
rect 13051 31438 13119 31494
rect 13175 31438 13243 31494
rect 13299 31438 13367 31494
rect 13423 31438 13491 31494
rect 13547 31438 13615 31494
rect 13671 31438 13739 31494
rect 13795 31438 13863 31494
rect 13919 31438 13987 31494
rect 14043 31438 14111 31494
rect 14167 31438 14235 31494
rect 14291 31438 14359 31494
rect 14415 31438 14483 31494
rect 14539 31438 14607 31494
rect 14663 31438 14673 31494
rect 12861 31370 14673 31438
rect 12861 31314 12871 31370
rect 12927 31314 12995 31370
rect 13051 31314 13119 31370
rect 13175 31314 13243 31370
rect 13299 31314 13367 31370
rect 13423 31314 13491 31370
rect 13547 31314 13615 31370
rect 13671 31314 13739 31370
rect 13795 31314 13863 31370
rect 13919 31314 13987 31370
rect 14043 31314 14111 31370
rect 14167 31314 14235 31370
rect 14291 31314 14359 31370
rect 14415 31314 14483 31370
rect 14539 31314 14607 31370
rect 14663 31314 14673 31370
rect 12861 31246 14673 31314
rect 12861 31190 12871 31246
rect 12927 31190 12995 31246
rect 13051 31190 13119 31246
rect 13175 31190 13243 31246
rect 13299 31190 13367 31246
rect 13423 31190 13491 31246
rect 13547 31190 13615 31246
rect 13671 31190 13739 31246
rect 13795 31190 13863 31246
rect 13919 31190 13987 31246
rect 14043 31190 14111 31246
rect 14167 31190 14235 31246
rect 14291 31190 14359 31246
rect 14415 31190 14483 31246
rect 14539 31190 14607 31246
rect 14663 31190 14673 31246
rect 12861 31122 14673 31190
rect 12861 31066 12871 31122
rect 12927 31066 12995 31122
rect 13051 31066 13119 31122
rect 13175 31066 13243 31122
rect 13299 31066 13367 31122
rect 13423 31066 13491 31122
rect 13547 31066 13615 31122
rect 13671 31066 13739 31122
rect 13795 31066 13863 31122
rect 13919 31066 13987 31122
rect 14043 31066 14111 31122
rect 14167 31066 14235 31122
rect 14291 31066 14359 31122
rect 14415 31066 14483 31122
rect 14539 31066 14607 31122
rect 14663 31066 14673 31122
rect 12861 30998 14673 31066
rect 12861 30942 12871 30998
rect 12927 30942 12995 30998
rect 13051 30942 13119 30998
rect 13175 30942 13243 30998
rect 13299 30942 13367 30998
rect 13423 30942 13491 30998
rect 13547 30942 13615 30998
rect 13671 30942 13739 30998
rect 13795 30942 13863 30998
rect 13919 30942 13987 30998
rect 14043 30942 14111 30998
rect 14167 30942 14235 30998
rect 14291 30942 14359 30998
rect 14415 30942 14483 30998
rect 14539 30942 14607 30998
rect 14663 30942 14673 30998
rect 12861 30874 14673 30942
rect 12861 30818 12871 30874
rect 12927 30818 12995 30874
rect 13051 30818 13119 30874
rect 13175 30818 13243 30874
rect 13299 30818 13367 30874
rect 13423 30818 13491 30874
rect 13547 30818 13615 30874
rect 13671 30818 13739 30874
rect 13795 30818 13863 30874
rect 13919 30818 13987 30874
rect 14043 30818 14111 30874
rect 14167 30818 14235 30874
rect 14291 30818 14359 30874
rect 14415 30818 14483 30874
rect 14539 30818 14607 30874
rect 14663 30818 14673 30874
rect 12861 30750 14673 30818
rect 12861 30694 12871 30750
rect 12927 30694 12995 30750
rect 13051 30694 13119 30750
rect 13175 30694 13243 30750
rect 13299 30694 13367 30750
rect 13423 30694 13491 30750
rect 13547 30694 13615 30750
rect 13671 30694 13739 30750
rect 13795 30694 13863 30750
rect 13919 30694 13987 30750
rect 14043 30694 14111 30750
rect 14167 30694 14235 30750
rect 14291 30694 14359 30750
rect 14415 30694 14483 30750
rect 14539 30694 14607 30750
rect 14663 30694 14673 30750
rect 12861 30626 14673 30694
rect 12861 30570 12871 30626
rect 12927 30570 12995 30626
rect 13051 30570 13119 30626
rect 13175 30570 13243 30626
rect 13299 30570 13367 30626
rect 13423 30570 13491 30626
rect 13547 30570 13615 30626
rect 13671 30570 13739 30626
rect 13795 30570 13863 30626
rect 13919 30570 13987 30626
rect 14043 30570 14111 30626
rect 14167 30570 14235 30626
rect 14291 30570 14359 30626
rect 14415 30570 14483 30626
rect 14539 30570 14607 30626
rect 14663 30570 14673 30626
rect 12861 30502 14673 30570
rect 12861 30446 12871 30502
rect 12927 30446 12995 30502
rect 13051 30446 13119 30502
rect 13175 30446 13243 30502
rect 13299 30446 13367 30502
rect 13423 30446 13491 30502
rect 13547 30446 13615 30502
rect 13671 30446 13739 30502
rect 13795 30446 13863 30502
rect 13919 30446 13987 30502
rect 14043 30446 14111 30502
rect 14167 30446 14235 30502
rect 14291 30446 14359 30502
rect 14415 30446 14483 30502
rect 14539 30446 14607 30502
rect 14663 30446 14673 30502
rect 12861 30436 14673 30446
rect 305 30148 2117 30158
rect 305 30092 315 30148
rect 371 30092 439 30148
rect 495 30092 563 30148
rect 619 30092 687 30148
rect 743 30092 811 30148
rect 867 30092 935 30148
rect 991 30092 1059 30148
rect 1115 30092 1183 30148
rect 1239 30092 1307 30148
rect 1363 30092 1431 30148
rect 1487 30092 1555 30148
rect 1611 30092 1679 30148
rect 1735 30092 1803 30148
rect 1859 30092 1927 30148
rect 1983 30092 2051 30148
rect 2107 30092 2117 30148
rect 305 30024 2117 30092
rect 305 29968 315 30024
rect 371 29968 439 30024
rect 495 29968 563 30024
rect 619 29968 687 30024
rect 743 29968 811 30024
rect 867 29968 935 30024
rect 991 29968 1059 30024
rect 1115 29968 1183 30024
rect 1239 29968 1307 30024
rect 1363 29968 1431 30024
rect 1487 29968 1555 30024
rect 1611 29968 1679 30024
rect 1735 29968 1803 30024
rect 1859 29968 1927 30024
rect 1983 29968 2051 30024
rect 2107 29968 2117 30024
rect 305 29900 2117 29968
rect 305 29844 315 29900
rect 371 29844 439 29900
rect 495 29844 563 29900
rect 619 29844 687 29900
rect 743 29844 811 29900
rect 867 29844 935 29900
rect 991 29844 1059 29900
rect 1115 29844 1183 29900
rect 1239 29844 1307 29900
rect 1363 29844 1431 29900
rect 1487 29844 1555 29900
rect 1611 29844 1679 29900
rect 1735 29844 1803 29900
rect 1859 29844 1927 29900
rect 1983 29844 2051 29900
rect 2107 29844 2117 29900
rect 305 29776 2117 29844
rect 305 29720 315 29776
rect 371 29720 439 29776
rect 495 29720 563 29776
rect 619 29720 687 29776
rect 743 29720 811 29776
rect 867 29720 935 29776
rect 991 29720 1059 29776
rect 1115 29720 1183 29776
rect 1239 29720 1307 29776
rect 1363 29720 1431 29776
rect 1487 29720 1555 29776
rect 1611 29720 1679 29776
rect 1735 29720 1803 29776
rect 1859 29720 1927 29776
rect 1983 29720 2051 29776
rect 2107 29720 2117 29776
rect 305 29652 2117 29720
rect 305 29596 315 29652
rect 371 29596 439 29652
rect 495 29596 563 29652
rect 619 29596 687 29652
rect 743 29596 811 29652
rect 867 29596 935 29652
rect 991 29596 1059 29652
rect 1115 29596 1183 29652
rect 1239 29596 1307 29652
rect 1363 29596 1431 29652
rect 1487 29596 1555 29652
rect 1611 29596 1679 29652
rect 1735 29596 1803 29652
rect 1859 29596 1927 29652
rect 1983 29596 2051 29652
rect 2107 29596 2117 29652
rect 305 29528 2117 29596
rect 305 29472 315 29528
rect 371 29472 439 29528
rect 495 29472 563 29528
rect 619 29472 687 29528
rect 743 29472 811 29528
rect 867 29472 935 29528
rect 991 29472 1059 29528
rect 1115 29472 1183 29528
rect 1239 29472 1307 29528
rect 1363 29472 1431 29528
rect 1487 29472 1555 29528
rect 1611 29472 1679 29528
rect 1735 29472 1803 29528
rect 1859 29472 1927 29528
rect 1983 29472 2051 29528
rect 2107 29472 2117 29528
rect 305 29404 2117 29472
rect 305 29348 315 29404
rect 371 29348 439 29404
rect 495 29348 563 29404
rect 619 29348 687 29404
rect 743 29348 811 29404
rect 867 29348 935 29404
rect 991 29348 1059 29404
rect 1115 29348 1183 29404
rect 1239 29348 1307 29404
rect 1363 29348 1431 29404
rect 1487 29348 1555 29404
rect 1611 29348 1679 29404
rect 1735 29348 1803 29404
rect 1859 29348 1927 29404
rect 1983 29348 2051 29404
rect 2107 29348 2117 29404
rect 305 29280 2117 29348
rect 305 29224 315 29280
rect 371 29224 439 29280
rect 495 29224 563 29280
rect 619 29224 687 29280
rect 743 29224 811 29280
rect 867 29224 935 29280
rect 991 29224 1059 29280
rect 1115 29224 1183 29280
rect 1239 29224 1307 29280
rect 1363 29224 1431 29280
rect 1487 29224 1555 29280
rect 1611 29224 1679 29280
rect 1735 29224 1803 29280
rect 1859 29224 1927 29280
rect 1983 29224 2051 29280
rect 2107 29224 2117 29280
rect 305 29156 2117 29224
rect 305 29100 315 29156
rect 371 29100 439 29156
rect 495 29100 563 29156
rect 619 29100 687 29156
rect 743 29100 811 29156
rect 867 29100 935 29156
rect 991 29100 1059 29156
rect 1115 29100 1183 29156
rect 1239 29100 1307 29156
rect 1363 29100 1431 29156
rect 1487 29100 1555 29156
rect 1611 29100 1679 29156
rect 1735 29100 1803 29156
rect 1859 29100 1927 29156
rect 1983 29100 2051 29156
rect 2107 29100 2117 29156
rect 305 29032 2117 29100
rect 305 28976 315 29032
rect 371 28976 439 29032
rect 495 28976 563 29032
rect 619 28976 687 29032
rect 743 28976 811 29032
rect 867 28976 935 29032
rect 991 28976 1059 29032
rect 1115 28976 1183 29032
rect 1239 28976 1307 29032
rect 1363 28976 1431 29032
rect 1487 28976 1555 29032
rect 1611 28976 1679 29032
rect 1735 28976 1803 29032
rect 1859 28976 1927 29032
rect 1983 28976 2051 29032
rect 2107 28976 2117 29032
rect 305 28908 2117 28976
rect 305 28852 315 28908
rect 371 28852 439 28908
rect 495 28852 563 28908
rect 619 28852 687 28908
rect 743 28852 811 28908
rect 867 28852 935 28908
rect 991 28852 1059 28908
rect 1115 28852 1183 28908
rect 1239 28852 1307 28908
rect 1363 28852 1431 28908
rect 1487 28852 1555 28908
rect 1611 28852 1679 28908
rect 1735 28852 1803 28908
rect 1859 28852 1927 28908
rect 1983 28852 2051 28908
rect 2107 28852 2117 28908
rect 305 28842 2117 28852
rect 2798 30148 4734 30158
rect 2798 30092 2808 30148
rect 2864 30092 2932 30148
rect 2988 30092 3056 30148
rect 3112 30092 3180 30148
rect 3236 30092 3304 30148
rect 3360 30092 3428 30148
rect 3484 30092 3552 30148
rect 3608 30092 3676 30148
rect 3732 30092 3800 30148
rect 3856 30092 3924 30148
rect 3980 30092 4048 30148
rect 4104 30092 4172 30148
rect 4228 30092 4296 30148
rect 4352 30092 4420 30148
rect 4476 30092 4544 30148
rect 4600 30092 4668 30148
rect 4724 30092 4734 30148
rect 2798 30024 4734 30092
rect 2798 29968 2808 30024
rect 2864 29968 2932 30024
rect 2988 29968 3056 30024
rect 3112 29968 3180 30024
rect 3236 29968 3304 30024
rect 3360 29968 3428 30024
rect 3484 29968 3552 30024
rect 3608 29968 3676 30024
rect 3732 29968 3800 30024
rect 3856 29968 3924 30024
rect 3980 29968 4048 30024
rect 4104 29968 4172 30024
rect 4228 29968 4296 30024
rect 4352 29968 4420 30024
rect 4476 29968 4544 30024
rect 4600 29968 4668 30024
rect 4724 29968 4734 30024
rect 2798 29900 4734 29968
rect 2798 29844 2808 29900
rect 2864 29844 2932 29900
rect 2988 29844 3056 29900
rect 3112 29844 3180 29900
rect 3236 29844 3304 29900
rect 3360 29844 3428 29900
rect 3484 29844 3552 29900
rect 3608 29844 3676 29900
rect 3732 29844 3800 29900
rect 3856 29844 3924 29900
rect 3980 29844 4048 29900
rect 4104 29844 4172 29900
rect 4228 29844 4296 29900
rect 4352 29844 4420 29900
rect 4476 29844 4544 29900
rect 4600 29844 4668 29900
rect 4724 29844 4734 29900
rect 2798 29776 4734 29844
rect 2798 29720 2808 29776
rect 2864 29720 2932 29776
rect 2988 29720 3056 29776
rect 3112 29720 3180 29776
rect 3236 29720 3304 29776
rect 3360 29720 3428 29776
rect 3484 29720 3552 29776
rect 3608 29720 3676 29776
rect 3732 29720 3800 29776
rect 3856 29720 3924 29776
rect 3980 29720 4048 29776
rect 4104 29720 4172 29776
rect 4228 29720 4296 29776
rect 4352 29720 4420 29776
rect 4476 29720 4544 29776
rect 4600 29720 4668 29776
rect 4724 29720 4734 29776
rect 2798 29652 4734 29720
rect 2798 29596 2808 29652
rect 2864 29596 2932 29652
rect 2988 29596 3056 29652
rect 3112 29596 3180 29652
rect 3236 29596 3304 29652
rect 3360 29596 3428 29652
rect 3484 29596 3552 29652
rect 3608 29596 3676 29652
rect 3732 29596 3800 29652
rect 3856 29596 3924 29652
rect 3980 29596 4048 29652
rect 4104 29596 4172 29652
rect 4228 29596 4296 29652
rect 4352 29596 4420 29652
rect 4476 29596 4544 29652
rect 4600 29596 4668 29652
rect 4724 29596 4734 29652
rect 2798 29528 4734 29596
rect 2798 29472 2808 29528
rect 2864 29472 2932 29528
rect 2988 29472 3056 29528
rect 3112 29472 3180 29528
rect 3236 29472 3304 29528
rect 3360 29472 3428 29528
rect 3484 29472 3552 29528
rect 3608 29472 3676 29528
rect 3732 29472 3800 29528
rect 3856 29472 3924 29528
rect 3980 29472 4048 29528
rect 4104 29472 4172 29528
rect 4228 29472 4296 29528
rect 4352 29472 4420 29528
rect 4476 29472 4544 29528
rect 4600 29472 4668 29528
rect 4724 29472 4734 29528
rect 2798 29404 4734 29472
rect 2798 29348 2808 29404
rect 2864 29348 2932 29404
rect 2988 29348 3056 29404
rect 3112 29348 3180 29404
rect 3236 29348 3304 29404
rect 3360 29348 3428 29404
rect 3484 29348 3552 29404
rect 3608 29348 3676 29404
rect 3732 29348 3800 29404
rect 3856 29348 3924 29404
rect 3980 29348 4048 29404
rect 4104 29348 4172 29404
rect 4228 29348 4296 29404
rect 4352 29348 4420 29404
rect 4476 29348 4544 29404
rect 4600 29348 4668 29404
rect 4724 29348 4734 29404
rect 2798 29280 4734 29348
rect 2798 29224 2808 29280
rect 2864 29224 2932 29280
rect 2988 29224 3056 29280
rect 3112 29224 3180 29280
rect 3236 29224 3304 29280
rect 3360 29224 3428 29280
rect 3484 29224 3552 29280
rect 3608 29224 3676 29280
rect 3732 29224 3800 29280
rect 3856 29224 3924 29280
rect 3980 29224 4048 29280
rect 4104 29224 4172 29280
rect 4228 29224 4296 29280
rect 4352 29224 4420 29280
rect 4476 29224 4544 29280
rect 4600 29224 4668 29280
rect 4724 29224 4734 29280
rect 2798 29156 4734 29224
rect 2798 29100 2808 29156
rect 2864 29100 2932 29156
rect 2988 29100 3056 29156
rect 3112 29100 3180 29156
rect 3236 29100 3304 29156
rect 3360 29100 3428 29156
rect 3484 29100 3552 29156
rect 3608 29100 3676 29156
rect 3732 29100 3800 29156
rect 3856 29100 3924 29156
rect 3980 29100 4048 29156
rect 4104 29100 4172 29156
rect 4228 29100 4296 29156
rect 4352 29100 4420 29156
rect 4476 29100 4544 29156
rect 4600 29100 4668 29156
rect 4724 29100 4734 29156
rect 2798 29032 4734 29100
rect 2798 28976 2808 29032
rect 2864 28976 2932 29032
rect 2988 28976 3056 29032
rect 3112 28976 3180 29032
rect 3236 28976 3304 29032
rect 3360 28976 3428 29032
rect 3484 28976 3552 29032
rect 3608 28976 3676 29032
rect 3732 28976 3800 29032
rect 3856 28976 3924 29032
rect 3980 28976 4048 29032
rect 4104 28976 4172 29032
rect 4228 28976 4296 29032
rect 4352 28976 4420 29032
rect 4476 28976 4544 29032
rect 4600 28976 4668 29032
rect 4724 28976 4734 29032
rect 2798 28908 4734 28976
rect 2798 28852 2808 28908
rect 2864 28852 2932 28908
rect 2988 28852 3056 28908
rect 3112 28852 3180 28908
rect 3236 28852 3304 28908
rect 3360 28852 3428 28908
rect 3484 28852 3552 28908
rect 3608 28852 3676 28908
rect 3732 28852 3800 28908
rect 3856 28852 3924 28908
rect 3980 28852 4048 28908
rect 4104 28852 4172 28908
rect 4228 28852 4296 28908
rect 4352 28852 4420 28908
rect 4476 28852 4544 28908
rect 4600 28852 4668 28908
rect 4724 28852 4734 28908
rect 2798 28842 4734 28852
rect 5168 30148 7104 30158
rect 5168 30092 5178 30148
rect 5234 30092 5302 30148
rect 5358 30092 5426 30148
rect 5482 30092 5550 30148
rect 5606 30092 5674 30148
rect 5730 30092 5798 30148
rect 5854 30092 5922 30148
rect 5978 30092 6046 30148
rect 6102 30092 6170 30148
rect 6226 30092 6294 30148
rect 6350 30092 6418 30148
rect 6474 30092 6542 30148
rect 6598 30092 6666 30148
rect 6722 30092 6790 30148
rect 6846 30092 6914 30148
rect 6970 30092 7038 30148
rect 7094 30092 7104 30148
rect 5168 30024 7104 30092
rect 5168 29968 5178 30024
rect 5234 29968 5302 30024
rect 5358 29968 5426 30024
rect 5482 29968 5550 30024
rect 5606 29968 5674 30024
rect 5730 29968 5798 30024
rect 5854 29968 5922 30024
rect 5978 29968 6046 30024
rect 6102 29968 6170 30024
rect 6226 29968 6294 30024
rect 6350 29968 6418 30024
rect 6474 29968 6542 30024
rect 6598 29968 6666 30024
rect 6722 29968 6790 30024
rect 6846 29968 6914 30024
rect 6970 29968 7038 30024
rect 7094 29968 7104 30024
rect 5168 29900 7104 29968
rect 5168 29844 5178 29900
rect 5234 29844 5302 29900
rect 5358 29844 5426 29900
rect 5482 29844 5550 29900
rect 5606 29844 5674 29900
rect 5730 29844 5798 29900
rect 5854 29844 5922 29900
rect 5978 29844 6046 29900
rect 6102 29844 6170 29900
rect 6226 29844 6294 29900
rect 6350 29844 6418 29900
rect 6474 29844 6542 29900
rect 6598 29844 6666 29900
rect 6722 29844 6790 29900
rect 6846 29844 6914 29900
rect 6970 29844 7038 29900
rect 7094 29844 7104 29900
rect 5168 29776 7104 29844
rect 5168 29720 5178 29776
rect 5234 29720 5302 29776
rect 5358 29720 5426 29776
rect 5482 29720 5550 29776
rect 5606 29720 5674 29776
rect 5730 29720 5798 29776
rect 5854 29720 5922 29776
rect 5978 29720 6046 29776
rect 6102 29720 6170 29776
rect 6226 29720 6294 29776
rect 6350 29720 6418 29776
rect 6474 29720 6542 29776
rect 6598 29720 6666 29776
rect 6722 29720 6790 29776
rect 6846 29720 6914 29776
rect 6970 29720 7038 29776
rect 7094 29720 7104 29776
rect 5168 29652 7104 29720
rect 5168 29596 5178 29652
rect 5234 29596 5302 29652
rect 5358 29596 5426 29652
rect 5482 29596 5550 29652
rect 5606 29596 5674 29652
rect 5730 29596 5798 29652
rect 5854 29596 5922 29652
rect 5978 29596 6046 29652
rect 6102 29596 6170 29652
rect 6226 29596 6294 29652
rect 6350 29596 6418 29652
rect 6474 29596 6542 29652
rect 6598 29596 6666 29652
rect 6722 29596 6790 29652
rect 6846 29596 6914 29652
rect 6970 29596 7038 29652
rect 7094 29596 7104 29652
rect 5168 29528 7104 29596
rect 5168 29472 5178 29528
rect 5234 29472 5302 29528
rect 5358 29472 5426 29528
rect 5482 29472 5550 29528
rect 5606 29472 5674 29528
rect 5730 29472 5798 29528
rect 5854 29472 5922 29528
rect 5978 29472 6046 29528
rect 6102 29472 6170 29528
rect 6226 29472 6294 29528
rect 6350 29472 6418 29528
rect 6474 29472 6542 29528
rect 6598 29472 6666 29528
rect 6722 29472 6790 29528
rect 6846 29472 6914 29528
rect 6970 29472 7038 29528
rect 7094 29472 7104 29528
rect 5168 29404 7104 29472
rect 5168 29348 5178 29404
rect 5234 29348 5302 29404
rect 5358 29348 5426 29404
rect 5482 29348 5550 29404
rect 5606 29348 5674 29404
rect 5730 29348 5798 29404
rect 5854 29348 5922 29404
rect 5978 29348 6046 29404
rect 6102 29348 6170 29404
rect 6226 29348 6294 29404
rect 6350 29348 6418 29404
rect 6474 29348 6542 29404
rect 6598 29348 6666 29404
rect 6722 29348 6790 29404
rect 6846 29348 6914 29404
rect 6970 29348 7038 29404
rect 7094 29348 7104 29404
rect 5168 29280 7104 29348
rect 5168 29224 5178 29280
rect 5234 29224 5302 29280
rect 5358 29224 5426 29280
rect 5482 29224 5550 29280
rect 5606 29224 5674 29280
rect 5730 29224 5798 29280
rect 5854 29224 5922 29280
rect 5978 29224 6046 29280
rect 6102 29224 6170 29280
rect 6226 29224 6294 29280
rect 6350 29224 6418 29280
rect 6474 29224 6542 29280
rect 6598 29224 6666 29280
rect 6722 29224 6790 29280
rect 6846 29224 6914 29280
rect 6970 29224 7038 29280
rect 7094 29224 7104 29280
rect 5168 29156 7104 29224
rect 5168 29100 5178 29156
rect 5234 29100 5302 29156
rect 5358 29100 5426 29156
rect 5482 29100 5550 29156
rect 5606 29100 5674 29156
rect 5730 29100 5798 29156
rect 5854 29100 5922 29156
rect 5978 29100 6046 29156
rect 6102 29100 6170 29156
rect 6226 29100 6294 29156
rect 6350 29100 6418 29156
rect 6474 29100 6542 29156
rect 6598 29100 6666 29156
rect 6722 29100 6790 29156
rect 6846 29100 6914 29156
rect 6970 29100 7038 29156
rect 7094 29100 7104 29156
rect 5168 29032 7104 29100
rect 5168 28976 5178 29032
rect 5234 28976 5302 29032
rect 5358 28976 5426 29032
rect 5482 28976 5550 29032
rect 5606 28976 5674 29032
rect 5730 28976 5798 29032
rect 5854 28976 5922 29032
rect 5978 28976 6046 29032
rect 6102 28976 6170 29032
rect 6226 28976 6294 29032
rect 6350 28976 6418 29032
rect 6474 28976 6542 29032
rect 6598 28976 6666 29032
rect 6722 28976 6790 29032
rect 6846 28976 6914 29032
rect 6970 28976 7038 29032
rect 7094 28976 7104 29032
rect 5168 28908 7104 28976
rect 5168 28852 5178 28908
rect 5234 28852 5302 28908
rect 5358 28852 5426 28908
rect 5482 28852 5550 28908
rect 5606 28852 5674 28908
rect 5730 28852 5798 28908
rect 5854 28852 5922 28908
rect 5978 28852 6046 28908
rect 6102 28852 6170 28908
rect 6226 28852 6294 28908
rect 6350 28852 6418 28908
rect 6474 28852 6542 28908
rect 6598 28852 6666 28908
rect 6722 28852 6790 28908
rect 6846 28852 6914 28908
rect 6970 28852 7038 28908
rect 7094 28852 7104 28908
rect 5168 28842 7104 28852
rect 7874 30148 9810 30158
rect 7874 30092 7884 30148
rect 7940 30092 8008 30148
rect 8064 30092 8132 30148
rect 8188 30092 8256 30148
rect 8312 30092 8380 30148
rect 8436 30092 8504 30148
rect 8560 30092 8628 30148
rect 8684 30092 8752 30148
rect 8808 30092 8876 30148
rect 8932 30092 9000 30148
rect 9056 30092 9124 30148
rect 9180 30092 9248 30148
rect 9304 30092 9372 30148
rect 9428 30092 9496 30148
rect 9552 30092 9620 30148
rect 9676 30092 9744 30148
rect 9800 30092 9810 30148
rect 7874 30024 9810 30092
rect 7874 29968 7884 30024
rect 7940 29968 8008 30024
rect 8064 29968 8132 30024
rect 8188 29968 8256 30024
rect 8312 29968 8380 30024
rect 8436 29968 8504 30024
rect 8560 29968 8628 30024
rect 8684 29968 8752 30024
rect 8808 29968 8876 30024
rect 8932 29968 9000 30024
rect 9056 29968 9124 30024
rect 9180 29968 9248 30024
rect 9304 29968 9372 30024
rect 9428 29968 9496 30024
rect 9552 29968 9620 30024
rect 9676 29968 9744 30024
rect 9800 29968 9810 30024
rect 7874 29900 9810 29968
rect 7874 29844 7884 29900
rect 7940 29844 8008 29900
rect 8064 29844 8132 29900
rect 8188 29844 8256 29900
rect 8312 29844 8380 29900
rect 8436 29844 8504 29900
rect 8560 29844 8628 29900
rect 8684 29844 8752 29900
rect 8808 29844 8876 29900
rect 8932 29844 9000 29900
rect 9056 29844 9124 29900
rect 9180 29844 9248 29900
rect 9304 29844 9372 29900
rect 9428 29844 9496 29900
rect 9552 29844 9620 29900
rect 9676 29844 9744 29900
rect 9800 29844 9810 29900
rect 7874 29776 9810 29844
rect 7874 29720 7884 29776
rect 7940 29720 8008 29776
rect 8064 29720 8132 29776
rect 8188 29720 8256 29776
rect 8312 29720 8380 29776
rect 8436 29720 8504 29776
rect 8560 29720 8628 29776
rect 8684 29720 8752 29776
rect 8808 29720 8876 29776
rect 8932 29720 9000 29776
rect 9056 29720 9124 29776
rect 9180 29720 9248 29776
rect 9304 29720 9372 29776
rect 9428 29720 9496 29776
rect 9552 29720 9620 29776
rect 9676 29720 9744 29776
rect 9800 29720 9810 29776
rect 7874 29652 9810 29720
rect 7874 29596 7884 29652
rect 7940 29596 8008 29652
rect 8064 29596 8132 29652
rect 8188 29596 8256 29652
rect 8312 29596 8380 29652
rect 8436 29596 8504 29652
rect 8560 29596 8628 29652
rect 8684 29596 8752 29652
rect 8808 29596 8876 29652
rect 8932 29596 9000 29652
rect 9056 29596 9124 29652
rect 9180 29596 9248 29652
rect 9304 29596 9372 29652
rect 9428 29596 9496 29652
rect 9552 29596 9620 29652
rect 9676 29596 9744 29652
rect 9800 29596 9810 29652
rect 7874 29528 9810 29596
rect 7874 29472 7884 29528
rect 7940 29472 8008 29528
rect 8064 29472 8132 29528
rect 8188 29472 8256 29528
rect 8312 29472 8380 29528
rect 8436 29472 8504 29528
rect 8560 29472 8628 29528
rect 8684 29472 8752 29528
rect 8808 29472 8876 29528
rect 8932 29472 9000 29528
rect 9056 29472 9124 29528
rect 9180 29472 9248 29528
rect 9304 29472 9372 29528
rect 9428 29472 9496 29528
rect 9552 29472 9620 29528
rect 9676 29472 9744 29528
rect 9800 29472 9810 29528
rect 7874 29404 9810 29472
rect 7874 29348 7884 29404
rect 7940 29348 8008 29404
rect 8064 29348 8132 29404
rect 8188 29348 8256 29404
rect 8312 29348 8380 29404
rect 8436 29348 8504 29404
rect 8560 29348 8628 29404
rect 8684 29348 8752 29404
rect 8808 29348 8876 29404
rect 8932 29348 9000 29404
rect 9056 29348 9124 29404
rect 9180 29348 9248 29404
rect 9304 29348 9372 29404
rect 9428 29348 9496 29404
rect 9552 29348 9620 29404
rect 9676 29348 9744 29404
rect 9800 29348 9810 29404
rect 7874 29280 9810 29348
rect 7874 29224 7884 29280
rect 7940 29224 8008 29280
rect 8064 29224 8132 29280
rect 8188 29224 8256 29280
rect 8312 29224 8380 29280
rect 8436 29224 8504 29280
rect 8560 29224 8628 29280
rect 8684 29224 8752 29280
rect 8808 29224 8876 29280
rect 8932 29224 9000 29280
rect 9056 29224 9124 29280
rect 9180 29224 9248 29280
rect 9304 29224 9372 29280
rect 9428 29224 9496 29280
rect 9552 29224 9620 29280
rect 9676 29224 9744 29280
rect 9800 29224 9810 29280
rect 7874 29156 9810 29224
rect 7874 29100 7884 29156
rect 7940 29100 8008 29156
rect 8064 29100 8132 29156
rect 8188 29100 8256 29156
rect 8312 29100 8380 29156
rect 8436 29100 8504 29156
rect 8560 29100 8628 29156
rect 8684 29100 8752 29156
rect 8808 29100 8876 29156
rect 8932 29100 9000 29156
rect 9056 29100 9124 29156
rect 9180 29100 9248 29156
rect 9304 29100 9372 29156
rect 9428 29100 9496 29156
rect 9552 29100 9620 29156
rect 9676 29100 9744 29156
rect 9800 29100 9810 29156
rect 7874 29032 9810 29100
rect 7874 28976 7884 29032
rect 7940 28976 8008 29032
rect 8064 28976 8132 29032
rect 8188 28976 8256 29032
rect 8312 28976 8380 29032
rect 8436 28976 8504 29032
rect 8560 28976 8628 29032
rect 8684 28976 8752 29032
rect 8808 28976 8876 29032
rect 8932 28976 9000 29032
rect 9056 28976 9124 29032
rect 9180 28976 9248 29032
rect 9304 28976 9372 29032
rect 9428 28976 9496 29032
rect 9552 28976 9620 29032
rect 9676 28976 9744 29032
rect 9800 28976 9810 29032
rect 7874 28908 9810 28976
rect 7874 28852 7884 28908
rect 7940 28852 8008 28908
rect 8064 28852 8132 28908
rect 8188 28852 8256 28908
rect 8312 28852 8380 28908
rect 8436 28852 8504 28908
rect 8560 28852 8628 28908
rect 8684 28852 8752 28908
rect 8808 28852 8876 28908
rect 8932 28852 9000 28908
rect 9056 28852 9124 28908
rect 9180 28852 9248 28908
rect 9304 28852 9372 28908
rect 9428 28852 9496 28908
rect 9552 28852 9620 28908
rect 9676 28852 9744 28908
rect 9800 28852 9810 28908
rect 7874 28842 9810 28852
rect 10244 30148 12180 30158
rect 10244 30092 10254 30148
rect 10310 30092 10378 30148
rect 10434 30092 10502 30148
rect 10558 30092 10626 30148
rect 10682 30092 10750 30148
rect 10806 30092 10874 30148
rect 10930 30092 10998 30148
rect 11054 30092 11122 30148
rect 11178 30092 11246 30148
rect 11302 30092 11370 30148
rect 11426 30092 11494 30148
rect 11550 30092 11618 30148
rect 11674 30092 11742 30148
rect 11798 30092 11866 30148
rect 11922 30092 11990 30148
rect 12046 30092 12114 30148
rect 12170 30092 12180 30148
rect 10244 30024 12180 30092
rect 10244 29968 10254 30024
rect 10310 29968 10378 30024
rect 10434 29968 10502 30024
rect 10558 29968 10626 30024
rect 10682 29968 10750 30024
rect 10806 29968 10874 30024
rect 10930 29968 10998 30024
rect 11054 29968 11122 30024
rect 11178 29968 11246 30024
rect 11302 29968 11370 30024
rect 11426 29968 11494 30024
rect 11550 29968 11618 30024
rect 11674 29968 11742 30024
rect 11798 29968 11866 30024
rect 11922 29968 11990 30024
rect 12046 29968 12114 30024
rect 12170 29968 12180 30024
rect 10244 29900 12180 29968
rect 10244 29844 10254 29900
rect 10310 29844 10378 29900
rect 10434 29844 10502 29900
rect 10558 29844 10626 29900
rect 10682 29844 10750 29900
rect 10806 29844 10874 29900
rect 10930 29844 10998 29900
rect 11054 29844 11122 29900
rect 11178 29844 11246 29900
rect 11302 29844 11370 29900
rect 11426 29844 11494 29900
rect 11550 29844 11618 29900
rect 11674 29844 11742 29900
rect 11798 29844 11866 29900
rect 11922 29844 11990 29900
rect 12046 29844 12114 29900
rect 12170 29844 12180 29900
rect 10244 29776 12180 29844
rect 10244 29720 10254 29776
rect 10310 29720 10378 29776
rect 10434 29720 10502 29776
rect 10558 29720 10626 29776
rect 10682 29720 10750 29776
rect 10806 29720 10874 29776
rect 10930 29720 10998 29776
rect 11054 29720 11122 29776
rect 11178 29720 11246 29776
rect 11302 29720 11370 29776
rect 11426 29720 11494 29776
rect 11550 29720 11618 29776
rect 11674 29720 11742 29776
rect 11798 29720 11866 29776
rect 11922 29720 11990 29776
rect 12046 29720 12114 29776
rect 12170 29720 12180 29776
rect 10244 29652 12180 29720
rect 10244 29596 10254 29652
rect 10310 29596 10378 29652
rect 10434 29596 10502 29652
rect 10558 29596 10626 29652
rect 10682 29596 10750 29652
rect 10806 29596 10874 29652
rect 10930 29596 10998 29652
rect 11054 29596 11122 29652
rect 11178 29596 11246 29652
rect 11302 29596 11370 29652
rect 11426 29596 11494 29652
rect 11550 29596 11618 29652
rect 11674 29596 11742 29652
rect 11798 29596 11866 29652
rect 11922 29596 11990 29652
rect 12046 29596 12114 29652
rect 12170 29596 12180 29652
rect 10244 29528 12180 29596
rect 10244 29472 10254 29528
rect 10310 29472 10378 29528
rect 10434 29472 10502 29528
rect 10558 29472 10626 29528
rect 10682 29472 10750 29528
rect 10806 29472 10874 29528
rect 10930 29472 10998 29528
rect 11054 29472 11122 29528
rect 11178 29472 11246 29528
rect 11302 29472 11370 29528
rect 11426 29472 11494 29528
rect 11550 29472 11618 29528
rect 11674 29472 11742 29528
rect 11798 29472 11866 29528
rect 11922 29472 11990 29528
rect 12046 29472 12114 29528
rect 12170 29472 12180 29528
rect 10244 29404 12180 29472
rect 10244 29348 10254 29404
rect 10310 29348 10378 29404
rect 10434 29348 10502 29404
rect 10558 29348 10626 29404
rect 10682 29348 10750 29404
rect 10806 29348 10874 29404
rect 10930 29348 10998 29404
rect 11054 29348 11122 29404
rect 11178 29348 11246 29404
rect 11302 29348 11370 29404
rect 11426 29348 11494 29404
rect 11550 29348 11618 29404
rect 11674 29348 11742 29404
rect 11798 29348 11866 29404
rect 11922 29348 11990 29404
rect 12046 29348 12114 29404
rect 12170 29348 12180 29404
rect 10244 29280 12180 29348
rect 10244 29224 10254 29280
rect 10310 29224 10378 29280
rect 10434 29224 10502 29280
rect 10558 29224 10626 29280
rect 10682 29224 10750 29280
rect 10806 29224 10874 29280
rect 10930 29224 10998 29280
rect 11054 29224 11122 29280
rect 11178 29224 11246 29280
rect 11302 29224 11370 29280
rect 11426 29224 11494 29280
rect 11550 29224 11618 29280
rect 11674 29224 11742 29280
rect 11798 29224 11866 29280
rect 11922 29224 11990 29280
rect 12046 29224 12114 29280
rect 12170 29224 12180 29280
rect 10244 29156 12180 29224
rect 10244 29100 10254 29156
rect 10310 29100 10378 29156
rect 10434 29100 10502 29156
rect 10558 29100 10626 29156
rect 10682 29100 10750 29156
rect 10806 29100 10874 29156
rect 10930 29100 10998 29156
rect 11054 29100 11122 29156
rect 11178 29100 11246 29156
rect 11302 29100 11370 29156
rect 11426 29100 11494 29156
rect 11550 29100 11618 29156
rect 11674 29100 11742 29156
rect 11798 29100 11866 29156
rect 11922 29100 11990 29156
rect 12046 29100 12114 29156
rect 12170 29100 12180 29156
rect 10244 29032 12180 29100
rect 10244 28976 10254 29032
rect 10310 28976 10378 29032
rect 10434 28976 10502 29032
rect 10558 28976 10626 29032
rect 10682 28976 10750 29032
rect 10806 28976 10874 29032
rect 10930 28976 10998 29032
rect 11054 28976 11122 29032
rect 11178 28976 11246 29032
rect 11302 28976 11370 29032
rect 11426 28976 11494 29032
rect 11550 28976 11618 29032
rect 11674 28976 11742 29032
rect 11798 28976 11866 29032
rect 11922 28976 11990 29032
rect 12046 28976 12114 29032
rect 12170 28976 12180 29032
rect 10244 28908 12180 28976
rect 10244 28852 10254 28908
rect 10310 28852 10378 28908
rect 10434 28852 10502 28908
rect 10558 28852 10626 28908
rect 10682 28852 10750 28908
rect 10806 28852 10874 28908
rect 10930 28852 10998 28908
rect 11054 28852 11122 28908
rect 11178 28852 11246 28908
rect 11302 28852 11370 28908
rect 11426 28852 11494 28908
rect 11550 28852 11618 28908
rect 11674 28852 11742 28908
rect 11798 28852 11866 28908
rect 11922 28852 11990 28908
rect 12046 28852 12114 28908
rect 12170 28852 12180 28908
rect 10244 28842 12180 28852
rect 12861 30148 14673 30158
rect 12861 30092 12871 30148
rect 12927 30092 12995 30148
rect 13051 30092 13119 30148
rect 13175 30092 13243 30148
rect 13299 30092 13367 30148
rect 13423 30092 13491 30148
rect 13547 30092 13615 30148
rect 13671 30092 13739 30148
rect 13795 30092 13863 30148
rect 13919 30092 13987 30148
rect 14043 30092 14111 30148
rect 14167 30092 14235 30148
rect 14291 30092 14359 30148
rect 14415 30092 14483 30148
rect 14539 30092 14607 30148
rect 14663 30092 14673 30148
rect 12861 30024 14673 30092
rect 12861 29968 12871 30024
rect 12927 29968 12995 30024
rect 13051 29968 13119 30024
rect 13175 29968 13243 30024
rect 13299 29968 13367 30024
rect 13423 29968 13491 30024
rect 13547 29968 13615 30024
rect 13671 29968 13739 30024
rect 13795 29968 13863 30024
rect 13919 29968 13987 30024
rect 14043 29968 14111 30024
rect 14167 29968 14235 30024
rect 14291 29968 14359 30024
rect 14415 29968 14483 30024
rect 14539 29968 14607 30024
rect 14663 29968 14673 30024
rect 12861 29900 14673 29968
rect 12861 29844 12871 29900
rect 12927 29844 12995 29900
rect 13051 29844 13119 29900
rect 13175 29844 13243 29900
rect 13299 29844 13367 29900
rect 13423 29844 13491 29900
rect 13547 29844 13615 29900
rect 13671 29844 13739 29900
rect 13795 29844 13863 29900
rect 13919 29844 13987 29900
rect 14043 29844 14111 29900
rect 14167 29844 14235 29900
rect 14291 29844 14359 29900
rect 14415 29844 14483 29900
rect 14539 29844 14607 29900
rect 14663 29844 14673 29900
rect 12861 29776 14673 29844
rect 12861 29720 12871 29776
rect 12927 29720 12995 29776
rect 13051 29720 13119 29776
rect 13175 29720 13243 29776
rect 13299 29720 13367 29776
rect 13423 29720 13491 29776
rect 13547 29720 13615 29776
rect 13671 29720 13739 29776
rect 13795 29720 13863 29776
rect 13919 29720 13987 29776
rect 14043 29720 14111 29776
rect 14167 29720 14235 29776
rect 14291 29720 14359 29776
rect 14415 29720 14483 29776
rect 14539 29720 14607 29776
rect 14663 29720 14673 29776
rect 12861 29652 14673 29720
rect 12861 29596 12871 29652
rect 12927 29596 12995 29652
rect 13051 29596 13119 29652
rect 13175 29596 13243 29652
rect 13299 29596 13367 29652
rect 13423 29596 13491 29652
rect 13547 29596 13615 29652
rect 13671 29596 13739 29652
rect 13795 29596 13863 29652
rect 13919 29596 13987 29652
rect 14043 29596 14111 29652
rect 14167 29596 14235 29652
rect 14291 29596 14359 29652
rect 14415 29596 14483 29652
rect 14539 29596 14607 29652
rect 14663 29596 14673 29652
rect 12861 29528 14673 29596
rect 12861 29472 12871 29528
rect 12927 29472 12995 29528
rect 13051 29472 13119 29528
rect 13175 29472 13243 29528
rect 13299 29472 13367 29528
rect 13423 29472 13491 29528
rect 13547 29472 13615 29528
rect 13671 29472 13739 29528
rect 13795 29472 13863 29528
rect 13919 29472 13987 29528
rect 14043 29472 14111 29528
rect 14167 29472 14235 29528
rect 14291 29472 14359 29528
rect 14415 29472 14483 29528
rect 14539 29472 14607 29528
rect 14663 29472 14673 29528
rect 12861 29404 14673 29472
rect 12861 29348 12871 29404
rect 12927 29348 12995 29404
rect 13051 29348 13119 29404
rect 13175 29348 13243 29404
rect 13299 29348 13367 29404
rect 13423 29348 13491 29404
rect 13547 29348 13615 29404
rect 13671 29348 13739 29404
rect 13795 29348 13863 29404
rect 13919 29348 13987 29404
rect 14043 29348 14111 29404
rect 14167 29348 14235 29404
rect 14291 29348 14359 29404
rect 14415 29348 14483 29404
rect 14539 29348 14607 29404
rect 14663 29348 14673 29404
rect 12861 29280 14673 29348
rect 12861 29224 12871 29280
rect 12927 29224 12995 29280
rect 13051 29224 13119 29280
rect 13175 29224 13243 29280
rect 13299 29224 13367 29280
rect 13423 29224 13491 29280
rect 13547 29224 13615 29280
rect 13671 29224 13739 29280
rect 13795 29224 13863 29280
rect 13919 29224 13987 29280
rect 14043 29224 14111 29280
rect 14167 29224 14235 29280
rect 14291 29224 14359 29280
rect 14415 29224 14483 29280
rect 14539 29224 14607 29280
rect 14663 29224 14673 29280
rect 12861 29156 14673 29224
rect 12861 29100 12871 29156
rect 12927 29100 12995 29156
rect 13051 29100 13119 29156
rect 13175 29100 13243 29156
rect 13299 29100 13367 29156
rect 13423 29100 13491 29156
rect 13547 29100 13615 29156
rect 13671 29100 13739 29156
rect 13795 29100 13863 29156
rect 13919 29100 13987 29156
rect 14043 29100 14111 29156
rect 14167 29100 14235 29156
rect 14291 29100 14359 29156
rect 14415 29100 14483 29156
rect 14539 29100 14607 29156
rect 14663 29100 14673 29156
rect 12861 29032 14673 29100
rect 12861 28976 12871 29032
rect 12927 28976 12995 29032
rect 13051 28976 13119 29032
rect 13175 28976 13243 29032
rect 13299 28976 13367 29032
rect 13423 28976 13491 29032
rect 13547 28976 13615 29032
rect 13671 28976 13739 29032
rect 13795 28976 13863 29032
rect 13919 28976 13987 29032
rect 14043 28976 14111 29032
rect 14167 28976 14235 29032
rect 14291 28976 14359 29032
rect 14415 28976 14483 29032
rect 14539 28976 14607 29032
rect 14663 28976 14673 29032
rect 12861 28908 14673 28976
rect 12861 28852 12871 28908
rect 12927 28852 12995 28908
rect 13051 28852 13119 28908
rect 13175 28852 13243 28908
rect 13299 28852 13367 28908
rect 13423 28852 13491 28908
rect 13547 28852 13615 28908
rect 13671 28852 13739 28908
rect 13795 28852 13863 28908
rect 13919 28852 13987 28908
rect 14043 28852 14111 28908
rect 14167 28852 14235 28908
rect 14291 28852 14359 28908
rect 14415 28852 14483 28908
rect 14539 28852 14607 28908
rect 14663 28852 14673 28908
rect 12861 28842 14673 28852
rect 2481 28548 2681 28558
rect 2481 28492 2491 28548
rect 2547 28492 2615 28548
rect 2671 28492 2681 28548
rect 2481 28424 2681 28492
rect 2481 28368 2491 28424
rect 2547 28368 2615 28424
rect 2671 28368 2681 28424
rect 2481 28300 2681 28368
rect 2481 28244 2491 28300
rect 2547 28244 2615 28300
rect 2671 28244 2681 28300
rect 2481 28176 2681 28244
rect 2481 28120 2491 28176
rect 2547 28120 2615 28176
rect 2671 28120 2681 28176
rect 2481 28052 2681 28120
rect 2481 27996 2491 28052
rect 2547 27996 2615 28052
rect 2671 27996 2681 28052
rect 2481 27928 2681 27996
rect 2481 27872 2491 27928
rect 2547 27872 2615 27928
rect 2671 27872 2681 27928
rect 2481 27804 2681 27872
rect 2481 27748 2491 27804
rect 2547 27748 2615 27804
rect 2671 27748 2681 27804
rect 2481 27680 2681 27748
rect 2481 27624 2491 27680
rect 2547 27624 2615 27680
rect 2671 27624 2681 27680
rect 2481 27556 2681 27624
rect 2481 27500 2491 27556
rect 2547 27500 2615 27556
rect 2671 27500 2681 27556
rect 2481 27432 2681 27500
rect 2481 27376 2491 27432
rect 2547 27376 2615 27432
rect 2671 27376 2681 27432
rect 2481 27308 2681 27376
rect 2481 27252 2491 27308
rect 2547 27252 2615 27308
rect 2671 27252 2681 27308
rect 2481 27242 2681 27252
rect 4851 28548 5051 28558
rect 4851 28492 4861 28548
rect 4917 28492 4985 28548
rect 5041 28492 5051 28548
rect 4851 28424 5051 28492
rect 4851 28368 4861 28424
rect 4917 28368 4985 28424
rect 5041 28368 5051 28424
rect 4851 28300 5051 28368
rect 4851 28244 4861 28300
rect 4917 28244 4985 28300
rect 5041 28244 5051 28300
rect 4851 28176 5051 28244
rect 4851 28120 4861 28176
rect 4917 28120 4985 28176
rect 5041 28120 5051 28176
rect 4851 28052 5051 28120
rect 4851 27996 4861 28052
rect 4917 27996 4985 28052
rect 5041 27996 5051 28052
rect 4851 27928 5051 27996
rect 4851 27872 4861 27928
rect 4917 27872 4985 27928
rect 5041 27872 5051 27928
rect 4851 27804 5051 27872
rect 4851 27748 4861 27804
rect 4917 27748 4985 27804
rect 5041 27748 5051 27804
rect 4851 27680 5051 27748
rect 4851 27624 4861 27680
rect 4917 27624 4985 27680
rect 5041 27624 5051 27680
rect 4851 27556 5051 27624
rect 4851 27500 4861 27556
rect 4917 27500 4985 27556
rect 5041 27500 5051 27556
rect 4851 27432 5051 27500
rect 4851 27376 4861 27432
rect 4917 27376 4985 27432
rect 5041 27376 5051 27432
rect 4851 27308 5051 27376
rect 4851 27252 4861 27308
rect 4917 27252 4985 27308
rect 5041 27252 5051 27308
rect 4851 27242 5051 27252
rect 7265 28548 7713 28558
rect 7265 28492 7275 28548
rect 7331 28492 7399 28548
rect 7455 28492 7523 28548
rect 7579 28492 7647 28548
rect 7703 28492 7713 28548
rect 7265 28424 7713 28492
rect 7265 28368 7275 28424
rect 7331 28368 7399 28424
rect 7455 28368 7523 28424
rect 7579 28368 7647 28424
rect 7703 28368 7713 28424
rect 7265 28300 7713 28368
rect 7265 28244 7275 28300
rect 7331 28244 7399 28300
rect 7455 28244 7523 28300
rect 7579 28244 7647 28300
rect 7703 28244 7713 28300
rect 7265 28176 7713 28244
rect 7265 28120 7275 28176
rect 7331 28120 7399 28176
rect 7455 28120 7523 28176
rect 7579 28120 7647 28176
rect 7703 28120 7713 28176
rect 7265 28052 7713 28120
rect 7265 27996 7275 28052
rect 7331 27996 7399 28052
rect 7455 27996 7523 28052
rect 7579 27996 7647 28052
rect 7703 27996 7713 28052
rect 7265 27928 7713 27996
rect 7265 27872 7275 27928
rect 7331 27872 7399 27928
rect 7455 27872 7523 27928
rect 7579 27872 7647 27928
rect 7703 27872 7713 27928
rect 7265 27804 7713 27872
rect 7265 27748 7275 27804
rect 7331 27748 7399 27804
rect 7455 27748 7523 27804
rect 7579 27748 7647 27804
rect 7703 27748 7713 27804
rect 7265 27680 7713 27748
rect 7265 27624 7275 27680
rect 7331 27624 7399 27680
rect 7455 27624 7523 27680
rect 7579 27624 7647 27680
rect 7703 27624 7713 27680
rect 7265 27556 7713 27624
rect 7265 27500 7275 27556
rect 7331 27500 7399 27556
rect 7455 27500 7523 27556
rect 7579 27500 7647 27556
rect 7703 27500 7713 27556
rect 7265 27432 7713 27500
rect 7265 27376 7275 27432
rect 7331 27376 7399 27432
rect 7455 27376 7523 27432
rect 7579 27376 7647 27432
rect 7703 27376 7713 27432
rect 7265 27308 7713 27376
rect 7265 27252 7275 27308
rect 7331 27252 7399 27308
rect 7455 27252 7523 27308
rect 7579 27252 7647 27308
rect 7703 27252 7713 27308
rect 7265 27242 7713 27252
rect 9927 28548 10127 28558
rect 9927 28492 9937 28548
rect 9993 28492 10061 28548
rect 10117 28492 10127 28548
rect 9927 28424 10127 28492
rect 9927 28368 9937 28424
rect 9993 28368 10061 28424
rect 10117 28368 10127 28424
rect 9927 28300 10127 28368
rect 9927 28244 9937 28300
rect 9993 28244 10061 28300
rect 10117 28244 10127 28300
rect 9927 28176 10127 28244
rect 9927 28120 9937 28176
rect 9993 28120 10061 28176
rect 10117 28120 10127 28176
rect 9927 28052 10127 28120
rect 9927 27996 9937 28052
rect 9993 27996 10061 28052
rect 10117 27996 10127 28052
rect 9927 27928 10127 27996
rect 9927 27872 9937 27928
rect 9993 27872 10061 27928
rect 10117 27872 10127 27928
rect 9927 27804 10127 27872
rect 9927 27748 9937 27804
rect 9993 27748 10061 27804
rect 10117 27748 10127 27804
rect 9927 27680 10127 27748
rect 9927 27624 9937 27680
rect 9993 27624 10061 27680
rect 10117 27624 10127 27680
rect 9927 27556 10127 27624
rect 9927 27500 9937 27556
rect 9993 27500 10061 27556
rect 10117 27500 10127 27556
rect 9927 27432 10127 27500
rect 9927 27376 9937 27432
rect 9993 27376 10061 27432
rect 10117 27376 10127 27432
rect 9927 27308 10127 27376
rect 9927 27252 9937 27308
rect 9993 27252 10061 27308
rect 10117 27252 10127 27308
rect 9927 27242 10127 27252
rect 12297 28548 12497 28558
rect 12297 28492 12307 28548
rect 12363 28492 12431 28548
rect 12487 28492 12497 28548
rect 12297 28424 12497 28492
rect 12297 28368 12307 28424
rect 12363 28368 12431 28424
rect 12487 28368 12497 28424
rect 12297 28300 12497 28368
rect 12297 28244 12307 28300
rect 12363 28244 12431 28300
rect 12487 28244 12497 28300
rect 12297 28176 12497 28244
rect 12297 28120 12307 28176
rect 12363 28120 12431 28176
rect 12487 28120 12497 28176
rect 12297 28052 12497 28120
rect 12297 27996 12307 28052
rect 12363 27996 12431 28052
rect 12487 27996 12497 28052
rect 12297 27928 12497 27996
rect 12297 27872 12307 27928
rect 12363 27872 12431 27928
rect 12487 27872 12497 27928
rect 12297 27804 12497 27872
rect 12297 27748 12307 27804
rect 12363 27748 12431 27804
rect 12487 27748 12497 27804
rect 12297 27680 12497 27748
rect 12297 27624 12307 27680
rect 12363 27624 12431 27680
rect 12487 27624 12497 27680
rect 12297 27556 12497 27624
rect 12297 27500 12307 27556
rect 12363 27500 12431 27556
rect 12487 27500 12497 27556
rect 12297 27432 12497 27500
rect 12297 27376 12307 27432
rect 12363 27376 12431 27432
rect 12487 27376 12497 27432
rect 12297 27308 12497 27376
rect 12297 27252 12307 27308
rect 12363 27252 12431 27308
rect 12487 27252 12497 27308
rect 12297 27242 12497 27252
rect 305 26954 2117 26964
rect 305 26898 315 26954
rect 371 26898 439 26954
rect 495 26898 563 26954
rect 619 26898 687 26954
rect 743 26898 811 26954
rect 867 26898 935 26954
rect 991 26898 1059 26954
rect 1115 26898 1183 26954
rect 1239 26898 1307 26954
rect 1363 26898 1431 26954
rect 1487 26898 1555 26954
rect 1611 26898 1679 26954
rect 1735 26898 1803 26954
rect 1859 26898 1927 26954
rect 1983 26898 2051 26954
rect 2107 26898 2117 26954
rect 305 26830 2117 26898
rect 305 26774 315 26830
rect 371 26774 439 26830
rect 495 26774 563 26830
rect 619 26774 687 26830
rect 743 26774 811 26830
rect 867 26774 935 26830
rect 991 26774 1059 26830
rect 1115 26774 1183 26830
rect 1239 26774 1307 26830
rect 1363 26774 1431 26830
rect 1487 26774 1555 26830
rect 1611 26774 1679 26830
rect 1735 26774 1803 26830
rect 1859 26774 1927 26830
rect 1983 26774 2051 26830
rect 2107 26774 2117 26830
rect 305 26706 2117 26774
rect 305 26650 315 26706
rect 371 26650 439 26706
rect 495 26650 563 26706
rect 619 26650 687 26706
rect 743 26650 811 26706
rect 867 26650 935 26706
rect 991 26650 1059 26706
rect 1115 26650 1183 26706
rect 1239 26650 1307 26706
rect 1363 26650 1431 26706
rect 1487 26650 1555 26706
rect 1611 26650 1679 26706
rect 1735 26650 1803 26706
rect 1859 26650 1927 26706
rect 1983 26650 2051 26706
rect 2107 26650 2117 26706
rect 305 26582 2117 26650
rect 305 26526 315 26582
rect 371 26526 439 26582
rect 495 26526 563 26582
rect 619 26526 687 26582
rect 743 26526 811 26582
rect 867 26526 935 26582
rect 991 26526 1059 26582
rect 1115 26526 1183 26582
rect 1239 26526 1307 26582
rect 1363 26526 1431 26582
rect 1487 26526 1555 26582
rect 1611 26526 1679 26582
rect 1735 26526 1803 26582
rect 1859 26526 1927 26582
rect 1983 26526 2051 26582
rect 2107 26526 2117 26582
rect 305 26458 2117 26526
rect 305 26402 315 26458
rect 371 26402 439 26458
rect 495 26402 563 26458
rect 619 26402 687 26458
rect 743 26402 811 26458
rect 867 26402 935 26458
rect 991 26402 1059 26458
rect 1115 26402 1183 26458
rect 1239 26402 1307 26458
rect 1363 26402 1431 26458
rect 1487 26402 1555 26458
rect 1611 26402 1679 26458
rect 1735 26402 1803 26458
rect 1859 26402 1927 26458
rect 1983 26402 2051 26458
rect 2107 26402 2117 26458
rect 305 26334 2117 26402
rect 305 26278 315 26334
rect 371 26278 439 26334
rect 495 26278 563 26334
rect 619 26278 687 26334
rect 743 26278 811 26334
rect 867 26278 935 26334
rect 991 26278 1059 26334
rect 1115 26278 1183 26334
rect 1239 26278 1307 26334
rect 1363 26278 1431 26334
rect 1487 26278 1555 26334
rect 1611 26278 1679 26334
rect 1735 26278 1803 26334
rect 1859 26278 1927 26334
rect 1983 26278 2051 26334
rect 2107 26278 2117 26334
rect 305 26210 2117 26278
rect 305 26154 315 26210
rect 371 26154 439 26210
rect 495 26154 563 26210
rect 619 26154 687 26210
rect 743 26154 811 26210
rect 867 26154 935 26210
rect 991 26154 1059 26210
rect 1115 26154 1183 26210
rect 1239 26154 1307 26210
rect 1363 26154 1431 26210
rect 1487 26154 1555 26210
rect 1611 26154 1679 26210
rect 1735 26154 1803 26210
rect 1859 26154 1927 26210
rect 1983 26154 2051 26210
rect 2107 26154 2117 26210
rect 305 26086 2117 26154
rect 305 26030 315 26086
rect 371 26030 439 26086
rect 495 26030 563 26086
rect 619 26030 687 26086
rect 743 26030 811 26086
rect 867 26030 935 26086
rect 991 26030 1059 26086
rect 1115 26030 1183 26086
rect 1239 26030 1307 26086
rect 1363 26030 1431 26086
rect 1487 26030 1555 26086
rect 1611 26030 1679 26086
rect 1735 26030 1803 26086
rect 1859 26030 1927 26086
rect 1983 26030 2051 26086
rect 2107 26030 2117 26086
rect 305 25962 2117 26030
rect 305 25906 315 25962
rect 371 25906 439 25962
rect 495 25906 563 25962
rect 619 25906 687 25962
rect 743 25906 811 25962
rect 867 25906 935 25962
rect 991 25906 1059 25962
rect 1115 25906 1183 25962
rect 1239 25906 1307 25962
rect 1363 25906 1431 25962
rect 1487 25906 1555 25962
rect 1611 25906 1679 25962
rect 1735 25906 1803 25962
rect 1859 25906 1927 25962
rect 1983 25906 2051 25962
rect 2107 25906 2117 25962
rect 305 25838 2117 25906
rect 305 25782 315 25838
rect 371 25782 439 25838
rect 495 25782 563 25838
rect 619 25782 687 25838
rect 743 25782 811 25838
rect 867 25782 935 25838
rect 991 25782 1059 25838
rect 1115 25782 1183 25838
rect 1239 25782 1307 25838
rect 1363 25782 1431 25838
rect 1487 25782 1555 25838
rect 1611 25782 1679 25838
rect 1735 25782 1803 25838
rect 1859 25782 1927 25838
rect 1983 25782 2051 25838
rect 2107 25782 2117 25838
rect 305 25714 2117 25782
rect 305 25658 315 25714
rect 371 25658 439 25714
rect 495 25658 563 25714
rect 619 25658 687 25714
rect 743 25658 811 25714
rect 867 25658 935 25714
rect 991 25658 1059 25714
rect 1115 25658 1183 25714
rect 1239 25658 1307 25714
rect 1363 25658 1431 25714
rect 1487 25658 1555 25714
rect 1611 25658 1679 25714
rect 1735 25658 1803 25714
rect 1859 25658 1927 25714
rect 1983 25658 2051 25714
rect 2107 25658 2117 25714
rect 305 25590 2117 25658
rect 305 25534 315 25590
rect 371 25534 439 25590
rect 495 25534 563 25590
rect 619 25534 687 25590
rect 743 25534 811 25590
rect 867 25534 935 25590
rect 991 25534 1059 25590
rect 1115 25534 1183 25590
rect 1239 25534 1307 25590
rect 1363 25534 1431 25590
rect 1487 25534 1555 25590
rect 1611 25534 1679 25590
rect 1735 25534 1803 25590
rect 1859 25534 1927 25590
rect 1983 25534 2051 25590
rect 2107 25534 2117 25590
rect 305 25466 2117 25534
rect 305 25410 315 25466
rect 371 25410 439 25466
rect 495 25410 563 25466
rect 619 25410 687 25466
rect 743 25410 811 25466
rect 867 25410 935 25466
rect 991 25410 1059 25466
rect 1115 25410 1183 25466
rect 1239 25410 1307 25466
rect 1363 25410 1431 25466
rect 1487 25410 1555 25466
rect 1611 25410 1679 25466
rect 1735 25410 1803 25466
rect 1859 25410 1927 25466
rect 1983 25410 2051 25466
rect 2107 25410 2117 25466
rect 305 25342 2117 25410
rect 305 25286 315 25342
rect 371 25286 439 25342
rect 495 25286 563 25342
rect 619 25286 687 25342
rect 743 25286 811 25342
rect 867 25286 935 25342
rect 991 25286 1059 25342
rect 1115 25286 1183 25342
rect 1239 25286 1307 25342
rect 1363 25286 1431 25342
rect 1487 25286 1555 25342
rect 1611 25286 1679 25342
rect 1735 25286 1803 25342
rect 1859 25286 1927 25342
rect 1983 25286 2051 25342
rect 2107 25286 2117 25342
rect 305 25218 2117 25286
rect 305 25162 315 25218
rect 371 25162 439 25218
rect 495 25162 563 25218
rect 619 25162 687 25218
rect 743 25162 811 25218
rect 867 25162 935 25218
rect 991 25162 1059 25218
rect 1115 25162 1183 25218
rect 1239 25162 1307 25218
rect 1363 25162 1431 25218
rect 1487 25162 1555 25218
rect 1611 25162 1679 25218
rect 1735 25162 1803 25218
rect 1859 25162 1927 25218
rect 1983 25162 2051 25218
rect 2107 25162 2117 25218
rect 305 25094 2117 25162
rect 305 25038 315 25094
rect 371 25038 439 25094
rect 495 25038 563 25094
rect 619 25038 687 25094
rect 743 25038 811 25094
rect 867 25038 935 25094
rect 991 25038 1059 25094
rect 1115 25038 1183 25094
rect 1239 25038 1307 25094
rect 1363 25038 1431 25094
rect 1487 25038 1555 25094
rect 1611 25038 1679 25094
rect 1735 25038 1803 25094
rect 1859 25038 1927 25094
rect 1983 25038 2051 25094
rect 2107 25038 2117 25094
rect 305 24970 2117 25038
rect 305 24914 315 24970
rect 371 24914 439 24970
rect 495 24914 563 24970
rect 619 24914 687 24970
rect 743 24914 811 24970
rect 867 24914 935 24970
rect 991 24914 1059 24970
rect 1115 24914 1183 24970
rect 1239 24914 1307 24970
rect 1363 24914 1431 24970
rect 1487 24914 1555 24970
rect 1611 24914 1679 24970
rect 1735 24914 1803 24970
rect 1859 24914 1927 24970
rect 1983 24914 2051 24970
rect 2107 24914 2117 24970
rect 305 24846 2117 24914
rect 305 24790 315 24846
rect 371 24790 439 24846
rect 495 24790 563 24846
rect 619 24790 687 24846
rect 743 24790 811 24846
rect 867 24790 935 24846
rect 991 24790 1059 24846
rect 1115 24790 1183 24846
rect 1239 24790 1307 24846
rect 1363 24790 1431 24846
rect 1487 24790 1555 24846
rect 1611 24790 1679 24846
rect 1735 24790 1803 24846
rect 1859 24790 1927 24846
rect 1983 24790 2051 24846
rect 2107 24790 2117 24846
rect 305 24722 2117 24790
rect 305 24666 315 24722
rect 371 24666 439 24722
rect 495 24666 563 24722
rect 619 24666 687 24722
rect 743 24666 811 24722
rect 867 24666 935 24722
rect 991 24666 1059 24722
rect 1115 24666 1183 24722
rect 1239 24666 1307 24722
rect 1363 24666 1431 24722
rect 1487 24666 1555 24722
rect 1611 24666 1679 24722
rect 1735 24666 1803 24722
rect 1859 24666 1927 24722
rect 1983 24666 2051 24722
rect 2107 24666 2117 24722
rect 305 24598 2117 24666
rect 305 24542 315 24598
rect 371 24542 439 24598
rect 495 24542 563 24598
rect 619 24542 687 24598
rect 743 24542 811 24598
rect 867 24542 935 24598
rect 991 24542 1059 24598
rect 1115 24542 1183 24598
rect 1239 24542 1307 24598
rect 1363 24542 1431 24598
rect 1487 24542 1555 24598
rect 1611 24542 1679 24598
rect 1735 24542 1803 24598
rect 1859 24542 1927 24598
rect 1983 24542 2051 24598
rect 2107 24542 2117 24598
rect 305 24474 2117 24542
rect 305 24418 315 24474
rect 371 24418 439 24474
rect 495 24418 563 24474
rect 619 24418 687 24474
rect 743 24418 811 24474
rect 867 24418 935 24474
rect 991 24418 1059 24474
rect 1115 24418 1183 24474
rect 1239 24418 1307 24474
rect 1363 24418 1431 24474
rect 1487 24418 1555 24474
rect 1611 24418 1679 24474
rect 1735 24418 1803 24474
rect 1859 24418 1927 24474
rect 1983 24418 2051 24474
rect 2107 24418 2117 24474
rect 305 24350 2117 24418
rect 305 24294 315 24350
rect 371 24294 439 24350
rect 495 24294 563 24350
rect 619 24294 687 24350
rect 743 24294 811 24350
rect 867 24294 935 24350
rect 991 24294 1059 24350
rect 1115 24294 1183 24350
rect 1239 24294 1307 24350
rect 1363 24294 1431 24350
rect 1487 24294 1555 24350
rect 1611 24294 1679 24350
rect 1735 24294 1803 24350
rect 1859 24294 1927 24350
rect 1983 24294 2051 24350
rect 2107 24294 2117 24350
rect 305 24226 2117 24294
rect 305 24170 315 24226
rect 371 24170 439 24226
rect 495 24170 563 24226
rect 619 24170 687 24226
rect 743 24170 811 24226
rect 867 24170 935 24226
rect 991 24170 1059 24226
rect 1115 24170 1183 24226
rect 1239 24170 1307 24226
rect 1363 24170 1431 24226
rect 1487 24170 1555 24226
rect 1611 24170 1679 24226
rect 1735 24170 1803 24226
rect 1859 24170 1927 24226
rect 1983 24170 2051 24226
rect 2107 24170 2117 24226
rect 305 24102 2117 24170
rect 305 24046 315 24102
rect 371 24046 439 24102
rect 495 24046 563 24102
rect 619 24046 687 24102
rect 743 24046 811 24102
rect 867 24046 935 24102
rect 991 24046 1059 24102
rect 1115 24046 1183 24102
rect 1239 24046 1307 24102
rect 1363 24046 1431 24102
rect 1487 24046 1555 24102
rect 1611 24046 1679 24102
rect 1735 24046 1803 24102
rect 1859 24046 1927 24102
rect 1983 24046 2051 24102
rect 2107 24046 2117 24102
rect 305 24036 2117 24046
rect 2798 26954 4734 26964
rect 2798 26898 2808 26954
rect 2864 26898 2932 26954
rect 2988 26898 3056 26954
rect 3112 26898 3180 26954
rect 3236 26898 3304 26954
rect 3360 26898 3428 26954
rect 3484 26898 3552 26954
rect 3608 26898 3676 26954
rect 3732 26898 3800 26954
rect 3856 26898 3924 26954
rect 3980 26898 4048 26954
rect 4104 26898 4172 26954
rect 4228 26898 4296 26954
rect 4352 26898 4420 26954
rect 4476 26898 4544 26954
rect 4600 26898 4668 26954
rect 4724 26898 4734 26954
rect 2798 26830 4734 26898
rect 2798 26774 2808 26830
rect 2864 26774 2932 26830
rect 2988 26774 3056 26830
rect 3112 26774 3180 26830
rect 3236 26774 3304 26830
rect 3360 26774 3428 26830
rect 3484 26774 3552 26830
rect 3608 26774 3676 26830
rect 3732 26774 3800 26830
rect 3856 26774 3924 26830
rect 3980 26774 4048 26830
rect 4104 26774 4172 26830
rect 4228 26774 4296 26830
rect 4352 26774 4420 26830
rect 4476 26774 4544 26830
rect 4600 26774 4668 26830
rect 4724 26774 4734 26830
rect 2798 26706 4734 26774
rect 2798 26650 2808 26706
rect 2864 26650 2932 26706
rect 2988 26650 3056 26706
rect 3112 26650 3180 26706
rect 3236 26650 3304 26706
rect 3360 26650 3428 26706
rect 3484 26650 3552 26706
rect 3608 26650 3676 26706
rect 3732 26650 3800 26706
rect 3856 26650 3924 26706
rect 3980 26650 4048 26706
rect 4104 26650 4172 26706
rect 4228 26650 4296 26706
rect 4352 26650 4420 26706
rect 4476 26650 4544 26706
rect 4600 26650 4668 26706
rect 4724 26650 4734 26706
rect 2798 26582 4734 26650
rect 2798 26526 2808 26582
rect 2864 26526 2932 26582
rect 2988 26526 3056 26582
rect 3112 26526 3180 26582
rect 3236 26526 3304 26582
rect 3360 26526 3428 26582
rect 3484 26526 3552 26582
rect 3608 26526 3676 26582
rect 3732 26526 3800 26582
rect 3856 26526 3924 26582
rect 3980 26526 4048 26582
rect 4104 26526 4172 26582
rect 4228 26526 4296 26582
rect 4352 26526 4420 26582
rect 4476 26526 4544 26582
rect 4600 26526 4668 26582
rect 4724 26526 4734 26582
rect 2798 26458 4734 26526
rect 2798 26402 2808 26458
rect 2864 26402 2932 26458
rect 2988 26402 3056 26458
rect 3112 26402 3180 26458
rect 3236 26402 3304 26458
rect 3360 26402 3428 26458
rect 3484 26402 3552 26458
rect 3608 26402 3676 26458
rect 3732 26402 3800 26458
rect 3856 26402 3924 26458
rect 3980 26402 4048 26458
rect 4104 26402 4172 26458
rect 4228 26402 4296 26458
rect 4352 26402 4420 26458
rect 4476 26402 4544 26458
rect 4600 26402 4668 26458
rect 4724 26402 4734 26458
rect 2798 26334 4734 26402
rect 2798 26278 2808 26334
rect 2864 26278 2932 26334
rect 2988 26278 3056 26334
rect 3112 26278 3180 26334
rect 3236 26278 3304 26334
rect 3360 26278 3428 26334
rect 3484 26278 3552 26334
rect 3608 26278 3676 26334
rect 3732 26278 3800 26334
rect 3856 26278 3924 26334
rect 3980 26278 4048 26334
rect 4104 26278 4172 26334
rect 4228 26278 4296 26334
rect 4352 26278 4420 26334
rect 4476 26278 4544 26334
rect 4600 26278 4668 26334
rect 4724 26278 4734 26334
rect 2798 26210 4734 26278
rect 2798 26154 2808 26210
rect 2864 26154 2932 26210
rect 2988 26154 3056 26210
rect 3112 26154 3180 26210
rect 3236 26154 3304 26210
rect 3360 26154 3428 26210
rect 3484 26154 3552 26210
rect 3608 26154 3676 26210
rect 3732 26154 3800 26210
rect 3856 26154 3924 26210
rect 3980 26154 4048 26210
rect 4104 26154 4172 26210
rect 4228 26154 4296 26210
rect 4352 26154 4420 26210
rect 4476 26154 4544 26210
rect 4600 26154 4668 26210
rect 4724 26154 4734 26210
rect 2798 26086 4734 26154
rect 2798 26030 2808 26086
rect 2864 26030 2932 26086
rect 2988 26030 3056 26086
rect 3112 26030 3180 26086
rect 3236 26030 3304 26086
rect 3360 26030 3428 26086
rect 3484 26030 3552 26086
rect 3608 26030 3676 26086
rect 3732 26030 3800 26086
rect 3856 26030 3924 26086
rect 3980 26030 4048 26086
rect 4104 26030 4172 26086
rect 4228 26030 4296 26086
rect 4352 26030 4420 26086
rect 4476 26030 4544 26086
rect 4600 26030 4668 26086
rect 4724 26030 4734 26086
rect 2798 25962 4734 26030
rect 2798 25906 2808 25962
rect 2864 25906 2932 25962
rect 2988 25906 3056 25962
rect 3112 25906 3180 25962
rect 3236 25906 3304 25962
rect 3360 25906 3428 25962
rect 3484 25906 3552 25962
rect 3608 25906 3676 25962
rect 3732 25906 3800 25962
rect 3856 25906 3924 25962
rect 3980 25906 4048 25962
rect 4104 25906 4172 25962
rect 4228 25906 4296 25962
rect 4352 25906 4420 25962
rect 4476 25906 4544 25962
rect 4600 25906 4668 25962
rect 4724 25906 4734 25962
rect 2798 25838 4734 25906
rect 2798 25782 2808 25838
rect 2864 25782 2932 25838
rect 2988 25782 3056 25838
rect 3112 25782 3180 25838
rect 3236 25782 3304 25838
rect 3360 25782 3428 25838
rect 3484 25782 3552 25838
rect 3608 25782 3676 25838
rect 3732 25782 3800 25838
rect 3856 25782 3924 25838
rect 3980 25782 4048 25838
rect 4104 25782 4172 25838
rect 4228 25782 4296 25838
rect 4352 25782 4420 25838
rect 4476 25782 4544 25838
rect 4600 25782 4668 25838
rect 4724 25782 4734 25838
rect 2798 25714 4734 25782
rect 2798 25658 2808 25714
rect 2864 25658 2932 25714
rect 2988 25658 3056 25714
rect 3112 25658 3180 25714
rect 3236 25658 3304 25714
rect 3360 25658 3428 25714
rect 3484 25658 3552 25714
rect 3608 25658 3676 25714
rect 3732 25658 3800 25714
rect 3856 25658 3924 25714
rect 3980 25658 4048 25714
rect 4104 25658 4172 25714
rect 4228 25658 4296 25714
rect 4352 25658 4420 25714
rect 4476 25658 4544 25714
rect 4600 25658 4668 25714
rect 4724 25658 4734 25714
rect 2798 25590 4734 25658
rect 2798 25534 2808 25590
rect 2864 25534 2932 25590
rect 2988 25534 3056 25590
rect 3112 25534 3180 25590
rect 3236 25534 3304 25590
rect 3360 25534 3428 25590
rect 3484 25534 3552 25590
rect 3608 25534 3676 25590
rect 3732 25534 3800 25590
rect 3856 25534 3924 25590
rect 3980 25534 4048 25590
rect 4104 25534 4172 25590
rect 4228 25534 4296 25590
rect 4352 25534 4420 25590
rect 4476 25534 4544 25590
rect 4600 25534 4668 25590
rect 4724 25534 4734 25590
rect 2798 25466 4734 25534
rect 2798 25410 2808 25466
rect 2864 25410 2932 25466
rect 2988 25410 3056 25466
rect 3112 25410 3180 25466
rect 3236 25410 3304 25466
rect 3360 25410 3428 25466
rect 3484 25410 3552 25466
rect 3608 25410 3676 25466
rect 3732 25410 3800 25466
rect 3856 25410 3924 25466
rect 3980 25410 4048 25466
rect 4104 25410 4172 25466
rect 4228 25410 4296 25466
rect 4352 25410 4420 25466
rect 4476 25410 4544 25466
rect 4600 25410 4668 25466
rect 4724 25410 4734 25466
rect 2798 25342 4734 25410
rect 2798 25286 2808 25342
rect 2864 25286 2932 25342
rect 2988 25286 3056 25342
rect 3112 25286 3180 25342
rect 3236 25286 3304 25342
rect 3360 25286 3428 25342
rect 3484 25286 3552 25342
rect 3608 25286 3676 25342
rect 3732 25286 3800 25342
rect 3856 25286 3924 25342
rect 3980 25286 4048 25342
rect 4104 25286 4172 25342
rect 4228 25286 4296 25342
rect 4352 25286 4420 25342
rect 4476 25286 4544 25342
rect 4600 25286 4668 25342
rect 4724 25286 4734 25342
rect 2798 25218 4734 25286
rect 2798 25162 2808 25218
rect 2864 25162 2932 25218
rect 2988 25162 3056 25218
rect 3112 25162 3180 25218
rect 3236 25162 3304 25218
rect 3360 25162 3428 25218
rect 3484 25162 3552 25218
rect 3608 25162 3676 25218
rect 3732 25162 3800 25218
rect 3856 25162 3924 25218
rect 3980 25162 4048 25218
rect 4104 25162 4172 25218
rect 4228 25162 4296 25218
rect 4352 25162 4420 25218
rect 4476 25162 4544 25218
rect 4600 25162 4668 25218
rect 4724 25162 4734 25218
rect 2798 25094 4734 25162
rect 2798 25038 2808 25094
rect 2864 25038 2932 25094
rect 2988 25038 3056 25094
rect 3112 25038 3180 25094
rect 3236 25038 3304 25094
rect 3360 25038 3428 25094
rect 3484 25038 3552 25094
rect 3608 25038 3676 25094
rect 3732 25038 3800 25094
rect 3856 25038 3924 25094
rect 3980 25038 4048 25094
rect 4104 25038 4172 25094
rect 4228 25038 4296 25094
rect 4352 25038 4420 25094
rect 4476 25038 4544 25094
rect 4600 25038 4668 25094
rect 4724 25038 4734 25094
rect 2798 24970 4734 25038
rect 2798 24914 2808 24970
rect 2864 24914 2932 24970
rect 2988 24914 3056 24970
rect 3112 24914 3180 24970
rect 3236 24914 3304 24970
rect 3360 24914 3428 24970
rect 3484 24914 3552 24970
rect 3608 24914 3676 24970
rect 3732 24914 3800 24970
rect 3856 24914 3924 24970
rect 3980 24914 4048 24970
rect 4104 24914 4172 24970
rect 4228 24914 4296 24970
rect 4352 24914 4420 24970
rect 4476 24914 4544 24970
rect 4600 24914 4668 24970
rect 4724 24914 4734 24970
rect 2798 24846 4734 24914
rect 2798 24790 2808 24846
rect 2864 24790 2932 24846
rect 2988 24790 3056 24846
rect 3112 24790 3180 24846
rect 3236 24790 3304 24846
rect 3360 24790 3428 24846
rect 3484 24790 3552 24846
rect 3608 24790 3676 24846
rect 3732 24790 3800 24846
rect 3856 24790 3924 24846
rect 3980 24790 4048 24846
rect 4104 24790 4172 24846
rect 4228 24790 4296 24846
rect 4352 24790 4420 24846
rect 4476 24790 4544 24846
rect 4600 24790 4668 24846
rect 4724 24790 4734 24846
rect 2798 24722 4734 24790
rect 2798 24666 2808 24722
rect 2864 24666 2932 24722
rect 2988 24666 3056 24722
rect 3112 24666 3180 24722
rect 3236 24666 3304 24722
rect 3360 24666 3428 24722
rect 3484 24666 3552 24722
rect 3608 24666 3676 24722
rect 3732 24666 3800 24722
rect 3856 24666 3924 24722
rect 3980 24666 4048 24722
rect 4104 24666 4172 24722
rect 4228 24666 4296 24722
rect 4352 24666 4420 24722
rect 4476 24666 4544 24722
rect 4600 24666 4668 24722
rect 4724 24666 4734 24722
rect 2798 24598 4734 24666
rect 2798 24542 2808 24598
rect 2864 24542 2932 24598
rect 2988 24542 3056 24598
rect 3112 24542 3180 24598
rect 3236 24542 3304 24598
rect 3360 24542 3428 24598
rect 3484 24542 3552 24598
rect 3608 24542 3676 24598
rect 3732 24542 3800 24598
rect 3856 24542 3924 24598
rect 3980 24542 4048 24598
rect 4104 24542 4172 24598
rect 4228 24542 4296 24598
rect 4352 24542 4420 24598
rect 4476 24542 4544 24598
rect 4600 24542 4668 24598
rect 4724 24542 4734 24598
rect 2798 24474 4734 24542
rect 2798 24418 2808 24474
rect 2864 24418 2932 24474
rect 2988 24418 3056 24474
rect 3112 24418 3180 24474
rect 3236 24418 3304 24474
rect 3360 24418 3428 24474
rect 3484 24418 3552 24474
rect 3608 24418 3676 24474
rect 3732 24418 3800 24474
rect 3856 24418 3924 24474
rect 3980 24418 4048 24474
rect 4104 24418 4172 24474
rect 4228 24418 4296 24474
rect 4352 24418 4420 24474
rect 4476 24418 4544 24474
rect 4600 24418 4668 24474
rect 4724 24418 4734 24474
rect 2798 24350 4734 24418
rect 2798 24294 2808 24350
rect 2864 24294 2932 24350
rect 2988 24294 3056 24350
rect 3112 24294 3180 24350
rect 3236 24294 3304 24350
rect 3360 24294 3428 24350
rect 3484 24294 3552 24350
rect 3608 24294 3676 24350
rect 3732 24294 3800 24350
rect 3856 24294 3924 24350
rect 3980 24294 4048 24350
rect 4104 24294 4172 24350
rect 4228 24294 4296 24350
rect 4352 24294 4420 24350
rect 4476 24294 4544 24350
rect 4600 24294 4668 24350
rect 4724 24294 4734 24350
rect 2798 24226 4734 24294
rect 2798 24170 2808 24226
rect 2864 24170 2932 24226
rect 2988 24170 3056 24226
rect 3112 24170 3180 24226
rect 3236 24170 3304 24226
rect 3360 24170 3428 24226
rect 3484 24170 3552 24226
rect 3608 24170 3676 24226
rect 3732 24170 3800 24226
rect 3856 24170 3924 24226
rect 3980 24170 4048 24226
rect 4104 24170 4172 24226
rect 4228 24170 4296 24226
rect 4352 24170 4420 24226
rect 4476 24170 4544 24226
rect 4600 24170 4668 24226
rect 4724 24170 4734 24226
rect 2798 24102 4734 24170
rect 2798 24046 2808 24102
rect 2864 24046 2932 24102
rect 2988 24046 3056 24102
rect 3112 24046 3180 24102
rect 3236 24046 3304 24102
rect 3360 24046 3428 24102
rect 3484 24046 3552 24102
rect 3608 24046 3676 24102
rect 3732 24046 3800 24102
rect 3856 24046 3924 24102
rect 3980 24046 4048 24102
rect 4104 24046 4172 24102
rect 4228 24046 4296 24102
rect 4352 24046 4420 24102
rect 4476 24046 4544 24102
rect 4600 24046 4668 24102
rect 4724 24046 4734 24102
rect 2798 24036 4734 24046
rect 5168 26954 7104 26964
rect 5168 26898 5178 26954
rect 5234 26898 5302 26954
rect 5358 26898 5426 26954
rect 5482 26898 5550 26954
rect 5606 26898 5674 26954
rect 5730 26898 5798 26954
rect 5854 26898 5922 26954
rect 5978 26898 6046 26954
rect 6102 26898 6170 26954
rect 6226 26898 6294 26954
rect 6350 26898 6418 26954
rect 6474 26898 6542 26954
rect 6598 26898 6666 26954
rect 6722 26898 6790 26954
rect 6846 26898 6914 26954
rect 6970 26898 7038 26954
rect 7094 26898 7104 26954
rect 5168 26830 7104 26898
rect 5168 26774 5178 26830
rect 5234 26774 5302 26830
rect 5358 26774 5426 26830
rect 5482 26774 5550 26830
rect 5606 26774 5674 26830
rect 5730 26774 5798 26830
rect 5854 26774 5922 26830
rect 5978 26774 6046 26830
rect 6102 26774 6170 26830
rect 6226 26774 6294 26830
rect 6350 26774 6418 26830
rect 6474 26774 6542 26830
rect 6598 26774 6666 26830
rect 6722 26774 6790 26830
rect 6846 26774 6914 26830
rect 6970 26774 7038 26830
rect 7094 26774 7104 26830
rect 5168 26706 7104 26774
rect 5168 26650 5178 26706
rect 5234 26650 5302 26706
rect 5358 26650 5426 26706
rect 5482 26650 5550 26706
rect 5606 26650 5674 26706
rect 5730 26650 5798 26706
rect 5854 26650 5922 26706
rect 5978 26650 6046 26706
rect 6102 26650 6170 26706
rect 6226 26650 6294 26706
rect 6350 26650 6418 26706
rect 6474 26650 6542 26706
rect 6598 26650 6666 26706
rect 6722 26650 6790 26706
rect 6846 26650 6914 26706
rect 6970 26650 7038 26706
rect 7094 26650 7104 26706
rect 5168 26582 7104 26650
rect 5168 26526 5178 26582
rect 5234 26526 5302 26582
rect 5358 26526 5426 26582
rect 5482 26526 5550 26582
rect 5606 26526 5674 26582
rect 5730 26526 5798 26582
rect 5854 26526 5922 26582
rect 5978 26526 6046 26582
rect 6102 26526 6170 26582
rect 6226 26526 6294 26582
rect 6350 26526 6418 26582
rect 6474 26526 6542 26582
rect 6598 26526 6666 26582
rect 6722 26526 6790 26582
rect 6846 26526 6914 26582
rect 6970 26526 7038 26582
rect 7094 26526 7104 26582
rect 5168 26458 7104 26526
rect 5168 26402 5178 26458
rect 5234 26402 5302 26458
rect 5358 26402 5426 26458
rect 5482 26402 5550 26458
rect 5606 26402 5674 26458
rect 5730 26402 5798 26458
rect 5854 26402 5922 26458
rect 5978 26402 6046 26458
rect 6102 26402 6170 26458
rect 6226 26402 6294 26458
rect 6350 26402 6418 26458
rect 6474 26402 6542 26458
rect 6598 26402 6666 26458
rect 6722 26402 6790 26458
rect 6846 26402 6914 26458
rect 6970 26402 7038 26458
rect 7094 26402 7104 26458
rect 5168 26334 7104 26402
rect 5168 26278 5178 26334
rect 5234 26278 5302 26334
rect 5358 26278 5426 26334
rect 5482 26278 5550 26334
rect 5606 26278 5674 26334
rect 5730 26278 5798 26334
rect 5854 26278 5922 26334
rect 5978 26278 6046 26334
rect 6102 26278 6170 26334
rect 6226 26278 6294 26334
rect 6350 26278 6418 26334
rect 6474 26278 6542 26334
rect 6598 26278 6666 26334
rect 6722 26278 6790 26334
rect 6846 26278 6914 26334
rect 6970 26278 7038 26334
rect 7094 26278 7104 26334
rect 5168 26210 7104 26278
rect 5168 26154 5178 26210
rect 5234 26154 5302 26210
rect 5358 26154 5426 26210
rect 5482 26154 5550 26210
rect 5606 26154 5674 26210
rect 5730 26154 5798 26210
rect 5854 26154 5922 26210
rect 5978 26154 6046 26210
rect 6102 26154 6170 26210
rect 6226 26154 6294 26210
rect 6350 26154 6418 26210
rect 6474 26154 6542 26210
rect 6598 26154 6666 26210
rect 6722 26154 6790 26210
rect 6846 26154 6914 26210
rect 6970 26154 7038 26210
rect 7094 26154 7104 26210
rect 5168 26086 7104 26154
rect 5168 26030 5178 26086
rect 5234 26030 5302 26086
rect 5358 26030 5426 26086
rect 5482 26030 5550 26086
rect 5606 26030 5674 26086
rect 5730 26030 5798 26086
rect 5854 26030 5922 26086
rect 5978 26030 6046 26086
rect 6102 26030 6170 26086
rect 6226 26030 6294 26086
rect 6350 26030 6418 26086
rect 6474 26030 6542 26086
rect 6598 26030 6666 26086
rect 6722 26030 6790 26086
rect 6846 26030 6914 26086
rect 6970 26030 7038 26086
rect 7094 26030 7104 26086
rect 5168 25962 7104 26030
rect 5168 25906 5178 25962
rect 5234 25906 5302 25962
rect 5358 25906 5426 25962
rect 5482 25906 5550 25962
rect 5606 25906 5674 25962
rect 5730 25906 5798 25962
rect 5854 25906 5922 25962
rect 5978 25906 6046 25962
rect 6102 25906 6170 25962
rect 6226 25906 6294 25962
rect 6350 25906 6418 25962
rect 6474 25906 6542 25962
rect 6598 25906 6666 25962
rect 6722 25906 6790 25962
rect 6846 25906 6914 25962
rect 6970 25906 7038 25962
rect 7094 25906 7104 25962
rect 5168 25838 7104 25906
rect 5168 25782 5178 25838
rect 5234 25782 5302 25838
rect 5358 25782 5426 25838
rect 5482 25782 5550 25838
rect 5606 25782 5674 25838
rect 5730 25782 5798 25838
rect 5854 25782 5922 25838
rect 5978 25782 6046 25838
rect 6102 25782 6170 25838
rect 6226 25782 6294 25838
rect 6350 25782 6418 25838
rect 6474 25782 6542 25838
rect 6598 25782 6666 25838
rect 6722 25782 6790 25838
rect 6846 25782 6914 25838
rect 6970 25782 7038 25838
rect 7094 25782 7104 25838
rect 5168 25714 7104 25782
rect 5168 25658 5178 25714
rect 5234 25658 5302 25714
rect 5358 25658 5426 25714
rect 5482 25658 5550 25714
rect 5606 25658 5674 25714
rect 5730 25658 5798 25714
rect 5854 25658 5922 25714
rect 5978 25658 6046 25714
rect 6102 25658 6170 25714
rect 6226 25658 6294 25714
rect 6350 25658 6418 25714
rect 6474 25658 6542 25714
rect 6598 25658 6666 25714
rect 6722 25658 6790 25714
rect 6846 25658 6914 25714
rect 6970 25658 7038 25714
rect 7094 25658 7104 25714
rect 5168 25590 7104 25658
rect 5168 25534 5178 25590
rect 5234 25534 5302 25590
rect 5358 25534 5426 25590
rect 5482 25534 5550 25590
rect 5606 25534 5674 25590
rect 5730 25534 5798 25590
rect 5854 25534 5922 25590
rect 5978 25534 6046 25590
rect 6102 25534 6170 25590
rect 6226 25534 6294 25590
rect 6350 25534 6418 25590
rect 6474 25534 6542 25590
rect 6598 25534 6666 25590
rect 6722 25534 6790 25590
rect 6846 25534 6914 25590
rect 6970 25534 7038 25590
rect 7094 25534 7104 25590
rect 5168 25466 7104 25534
rect 5168 25410 5178 25466
rect 5234 25410 5302 25466
rect 5358 25410 5426 25466
rect 5482 25410 5550 25466
rect 5606 25410 5674 25466
rect 5730 25410 5798 25466
rect 5854 25410 5922 25466
rect 5978 25410 6046 25466
rect 6102 25410 6170 25466
rect 6226 25410 6294 25466
rect 6350 25410 6418 25466
rect 6474 25410 6542 25466
rect 6598 25410 6666 25466
rect 6722 25410 6790 25466
rect 6846 25410 6914 25466
rect 6970 25410 7038 25466
rect 7094 25410 7104 25466
rect 5168 25342 7104 25410
rect 5168 25286 5178 25342
rect 5234 25286 5302 25342
rect 5358 25286 5426 25342
rect 5482 25286 5550 25342
rect 5606 25286 5674 25342
rect 5730 25286 5798 25342
rect 5854 25286 5922 25342
rect 5978 25286 6046 25342
rect 6102 25286 6170 25342
rect 6226 25286 6294 25342
rect 6350 25286 6418 25342
rect 6474 25286 6542 25342
rect 6598 25286 6666 25342
rect 6722 25286 6790 25342
rect 6846 25286 6914 25342
rect 6970 25286 7038 25342
rect 7094 25286 7104 25342
rect 5168 25218 7104 25286
rect 5168 25162 5178 25218
rect 5234 25162 5302 25218
rect 5358 25162 5426 25218
rect 5482 25162 5550 25218
rect 5606 25162 5674 25218
rect 5730 25162 5798 25218
rect 5854 25162 5922 25218
rect 5978 25162 6046 25218
rect 6102 25162 6170 25218
rect 6226 25162 6294 25218
rect 6350 25162 6418 25218
rect 6474 25162 6542 25218
rect 6598 25162 6666 25218
rect 6722 25162 6790 25218
rect 6846 25162 6914 25218
rect 6970 25162 7038 25218
rect 7094 25162 7104 25218
rect 5168 25094 7104 25162
rect 5168 25038 5178 25094
rect 5234 25038 5302 25094
rect 5358 25038 5426 25094
rect 5482 25038 5550 25094
rect 5606 25038 5674 25094
rect 5730 25038 5798 25094
rect 5854 25038 5922 25094
rect 5978 25038 6046 25094
rect 6102 25038 6170 25094
rect 6226 25038 6294 25094
rect 6350 25038 6418 25094
rect 6474 25038 6542 25094
rect 6598 25038 6666 25094
rect 6722 25038 6790 25094
rect 6846 25038 6914 25094
rect 6970 25038 7038 25094
rect 7094 25038 7104 25094
rect 5168 24970 7104 25038
rect 5168 24914 5178 24970
rect 5234 24914 5302 24970
rect 5358 24914 5426 24970
rect 5482 24914 5550 24970
rect 5606 24914 5674 24970
rect 5730 24914 5798 24970
rect 5854 24914 5922 24970
rect 5978 24914 6046 24970
rect 6102 24914 6170 24970
rect 6226 24914 6294 24970
rect 6350 24914 6418 24970
rect 6474 24914 6542 24970
rect 6598 24914 6666 24970
rect 6722 24914 6790 24970
rect 6846 24914 6914 24970
rect 6970 24914 7038 24970
rect 7094 24914 7104 24970
rect 5168 24846 7104 24914
rect 5168 24790 5178 24846
rect 5234 24790 5302 24846
rect 5358 24790 5426 24846
rect 5482 24790 5550 24846
rect 5606 24790 5674 24846
rect 5730 24790 5798 24846
rect 5854 24790 5922 24846
rect 5978 24790 6046 24846
rect 6102 24790 6170 24846
rect 6226 24790 6294 24846
rect 6350 24790 6418 24846
rect 6474 24790 6542 24846
rect 6598 24790 6666 24846
rect 6722 24790 6790 24846
rect 6846 24790 6914 24846
rect 6970 24790 7038 24846
rect 7094 24790 7104 24846
rect 5168 24722 7104 24790
rect 5168 24666 5178 24722
rect 5234 24666 5302 24722
rect 5358 24666 5426 24722
rect 5482 24666 5550 24722
rect 5606 24666 5674 24722
rect 5730 24666 5798 24722
rect 5854 24666 5922 24722
rect 5978 24666 6046 24722
rect 6102 24666 6170 24722
rect 6226 24666 6294 24722
rect 6350 24666 6418 24722
rect 6474 24666 6542 24722
rect 6598 24666 6666 24722
rect 6722 24666 6790 24722
rect 6846 24666 6914 24722
rect 6970 24666 7038 24722
rect 7094 24666 7104 24722
rect 5168 24598 7104 24666
rect 5168 24542 5178 24598
rect 5234 24542 5302 24598
rect 5358 24542 5426 24598
rect 5482 24542 5550 24598
rect 5606 24542 5674 24598
rect 5730 24542 5798 24598
rect 5854 24542 5922 24598
rect 5978 24542 6046 24598
rect 6102 24542 6170 24598
rect 6226 24542 6294 24598
rect 6350 24542 6418 24598
rect 6474 24542 6542 24598
rect 6598 24542 6666 24598
rect 6722 24542 6790 24598
rect 6846 24542 6914 24598
rect 6970 24542 7038 24598
rect 7094 24542 7104 24598
rect 5168 24474 7104 24542
rect 5168 24418 5178 24474
rect 5234 24418 5302 24474
rect 5358 24418 5426 24474
rect 5482 24418 5550 24474
rect 5606 24418 5674 24474
rect 5730 24418 5798 24474
rect 5854 24418 5922 24474
rect 5978 24418 6046 24474
rect 6102 24418 6170 24474
rect 6226 24418 6294 24474
rect 6350 24418 6418 24474
rect 6474 24418 6542 24474
rect 6598 24418 6666 24474
rect 6722 24418 6790 24474
rect 6846 24418 6914 24474
rect 6970 24418 7038 24474
rect 7094 24418 7104 24474
rect 5168 24350 7104 24418
rect 5168 24294 5178 24350
rect 5234 24294 5302 24350
rect 5358 24294 5426 24350
rect 5482 24294 5550 24350
rect 5606 24294 5674 24350
rect 5730 24294 5798 24350
rect 5854 24294 5922 24350
rect 5978 24294 6046 24350
rect 6102 24294 6170 24350
rect 6226 24294 6294 24350
rect 6350 24294 6418 24350
rect 6474 24294 6542 24350
rect 6598 24294 6666 24350
rect 6722 24294 6790 24350
rect 6846 24294 6914 24350
rect 6970 24294 7038 24350
rect 7094 24294 7104 24350
rect 5168 24226 7104 24294
rect 5168 24170 5178 24226
rect 5234 24170 5302 24226
rect 5358 24170 5426 24226
rect 5482 24170 5550 24226
rect 5606 24170 5674 24226
rect 5730 24170 5798 24226
rect 5854 24170 5922 24226
rect 5978 24170 6046 24226
rect 6102 24170 6170 24226
rect 6226 24170 6294 24226
rect 6350 24170 6418 24226
rect 6474 24170 6542 24226
rect 6598 24170 6666 24226
rect 6722 24170 6790 24226
rect 6846 24170 6914 24226
rect 6970 24170 7038 24226
rect 7094 24170 7104 24226
rect 5168 24102 7104 24170
rect 5168 24046 5178 24102
rect 5234 24046 5302 24102
rect 5358 24046 5426 24102
rect 5482 24046 5550 24102
rect 5606 24046 5674 24102
rect 5730 24046 5798 24102
rect 5854 24046 5922 24102
rect 5978 24046 6046 24102
rect 6102 24046 6170 24102
rect 6226 24046 6294 24102
rect 6350 24046 6418 24102
rect 6474 24046 6542 24102
rect 6598 24046 6666 24102
rect 6722 24046 6790 24102
rect 6846 24046 6914 24102
rect 6970 24046 7038 24102
rect 7094 24046 7104 24102
rect 5168 24036 7104 24046
rect 7874 26954 9810 26964
rect 7874 26898 7884 26954
rect 7940 26898 8008 26954
rect 8064 26898 8132 26954
rect 8188 26898 8256 26954
rect 8312 26898 8380 26954
rect 8436 26898 8504 26954
rect 8560 26898 8628 26954
rect 8684 26898 8752 26954
rect 8808 26898 8876 26954
rect 8932 26898 9000 26954
rect 9056 26898 9124 26954
rect 9180 26898 9248 26954
rect 9304 26898 9372 26954
rect 9428 26898 9496 26954
rect 9552 26898 9620 26954
rect 9676 26898 9744 26954
rect 9800 26898 9810 26954
rect 7874 26830 9810 26898
rect 7874 26774 7884 26830
rect 7940 26774 8008 26830
rect 8064 26774 8132 26830
rect 8188 26774 8256 26830
rect 8312 26774 8380 26830
rect 8436 26774 8504 26830
rect 8560 26774 8628 26830
rect 8684 26774 8752 26830
rect 8808 26774 8876 26830
rect 8932 26774 9000 26830
rect 9056 26774 9124 26830
rect 9180 26774 9248 26830
rect 9304 26774 9372 26830
rect 9428 26774 9496 26830
rect 9552 26774 9620 26830
rect 9676 26774 9744 26830
rect 9800 26774 9810 26830
rect 7874 26706 9810 26774
rect 7874 26650 7884 26706
rect 7940 26650 8008 26706
rect 8064 26650 8132 26706
rect 8188 26650 8256 26706
rect 8312 26650 8380 26706
rect 8436 26650 8504 26706
rect 8560 26650 8628 26706
rect 8684 26650 8752 26706
rect 8808 26650 8876 26706
rect 8932 26650 9000 26706
rect 9056 26650 9124 26706
rect 9180 26650 9248 26706
rect 9304 26650 9372 26706
rect 9428 26650 9496 26706
rect 9552 26650 9620 26706
rect 9676 26650 9744 26706
rect 9800 26650 9810 26706
rect 7874 26582 9810 26650
rect 7874 26526 7884 26582
rect 7940 26526 8008 26582
rect 8064 26526 8132 26582
rect 8188 26526 8256 26582
rect 8312 26526 8380 26582
rect 8436 26526 8504 26582
rect 8560 26526 8628 26582
rect 8684 26526 8752 26582
rect 8808 26526 8876 26582
rect 8932 26526 9000 26582
rect 9056 26526 9124 26582
rect 9180 26526 9248 26582
rect 9304 26526 9372 26582
rect 9428 26526 9496 26582
rect 9552 26526 9620 26582
rect 9676 26526 9744 26582
rect 9800 26526 9810 26582
rect 7874 26458 9810 26526
rect 7874 26402 7884 26458
rect 7940 26402 8008 26458
rect 8064 26402 8132 26458
rect 8188 26402 8256 26458
rect 8312 26402 8380 26458
rect 8436 26402 8504 26458
rect 8560 26402 8628 26458
rect 8684 26402 8752 26458
rect 8808 26402 8876 26458
rect 8932 26402 9000 26458
rect 9056 26402 9124 26458
rect 9180 26402 9248 26458
rect 9304 26402 9372 26458
rect 9428 26402 9496 26458
rect 9552 26402 9620 26458
rect 9676 26402 9744 26458
rect 9800 26402 9810 26458
rect 7874 26334 9810 26402
rect 7874 26278 7884 26334
rect 7940 26278 8008 26334
rect 8064 26278 8132 26334
rect 8188 26278 8256 26334
rect 8312 26278 8380 26334
rect 8436 26278 8504 26334
rect 8560 26278 8628 26334
rect 8684 26278 8752 26334
rect 8808 26278 8876 26334
rect 8932 26278 9000 26334
rect 9056 26278 9124 26334
rect 9180 26278 9248 26334
rect 9304 26278 9372 26334
rect 9428 26278 9496 26334
rect 9552 26278 9620 26334
rect 9676 26278 9744 26334
rect 9800 26278 9810 26334
rect 7874 26210 9810 26278
rect 7874 26154 7884 26210
rect 7940 26154 8008 26210
rect 8064 26154 8132 26210
rect 8188 26154 8256 26210
rect 8312 26154 8380 26210
rect 8436 26154 8504 26210
rect 8560 26154 8628 26210
rect 8684 26154 8752 26210
rect 8808 26154 8876 26210
rect 8932 26154 9000 26210
rect 9056 26154 9124 26210
rect 9180 26154 9248 26210
rect 9304 26154 9372 26210
rect 9428 26154 9496 26210
rect 9552 26154 9620 26210
rect 9676 26154 9744 26210
rect 9800 26154 9810 26210
rect 7874 26086 9810 26154
rect 7874 26030 7884 26086
rect 7940 26030 8008 26086
rect 8064 26030 8132 26086
rect 8188 26030 8256 26086
rect 8312 26030 8380 26086
rect 8436 26030 8504 26086
rect 8560 26030 8628 26086
rect 8684 26030 8752 26086
rect 8808 26030 8876 26086
rect 8932 26030 9000 26086
rect 9056 26030 9124 26086
rect 9180 26030 9248 26086
rect 9304 26030 9372 26086
rect 9428 26030 9496 26086
rect 9552 26030 9620 26086
rect 9676 26030 9744 26086
rect 9800 26030 9810 26086
rect 7874 25962 9810 26030
rect 7874 25906 7884 25962
rect 7940 25906 8008 25962
rect 8064 25906 8132 25962
rect 8188 25906 8256 25962
rect 8312 25906 8380 25962
rect 8436 25906 8504 25962
rect 8560 25906 8628 25962
rect 8684 25906 8752 25962
rect 8808 25906 8876 25962
rect 8932 25906 9000 25962
rect 9056 25906 9124 25962
rect 9180 25906 9248 25962
rect 9304 25906 9372 25962
rect 9428 25906 9496 25962
rect 9552 25906 9620 25962
rect 9676 25906 9744 25962
rect 9800 25906 9810 25962
rect 7874 25838 9810 25906
rect 7874 25782 7884 25838
rect 7940 25782 8008 25838
rect 8064 25782 8132 25838
rect 8188 25782 8256 25838
rect 8312 25782 8380 25838
rect 8436 25782 8504 25838
rect 8560 25782 8628 25838
rect 8684 25782 8752 25838
rect 8808 25782 8876 25838
rect 8932 25782 9000 25838
rect 9056 25782 9124 25838
rect 9180 25782 9248 25838
rect 9304 25782 9372 25838
rect 9428 25782 9496 25838
rect 9552 25782 9620 25838
rect 9676 25782 9744 25838
rect 9800 25782 9810 25838
rect 7874 25714 9810 25782
rect 7874 25658 7884 25714
rect 7940 25658 8008 25714
rect 8064 25658 8132 25714
rect 8188 25658 8256 25714
rect 8312 25658 8380 25714
rect 8436 25658 8504 25714
rect 8560 25658 8628 25714
rect 8684 25658 8752 25714
rect 8808 25658 8876 25714
rect 8932 25658 9000 25714
rect 9056 25658 9124 25714
rect 9180 25658 9248 25714
rect 9304 25658 9372 25714
rect 9428 25658 9496 25714
rect 9552 25658 9620 25714
rect 9676 25658 9744 25714
rect 9800 25658 9810 25714
rect 7874 25590 9810 25658
rect 7874 25534 7884 25590
rect 7940 25534 8008 25590
rect 8064 25534 8132 25590
rect 8188 25534 8256 25590
rect 8312 25534 8380 25590
rect 8436 25534 8504 25590
rect 8560 25534 8628 25590
rect 8684 25534 8752 25590
rect 8808 25534 8876 25590
rect 8932 25534 9000 25590
rect 9056 25534 9124 25590
rect 9180 25534 9248 25590
rect 9304 25534 9372 25590
rect 9428 25534 9496 25590
rect 9552 25534 9620 25590
rect 9676 25534 9744 25590
rect 9800 25534 9810 25590
rect 7874 25466 9810 25534
rect 7874 25410 7884 25466
rect 7940 25410 8008 25466
rect 8064 25410 8132 25466
rect 8188 25410 8256 25466
rect 8312 25410 8380 25466
rect 8436 25410 8504 25466
rect 8560 25410 8628 25466
rect 8684 25410 8752 25466
rect 8808 25410 8876 25466
rect 8932 25410 9000 25466
rect 9056 25410 9124 25466
rect 9180 25410 9248 25466
rect 9304 25410 9372 25466
rect 9428 25410 9496 25466
rect 9552 25410 9620 25466
rect 9676 25410 9744 25466
rect 9800 25410 9810 25466
rect 7874 25342 9810 25410
rect 7874 25286 7884 25342
rect 7940 25286 8008 25342
rect 8064 25286 8132 25342
rect 8188 25286 8256 25342
rect 8312 25286 8380 25342
rect 8436 25286 8504 25342
rect 8560 25286 8628 25342
rect 8684 25286 8752 25342
rect 8808 25286 8876 25342
rect 8932 25286 9000 25342
rect 9056 25286 9124 25342
rect 9180 25286 9248 25342
rect 9304 25286 9372 25342
rect 9428 25286 9496 25342
rect 9552 25286 9620 25342
rect 9676 25286 9744 25342
rect 9800 25286 9810 25342
rect 7874 25218 9810 25286
rect 7874 25162 7884 25218
rect 7940 25162 8008 25218
rect 8064 25162 8132 25218
rect 8188 25162 8256 25218
rect 8312 25162 8380 25218
rect 8436 25162 8504 25218
rect 8560 25162 8628 25218
rect 8684 25162 8752 25218
rect 8808 25162 8876 25218
rect 8932 25162 9000 25218
rect 9056 25162 9124 25218
rect 9180 25162 9248 25218
rect 9304 25162 9372 25218
rect 9428 25162 9496 25218
rect 9552 25162 9620 25218
rect 9676 25162 9744 25218
rect 9800 25162 9810 25218
rect 7874 25094 9810 25162
rect 7874 25038 7884 25094
rect 7940 25038 8008 25094
rect 8064 25038 8132 25094
rect 8188 25038 8256 25094
rect 8312 25038 8380 25094
rect 8436 25038 8504 25094
rect 8560 25038 8628 25094
rect 8684 25038 8752 25094
rect 8808 25038 8876 25094
rect 8932 25038 9000 25094
rect 9056 25038 9124 25094
rect 9180 25038 9248 25094
rect 9304 25038 9372 25094
rect 9428 25038 9496 25094
rect 9552 25038 9620 25094
rect 9676 25038 9744 25094
rect 9800 25038 9810 25094
rect 7874 24970 9810 25038
rect 7874 24914 7884 24970
rect 7940 24914 8008 24970
rect 8064 24914 8132 24970
rect 8188 24914 8256 24970
rect 8312 24914 8380 24970
rect 8436 24914 8504 24970
rect 8560 24914 8628 24970
rect 8684 24914 8752 24970
rect 8808 24914 8876 24970
rect 8932 24914 9000 24970
rect 9056 24914 9124 24970
rect 9180 24914 9248 24970
rect 9304 24914 9372 24970
rect 9428 24914 9496 24970
rect 9552 24914 9620 24970
rect 9676 24914 9744 24970
rect 9800 24914 9810 24970
rect 7874 24846 9810 24914
rect 7874 24790 7884 24846
rect 7940 24790 8008 24846
rect 8064 24790 8132 24846
rect 8188 24790 8256 24846
rect 8312 24790 8380 24846
rect 8436 24790 8504 24846
rect 8560 24790 8628 24846
rect 8684 24790 8752 24846
rect 8808 24790 8876 24846
rect 8932 24790 9000 24846
rect 9056 24790 9124 24846
rect 9180 24790 9248 24846
rect 9304 24790 9372 24846
rect 9428 24790 9496 24846
rect 9552 24790 9620 24846
rect 9676 24790 9744 24846
rect 9800 24790 9810 24846
rect 7874 24722 9810 24790
rect 7874 24666 7884 24722
rect 7940 24666 8008 24722
rect 8064 24666 8132 24722
rect 8188 24666 8256 24722
rect 8312 24666 8380 24722
rect 8436 24666 8504 24722
rect 8560 24666 8628 24722
rect 8684 24666 8752 24722
rect 8808 24666 8876 24722
rect 8932 24666 9000 24722
rect 9056 24666 9124 24722
rect 9180 24666 9248 24722
rect 9304 24666 9372 24722
rect 9428 24666 9496 24722
rect 9552 24666 9620 24722
rect 9676 24666 9744 24722
rect 9800 24666 9810 24722
rect 7874 24598 9810 24666
rect 7874 24542 7884 24598
rect 7940 24542 8008 24598
rect 8064 24542 8132 24598
rect 8188 24542 8256 24598
rect 8312 24542 8380 24598
rect 8436 24542 8504 24598
rect 8560 24542 8628 24598
rect 8684 24542 8752 24598
rect 8808 24542 8876 24598
rect 8932 24542 9000 24598
rect 9056 24542 9124 24598
rect 9180 24542 9248 24598
rect 9304 24542 9372 24598
rect 9428 24542 9496 24598
rect 9552 24542 9620 24598
rect 9676 24542 9744 24598
rect 9800 24542 9810 24598
rect 7874 24474 9810 24542
rect 7874 24418 7884 24474
rect 7940 24418 8008 24474
rect 8064 24418 8132 24474
rect 8188 24418 8256 24474
rect 8312 24418 8380 24474
rect 8436 24418 8504 24474
rect 8560 24418 8628 24474
rect 8684 24418 8752 24474
rect 8808 24418 8876 24474
rect 8932 24418 9000 24474
rect 9056 24418 9124 24474
rect 9180 24418 9248 24474
rect 9304 24418 9372 24474
rect 9428 24418 9496 24474
rect 9552 24418 9620 24474
rect 9676 24418 9744 24474
rect 9800 24418 9810 24474
rect 7874 24350 9810 24418
rect 7874 24294 7884 24350
rect 7940 24294 8008 24350
rect 8064 24294 8132 24350
rect 8188 24294 8256 24350
rect 8312 24294 8380 24350
rect 8436 24294 8504 24350
rect 8560 24294 8628 24350
rect 8684 24294 8752 24350
rect 8808 24294 8876 24350
rect 8932 24294 9000 24350
rect 9056 24294 9124 24350
rect 9180 24294 9248 24350
rect 9304 24294 9372 24350
rect 9428 24294 9496 24350
rect 9552 24294 9620 24350
rect 9676 24294 9744 24350
rect 9800 24294 9810 24350
rect 7874 24226 9810 24294
rect 7874 24170 7884 24226
rect 7940 24170 8008 24226
rect 8064 24170 8132 24226
rect 8188 24170 8256 24226
rect 8312 24170 8380 24226
rect 8436 24170 8504 24226
rect 8560 24170 8628 24226
rect 8684 24170 8752 24226
rect 8808 24170 8876 24226
rect 8932 24170 9000 24226
rect 9056 24170 9124 24226
rect 9180 24170 9248 24226
rect 9304 24170 9372 24226
rect 9428 24170 9496 24226
rect 9552 24170 9620 24226
rect 9676 24170 9744 24226
rect 9800 24170 9810 24226
rect 7874 24102 9810 24170
rect 7874 24046 7884 24102
rect 7940 24046 8008 24102
rect 8064 24046 8132 24102
rect 8188 24046 8256 24102
rect 8312 24046 8380 24102
rect 8436 24046 8504 24102
rect 8560 24046 8628 24102
rect 8684 24046 8752 24102
rect 8808 24046 8876 24102
rect 8932 24046 9000 24102
rect 9056 24046 9124 24102
rect 9180 24046 9248 24102
rect 9304 24046 9372 24102
rect 9428 24046 9496 24102
rect 9552 24046 9620 24102
rect 9676 24046 9744 24102
rect 9800 24046 9810 24102
rect 7874 24036 9810 24046
rect 10244 26954 12180 26964
rect 10244 26898 10254 26954
rect 10310 26898 10378 26954
rect 10434 26898 10502 26954
rect 10558 26898 10626 26954
rect 10682 26898 10750 26954
rect 10806 26898 10874 26954
rect 10930 26898 10998 26954
rect 11054 26898 11122 26954
rect 11178 26898 11246 26954
rect 11302 26898 11370 26954
rect 11426 26898 11494 26954
rect 11550 26898 11618 26954
rect 11674 26898 11742 26954
rect 11798 26898 11866 26954
rect 11922 26898 11990 26954
rect 12046 26898 12114 26954
rect 12170 26898 12180 26954
rect 10244 26830 12180 26898
rect 10244 26774 10254 26830
rect 10310 26774 10378 26830
rect 10434 26774 10502 26830
rect 10558 26774 10626 26830
rect 10682 26774 10750 26830
rect 10806 26774 10874 26830
rect 10930 26774 10998 26830
rect 11054 26774 11122 26830
rect 11178 26774 11246 26830
rect 11302 26774 11370 26830
rect 11426 26774 11494 26830
rect 11550 26774 11618 26830
rect 11674 26774 11742 26830
rect 11798 26774 11866 26830
rect 11922 26774 11990 26830
rect 12046 26774 12114 26830
rect 12170 26774 12180 26830
rect 10244 26706 12180 26774
rect 10244 26650 10254 26706
rect 10310 26650 10378 26706
rect 10434 26650 10502 26706
rect 10558 26650 10626 26706
rect 10682 26650 10750 26706
rect 10806 26650 10874 26706
rect 10930 26650 10998 26706
rect 11054 26650 11122 26706
rect 11178 26650 11246 26706
rect 11302 26650 11370 26706
rect 11426 26650 11494 26706
rect 11550 26650 11618 26706
rect 11674 26650 11742 26706
rect 11798 26650 11866 26706
rect 11922 26650 11990 26706
rect 12046 26650 12114 26706
rect 12170 26650 12180 26706
rect 10244 26582 12180 26650
rect 10244 26526 10254 26582
rect 10310 26526 10378 26582
rect 10434 26526 10502 26582
rect 10558 26526 10626 26582
rect 10682 26526 10750 26582
rect 10806 26526 10874 26582
rect 10930 26526 10998 26582
rect 11054 26526 11122 26582
rect 11178 26526 11246 26582
rect 11302 26526 11370 26582
rect 11426 26526 11494 26582
rect 11550 26526 11618 26582
rect 11674 26526 11742 26582
rect 11798 26526 11866 26582
rect 11922 26526 11990 26582
rect 12046 26526 12114 26582
rect 12170 26526 12180 26582
rect 10244 26458 12180 26526
rect 10244 26402 10254 26458
rect 10310 26402 10378 26458
rect 10434 26402 10502 26458
rect 10558 26402 10626 26458
rect 10682 26402 10750 26458
rect 10806 26402 10874 26458
rect 10930 26402 10998 26458
rect 11054 26402 11122 26458
rect 11178 26402 11246 26458
rect 11302 26402 11370 26458
rect 11426 26402 11494 26458
rect 11550 26402 11618 26458
rect 11674 26402 11742 26458
rect 11798 26402 11866 26458
rect 11922 26402 11990 26458
rect 12046 26402 12114 26458
rect 12170 26402 12180 26458
rect 10244 26334 12180 26402
rect 10244 26278 10254 26334
rect 10310 26278 10378 26334
rect 10434 26278 10502 26334
rect 10558 26278 10626 26334
rect 10682 26278 10750 26334
rect 10806 26278 10874 26334
rect 10930 26278 10998 26334
rect 11054 26278 11122 26334
rect 11178 26278 11246 26334
rect 11302 26278 11370 26334
rect 11426 26278 11494 26334
rect 11550 26278 11618 26334
rect 11674 26278 11742 26334
rect 11798 26278 11866 26334
rect 11922 26278 11990 26334
rect 12046 26278 12114 26334
rect 12170 26278 12180 26334
rect 10244 26210 12180 26278
rect 10244 26154 10254 26210
rect 10310 26154 10378 26210
rect 10434 26154 10502 26210
rect 10558 26154 10626 26210
rect 10682 26154 10750 26210
rect 10806 26154 10874 26210
rect 10930 26154 10998 26210
rect 11054 26154 11122 26210
rect 11178 26154 11246 26210
rect 11302 26154 11370 26210
rect 11426 26154 11494 26210
rect 11550 26154 11618 26210
rect 11674 26154 11742 26210
rect 11798 26154 11866 26210
rect 11922 26154 11990 26210
rect 12046 26154 12114 26210
rect 12170 26154 12180 26210
rect 10244 26086 12180 26154
rect 10244 26030 10254 26086
rect 10310 26030 10378 26086
rect 10434 26030 10502 26086
rect 10558 26030 10626 26086
rect 10682 26030 10750 26086
rect 10806 26030 10874 26086
rect 10930 26030 10998 26086
rect 11054 26030 11122 26086
rect 11178 26030 11246 26086
rect 11302 26030 11370 26086
rect 11426 26030 11494 26086
rect 11550 26030 11618 26086
rect 11674 26030 11742 26086
rect 11798 26030 11866 26086
rect 11922 26030 11990 26086
rect 12046 26030 12114 26086
rect 12170 26030 12180 26086
rect 10244 25962 12180 26030
rect 10244 25906 10254 25962
rect 10310 25906 10378 25962
rect 10434 25906 10502 25962
rect 10558 25906 10626 25962
rect 10682 25906 10750 25962
rect 10806 25906 10874 25962
rect 10930 25906 10998 25962
rect 11054 25906 11122 25962
rect 11178 25906 11246 25962
rect 11302 25906 11370 25962
rect 11426 25906 11494 25962
rect 11550 25906 11618 25962
rect 11674 25906 11742 25962
rect 11798 25906 11866 25962
rect 11922 25906 11990 25962
rect 12046 25906 12114 25962
rect 12170 25906 12180 25962
rect 10244 25838 12180 25906
rect 10244 25782 10254 25838
rect 10310 25782 10378 25838
rect 10434 25782 10502 25838
rect 10558 25782 10626 25838
rect 10682 25782 10750 25838
rect 10806 25782 10874 25838
rect 10930 25782 10998 25838
rect 11054 25782 11122 25838
rect 11178 25782 11246 25838
rect 11302 25782 11370 25838
rect 11426 25782 11494 25838
rect 11550 25782 11618 25838
rect 11674 25782 11742 25838
rect 11798 25782 11866 25838
rect 11922 25782 11990 25838
rect 12046 25782 12114 25838
rect 12170 25782 12180 25838
rect 10244 25714 12180 25782
rect 10244 25658 10254 25714
rect 10310 25658 10378 25714
rect 10434 25658 10502 25714
rect 10558 25658 10626 25714
rect 10682 25658 10750 25714
rect 10806 25658 10874 25714
rect 10930 25658 10998 25714
rect 11054 25658 11122 25714
rect 11178 25658 11246 25714
rect 11302 25658 11370 25714
rect 11426 25658 11494 25714
rect 11550 25658 11618 25714
rect 11674 25658 11742 25714
rect 11798 25658 11866 25714
rect 11922 25658 11990 25714
rect 12046 25658 12114 25714
rect 12170 25658 12180 25714
rect 10244 25590 12180 25658
rect 10244 25534 10254 25590
rect 10310 25534 10378 25590
rect 10434 25534 10502 25590
rect 10558 25534 10626 25590
rect 10682 25534 10750 25590
rect 10806 25534 10874 25590
rect 10930 25534 10998 25590
rect 11054 25534 11122 25590
rect 11178 25534 11246 25590
rect 11302 25534 11370 25590
rect 11426 25534 11494 25590
rect 11550 25534 11618 25590
rect 11674 25534 11742 25590
rect 11798 25534 11866 25590
rect 11922 25534 11990 25590
rect 12046 25534 12114 25590
rect 12170 25534 12180 25590
rect 10244 25466 12180 25534
rect 10244 25410 10254 25466
rect 10310 25410 10378 25466
rect 10434 25410 10502 25466
rect 10558 25410 10626 25466
rect 10682 25410 10750 25466
rect 10806 25410 10874 25466
rect 10930 25410 10998 25466
rect 11054 25410 11122 25466
rect 11178 25410 11246 25466
rect 11302 25410 11370 25466
rect 11426 25410 11494 25466
rect 11550 25410 11618 25466
rect 11674 25410 11742 25466
rect 11798 25410 11866 25466
rect 11922 25410 11990 25466
rect 12046 25410 12114 25466
rect 12170 25410 12180 25466
rect 10244 25342 12180 25410
rect 10244 25286 10254 25342
rect 10310 25286 10378 25342
rect 10434 25286 10502 25342
rect 10558 25286 10626 25342
rect 10682 25286 10750 25342
rect 10806 25286 10874 25342
rect 10930 25286 10998 25342
rect 11054 25286 11122 25342
rect 11178 25286 11246 25342
rect 11302 25286 11370 25342
rect 11426 25286 11494 25342
rect 11550 25286 11618 25342
rect 11674 25286 11742 25342
rect 11798 25286 11866 25342
rect 11922 25286 11990 25342
rect 12046 25286 12114 25342
rect 12170 25286 12180 25342
rect 10244 25218 12180 25286
rect 10244 25162 10254 25218
rect 10310 25162 10378 25218
rect 10434 25162 10502 25218
rect 10558 25162 10626 25218
rect 10682 25162 10750 25218
rect 10806 25162 10874 25218
rect 10930 25162 10998 25218
rect 11054 25162 11122 25218
rect 11178 25162 11246 25218
rect 11302 25162 11370 25218
rect 11426 25162 11494 25218
rect 11550 25162 11618 25218
rect 11674 25162 11742 25218
rect 11798 25162 11866 25218
rect 11922 25162 11990 25218
rect 12046 25162 12114 25218
rect 12170 25162 12180 25218
rect 10244 25094 12180 25162
rect 10244 25038 10254 25094
rect 10310 25038 10378 25094
rect 10434 25038 10502 25094
rect 10558 25038 10626 25094
rect 10682 25038 10750 25094
rect 10806 25038 10874 25094
rect 10930 25038 10998 25094
rect 11054 25038 11122 25094
rect 11178 25038 11246 25094
rect 11302 25038 11370 25094
rect 11426 25038 11494 25094
rect 11550 25038 11618 25094
rect 11674 25038 11742 25094
rect 11798 25038 11866 25094
rect 11922 25038 11990 25094
rect 12046 25038 12114 25094
rect 12170 25038 12180 25094
rect 10244 24970 12180 25038
rect 10244 24914 10254 24970
rect 10310 24914 10378 24970
rect 10434 24914 10502 24970
rect 10558 24914 10626 24970
rect 10682 24914 10750 24970
rect 10806 24914 10874 24970
rect 10930 24914 10998 24970
rect 11054 24914 11122 24970
rect 11178 24914 11246 24970
rect 11302 24914 11370 24970
rect 11426 24914 11494 24970
rect 11550 24914 11618 24970
rect 11674 24914 11742 24970
rect 11798 24914 11866 24970
rect 11922 24914 11990 24970
rect 12046 24914 12114 24970
rect 12170 24914 12180 24970
rect 10244 24846 12180 24914
rect 10244 24790 10254 24846
rect 10310 24790 10378 24846
rect 10434 24790 10502 24846
rect 10558 24790 10626 24846
rect 10682 24790 10750 24846
rect 10806 24790 10874 24846
rect 10930 24790 10998 24846
rect 11054 24790 11122 24846
rect 11178 24790 11246 24846
rect 11302 24790 11370 24846
rect 11426 24790 11494 24846
rect 11550 24790 11618 24846
rect 11674 24790 11742 24846
rect 11798 24790 11866 24846
rect 11922 24790 11990 24846
rect 12046 24790 12114 24846
rect 12170 24790 12180 24846
rect 10244 24722 12180 24790
rect 10244 24666 10254 24722
rect 10310 24666 10378 24722
rect 10434 24666 10502 24722
rect 10558 24666 10626 24722
rect 10682 24666 10750 24722
rect 10806 24666 10874 24722
rect 10930 24666 10998 24722
rect 11054 24666 11122 24722
rect 11178 24666 11246 24722
rect 11302 24666 11370 24722
rect 11426 24666 11494 24722
rect 11550 24666 11618 24722
rect 11674 24666 11742 24722
rect 11798 24666 11866 24722
rect 11922 24666 11990 24722
rect 12046 24666 12114 24722
rect 12170 24666 12180 24722
rect 10244 24598 12180 24666
rect 10244 24542 10254 24598
rect 10310 24542 10378 24598
rect 10434 24542 10502 24598
rect 10558 24542 10626 24598
rect 10682 24542 10750 24598
rect 10806 24542 10874 24598
rect 10930 24542 10998 24598
rect 11054 24542 11122 24598
rect 11178 24542 11246 24598
rect 11302 24542 11370 24598
rect 11426 24542 11494 24598
rect 11550 24542 11618 24598
rect 11674 24542 11742 24598
rect 11798 24542 11866 24598
rect 11922 24542 11990 24598
rect 12046 24542 12114 24598
rect 12170 24542 12180 24598
rect 10244 24474 12180 24542
rect 10244 24418 10254 24474
rect 10310 24418 10378 24474
rect 10434 24418 10502 24474
rect 10558 24418 10626 24474
rect 10682 24418 10750 24474
rect 10806 24418 10874 24474
rect 10930 24418 10998 24474
rect 11054 24418 11122 24474
rect 11178 24418 11246 24474
rect 11302 24418 11370 24474
rect 11426 24418 11494 24474
rect 11550 24418 11618 24474
rect 11674 24418 11742 24474
rect 11798 24418 11866 24474
rect 11922 24418 11990 24474
rect 12046 24418 12114 24474
rect 12170 24418 12180 24474
rect 10244 24350 12180 24418
rect 10244 24294 10254 24350
rect 10310 24294 10378 24350
rect 10434 24294 10502 24350
rect 10558 24294 10626 24350
rect 10682 24294 10750 24350
rect 10806 24294 10874 24350
rect 10930 24294 10998 24350
rect 11054 24294 11122 24350
rect 11178 24294 11246 24350
rect 11302 24294 11370 24350
rect 11426 24294 11494 24350
rect 11550 24294 11618 24350
rect 11674 24294 11742 24350
rect 11798 24294 11866 24350
rect 11922 24294 11990 24350
rect 12046 24294 12114 24350
rect 12170 24294 12180 24350
rect 10244 24226 12180 24294
rect 10244 24170 10254 24226
rect 10310 24170 10378 24226
rect 10434 24170 10502 24226
rect 10558 24170 10626 24226
rect 10682 24170 10750 24226
rect 10806 24170 10874 24226
rect 10930 24170 10998 24226
rect 11054 24170 11122 24226
rect 11178 24170 11246 24226
rect 11302 24170 11370 24226
rect 11426 24170 11494 24226
rect 11550 24170 11618 24226
rect 11674 24170 11742 24226
rect 11798 24170 11866 24226
rect 11922 24170 11990 24226
rect 12046 24170 12114 24226
rect 12170 24170 12180 24226
rect 10244 24102 12180 24170
rect 10244 24046 10254 24102
rect 10310 24046 10378 24102
rect 10434 24046 10502 24102
rect 10558 24046 10626 24102
rect 10682 24046 10750 24102
rect 10806 24046 10874 24102
rect 10930 24046 10998 24102
rect 11054 24046 11122 24102
rect 11178 24046 11246 24102
rect 11302 24046 11370 24102
rect 11426 24046 11494 24102
rect 11550 24046 11618 24102
rect 11674 24046 11742 24102
rect 11798 24046 11866 24102
rect 11922 24046 11990 24102
rect 12046 24046 12114 24102
rect 12170 24046 12180 24102
rect 10244 24036 12180 24046
rect 12861 26954 14673 26964
rect 12861 26898 12871 26954
rect 12927 26898 12995 26954
rect 13051 26898 13119 26954
rect 13175 26898 13243 26954
rect 13299 26898 13367 26954
rect 13423 26898 13491 26954
rect 13547 26898 13615 26954
rect 13671 26898 13739 26954
rect 13795 26898 13863 26954
rect 13919 26898 13987 26954
rect 14043 26898 14111 26954
rect 14167 26898 14235 26954
rect 14291 26898 14359 26954
rect 14415 26898 14483 26954
rect 14539 26898 14607 26954
rect 14663 26898 14673 26954
rect 12861 26830 14673 26898
rect 12861 26774 12871 26830
rect 12927 26774 12995 26830
rect 13051 26774 13119 26830
rect 13175 26774 13243 26830
rect 13299 26774 13367 26830
rect 13423 26774 13491 26830
rect 13547 26774 13615 26830
rect 13671 26774 13739 26830
rect 13795 26774 13863 26830
rect 13919 26774 13987 26830
rect 14043 26774 14111 26830
rect 14167 26774 14235 26830
rect 14291 26774 14359 26830
rect 14415 26774 14483 26830
rect 14539 26774 14607 26830
rect 14663 26774 14673 26830
rect 12861 26706 14673 26774
rect 12861 26650 12871 26706
rect 12927 26650 12995 26706
rect 13051 26650 13119 26706
rect 13175 26650 13243 26706
rect 13299 26650 13367 26706
rect 13423 26650 13491 26706
rect 13547 26650 13615 26706
rect 13671 26650 13739 26706
rect 13795 26650 13863 26706
rect 13919 26650 13987 26706
rect 14043 26650 14111 26706
rect 14167 26650 14235 26706
rect 14291 26650 14359 26706
rect 14415 26650 14483 26706
rect 14539 26650 14607 26706
rect 14663 26650 14673 26706
rect 12861 26582 14673 26650
rect 12861 26526 12871 26582
rect 12927 26526 12995 26582
rect 13051 26526 13119 26582
rect 13175 26526 13243 26582
rect 13299 26526 13367 26582
rect 13423 26526 13491 26582
rect 13547 26526 13615 26582
rect 13671 26526 13739 26582
rect 13795 26526 13863 26582
rect 13919 26526 13987 26582
rect 14043 26526 14111 26582
rect 14167 26526 14235 26582
rect 14291 26526 14359 26582
rect 14415 26526 14483 26582
rect 14539 26526 14607 26582
rect 14663 26526 14673 26582
rect 12861 26458 14673 26526
rect 12861 26402 12871 26458
rect 12927 26402 12995 26458
rect 13051 26402 13119 26458
rect 13175 26402 13243 26458
rect 13299 26402 13367 26458
rect 13423 26402 13491 26458
rect 13547 26402 13615 26458
rect 13671 26402 13739 26458
rect 13795 26402 13863 26458
rect 13919 26402 13987 26458
rect 14043 26402 14111 26458
rect 14167 26402 14235 26458
rect 14291 26402 14359 26458
rect 14415 26402 14483 26458
rect 14539 26402 14607 26458
rect 14663 26402 14673 26458
rect 12861 26334 14673 26402
rect 12861 26278 12871 26334
rect 12927 26278 12995 26334
rect 13051 26278 13119 26334
rect 13175 26278 13243 26334
rect 13299 26278 13367 26334
rect 13423 26278 13491 26334
rect 13547 26278 13615 26334
rect 13671 26278 13739 26334
rect 13795 26278 13863 26334
rect 13919 26278 13987 26334
rect 14043 26278 14111 26334
rect 14167 26278 14235 26334
rect 14291 26278 14359 26334
rect 14415 26278 14483 26334
rect 14539 26278 14607 26334
rect 14663 26278 14673 26334
rect 12861 26210 14673 26278
rect 12861 26154 12871 26210
rect 12927 26154 12995 26210
rect 13051 26154 13119 26210
rect 13175 26154 13243 26210
rect 13299 26154 13367 26210
rect 13423 26154 13491 26210
rect 13547 26154 13615 26210
rect 13671 26154 13739 26210
rect 13795 26154 13863 26210
rect 13919 26154 13987 26210
rect 14043 26154 14111 26210
rect 14167 26154 14235 26210
rect 14291 26154 14359 26210
rect 14415 26154 14483 26210
rect 14539 26154 14607 26210
rect 14663 26154 14673 26210
rect 12861 26086 14673 26154
rect 12861 26030 12871 26086
rect 12927 26030 12995 26086
rect 13051 26030 13119 26086
rect 13175 26030 13243 26086
rect 13299 26030 13367 26086
rect 13423 26030 13491 26086
rect 13547 26030 13615 26086
rect 13671 26030 13739 26086
rect 13795 26030 13863 26086
rect 13919 26030 13987 26086
rect 14043 26030 14111 26086
rect 14167 26030 14235 26086
rect 14291 26030 14359 26086
rect 14415 26030 14483 26086
rect 14539 26030 14607 26086
rect 14663 26030 14673 26086
rect 12861 25962 14673 26030
rect 12861 25906 12871 25962
rect 12927 25906 12995 25962
rect 13051 25906 13119 25962
rect 13175 25906 13243 25962
rect 13299 25906 13367 25962
rect 13423 25906 13491 25962
rect 13547 25906 13615 25962
rect 13671 25906 13739 25962
rect 13795 25906 13863 25962
rect 13919 25906 13987 25962
rect 14043 25906 14111 25962
rect 14167 25906 14235 25962
rect 14291 25906 14359 25962
rect 14415 25906 14483 25962
rect 14539 25906 14607 25962
rect 14663 25906 14673 25962
rect 12861 25838 14673 25906
rect 12861 25782 12871 25838
rect 12927 25782 12995 25838
rect 13051 25782 13119 25838
rect 13175 25782 13243 25838
rect 13299 25782 13367 25838
rect 13423 25782 13491 25838
rect 13547 25782 13615 25838
rect 13671 25782 13739 25838
rect 13795 25782 13863 25838
rect 13919 25782 13987 25838
rect 14043 25782 14111 25838
rect 14167 25782 14235 25838
rect 14291 25782 14359 25838
rect 14415 25782 14483 25838
rect 14539 25782 14607 25838
rect 14663 25782 14673 25838
rect 12861 25714 14673 25782
rect 12861 25658 12871 25714
rect 12927 25658 12995 25714
rect 13051 25658 13119 25714
rect 13175 25658 13243 25714
rect 13299 25658 13367 25714
rect 13423 25658 13491 25714
rect 13547 25658 13615 25714
rect 13671 25658 13739 25714
rect 13795 25658 13863 25714
rect 13919 25658 13987 25714
rect 14043 25658 14111 25714
rect 14167 25658 14235 25714
rect 14291 25658 14359 25714
rect 14415 25658 14483 25714
rect 14539 25658 14607 25714
rect 14663 25658 14673 25714
rect 12861 25590 14673 25658
rect 12861 25534 12871 25590
rect 12927 25534 12995 25590
rect 13051 25534 13119 25590
rect 13175 25534 13243 25590
rect 13299 25534 13367 25590
rect 13423 25534 13491 25590
rect 13547 25534 13615 25590
rect 13671 25534 13739 25590
rect 13795 25534 13863 25590
rect 13919 25534 13987 25590
rect 14043 25534 14111 25590
rect 14167 25534 14235 25590
rect 14291 25534 14359 25590
rect 14415 25534 14483 25590
rect 14539 25534 14607 25590
rect 14663 25534 14673 25590
rect 12861 25466 14673 25534
rect 12861 25410 12871 25466
rect 12927 25410 12995 25466
rect 13051 25410 13119 25466
rect 13175 25410 13243 25466
rect 13299 25410 13367 25466
rect 13423 25410 13491 25466
rect 13547 25410 13615 25466
rect 13671 25410 13739 25466
rect 13795 25410 13863 25466
rect 13919 25410 13987 25466
rect 14043 25410 14111 25466
rect 14167 25410 14235 25466
rect 14291 25410 14359 25466
rect 14415 25410 14483 25466
rect 14539 25410 14607 25466
rect 14663 25410 14673 25466
rect 12861 25342 14673 25410
rect 12861 25286 12871 25342
rect 12927 25286 12995 25342
rect 13051 25286 13119 25342
rect 13175 25286 13243 25342
rect 13299 25286 13367 25342
rect 13423 25286 13491 25342
rect 13547 25286 13615 25342
rect 13671 25286 13739 25342
rect 13795 25286 13863 25342
rect 13919 25286 13987 25342
rect 14043 25286 14111 25342
rect 14167 25286 14235 25342
rect 14291 25286 14359 25342
rect 14415 25286 14483 25342
rect 14539 25286 14607 25342
rect 14663 25286 14673 25342
rect 12861 25218 14673 25286
rect 12861 25162 12871 25218
rect 12927 25162 12995 25218
rect 13051 25162 13119 25218
rect 13175 25162 13243 25218
rect 13299 25162 13367 25218
rect 13423 25162 13491 25218
rect 13547 25162 13615 25218
rect 13671 25162 13739 25218
rect 13795 25162 13863 25218
rect 13919 25162 13987 25218
rect 14043 25162 14111 25218
rect 14167 25162 14235 25218
rect 14291 25162 14359 25218
rect 14415 25162 14483 25218
rect 14539 25162 14607 25218
rect 14663 25162 14673 25218
rect 12861 25094 14673 25162
rect 12861 25038 12871 25094
rect 12927 25038 12995 25094
rect 13051 25038 13119 25094
rect 13175 25038 13243 25094
rect 13299 25038 13367 25094
rect 13423 25038 13491 25094
rect 13547 25038 13615 25094
rect 13671 25038 13739 25094
rect 13795 25038 13863 25094
rect 13919 25038 13987 25094
rect 14043 25038 14111 25094
rect 14167 25038 14235 25094
rect 14291 25038 14359 25094
rect 14415 25038 14483 25094
rect 14539 25038 14607 25094
rect 14663 25038 14673 25094
rect 12861 24970 14673 25038
rect 12861 24914 12871 24970
rect 12927 24914 12995 24970
rect 13051 24914 13119 24970
rect 13175 24914 13243 24970
rect 13299 24914 13367 24970
rect 13423 24914 13491 24970
rect 13547 24914 13615 24970
rect 13671 24914 13739 24970
rect 13795 24914 13863 24970
rect 13919 24914 13987 24970
rect 14043 24914 14111 24970
rect 14167 24914 14235 24970
rect 14291 24914 14359 24970
rect 14415 24914 14483 24970
rect 14539 24914 14607 24970
rect 14663 24914 14673 24970
rect 12861 24846 14673 24914
rect 12861 24790 12871 24846
rect 12927 24790 12995 24846
rect 13051 24790 13119 24846
rect 13175 24790 13243 24846
rect 13299 24790 13367 24846
rect 13423 24790 13491 24846
rect 13547 24790 13615 24846
rect 13671 24790 13739 24846
rect 13795 24790 13863 24846
rect 13919 24790 13987 24846
rect 14043 24790 14111 24846
rect 14167 24790 14235 24846
rect 14291 24790 14359 24846
rect 14415 24790 14483 24846
rect 14539 24790 14607 24846
rect 14663 24790 14673 24846
rect 12861 24722 14673 24790
rect 12861 24666 12871 24722
rect 12927 24666 12995 24722
rect 13051 24666 13119 24722
rect 13175 24666 13243 24722
rect 13299 24666 13367 24722
rect 13423 24666 13491 24722
rect 13547 24666 13615 24722
rect 13671 24666 13739 24722
rect 13795 24666 13863 24722
rect 13919 24666 13987 24722
rect 14043 24666 14111 24722
rect 14167 24666 14235 24722
rect 14291 24666 14359 24722
rect 14415 24666 14483 24722
rect 14539 24666 14607 24722
rect 14663 24666 14673 24722
rect 12861 24598 14673 24666
rect 12861 24542 12871 24598
rect 12927 24542 12995 24598
rect 13051 24542 13119 24598
rect 13175 24542 13243 24598
rect 13299 24542 13367 24598
rect 13423 24542 13491 24598
rect 13547 24542 13615 24598
rect 13671 24542 13739 24598
rect 13795 24542 13863 24598
rect 13919 24542 13987 24598
rect 14043 24542 14111 24598
rect 14167 24542 14235 24598
rect 14291 24542 14359 24598
rect 14415 24542 14483 24598
rect 14539 24542 14607 24598
rect 14663 24542 14673 24598
rect 12861 24474 14673 24542
rect 12861 24418 12871 24474
rect 12927 24418 12995 24474
rect 13051 24418 13119 24474
rect 13175 24418 13243 24474
rect 13299 24418 13367 24474
rect 13423 24418 13491 24474
rect 13547 24418 13615 24474
rect 13671 24418 13739 24474
rect 13795 24418 13863 24474
rect 13919 24418 13987 24474
rect 14043 24418 14111 24474
rect 14167 24418 14235 24474
rect 14291 24418 14359 24474
rect 14415 24418 14483 24474
rect 14539 24418 14607 24474
rect 14663 24418 14673 24474
rect 12861 24350 14673 24418
rect 12861 24294 12871 24350
rect 12927 24294 12995 24350
rect 13051 24294 13119 24350
rect 13175 24294 13243 24350
rect 13299 24294 13367 24350
rect 13423 24294 13491 24350
rect 13547 24294 13615 24350
rect 13671 24294 13739 24350
rect 13795 24294 13863 24350
rect 13919 24294 13987 24350
rect 14043 24294 14111 24350
rect 14167 24294 14235 24350
rect 14291 24294 14359 24350
rect 14415 24294 14483 24350
rect 14539 24294 14607 24350
rect 14663 24294 14673 24350
rect 12861 24226 14673 24294
rect 12861 24170 12871 24226
rect 12927 24170 12995 24226
rect 13051 24170 13119 24226
rect 13175 24170 13243 24226
rect 13299 24170 13367 24226
rect 13423 24170 13491 24226
rect 13547 24170 13615 24226
rect 13671 24170 13739 24226
rect 13795 24170 13863 24226
rect 13919 24170 13987 24226
rect 14043 24170 14111 24226
rect 14167 24170 14235 24226
rect 14291 24170 14359 24226
rect 14415 24170 14483 24226
rect 14539 24170 14607 24226
rect 14663 24170 14673 24226
rect 12861 24102 14673 24170
rect 12861 24046 12871 24102
rect 12927 24046 12995 24102
rect 13051 24046 13119 24102
rect 13175 24046 13243 24102
rect 13299 24046 13367 24102
rect 13423 24046 13491 24102
rect 13547 24046 13615 24102
rect 13671 24046 13739 24102
rect 13795 24046 13863 24102
rect 13919 24046 13987 24102
rect 14043 24046 14111 24102
rect 14167 24046 14235 24102
rect 14291 24046 14359 24102
rect 14415 24046 14483 24102
rect 14539 24046 14607 24102
rect 14663 24046 14673 24102
rect 12861 24036 14673 24046
rect 305 23754 2117 23764
rect 305 23698 315 23754
rect 371 23698 439 23754
rect 495 23698 563 23754
rect 619 23698 687 23754
rect 743 23698 811 23754
rect 867 23698 935 23754
rect 991 23698 1059 23754
rect 1115 23698 1183 23754
rect 1239 23698 1307 23754
rect 1363 23698 1431 23754
rect 1487 23698 1555 23754
rect 1611 23698 1679 23754
rect 1735 23698 1803 23754
rect 1859 23698 1927 23754
rect 1983 23698 2051 23754
rect 2107 23698 2117 23754
rect 305 23630 2117 23698
rect 305 23574 315 23630
rect 371 23574 439 23630
rect 495 23574 563 23630
rect 619 23574 687 23630
rect 743 23574 811 23630
rect 867 23574 935 23630
rect 991 23574 1059 23630
rect 1115 23574 1183 23630
rect 1239 23574 1307 23630
rect 1363 23574 1431 23630
rect 1487 23574 1555 23630
rect 1611 23574 1679 23630
rect 1735 23574 1803 23630
rect 1859 23574 1927 23630
rect 1983 23574 2051 23630
rect 2107 23574 2117 23630
rect 305 23506 2117 23574
rect 305 23450 315 23506
rect 371 23450 439 23506
rect 495 23450 563 23506
rect 619 23450 687 23506
rect 743 23450 811 23506
rect 867 23450 935 23506
rect 991 23450 1059 23506
rect 1115 23450 1183 23506
rect 1239 23450 1307 23506
rect 1363 23450 1431 23506
rect 1487 23450 1555 23506
rect 1611 23450 1679 23506
rect 1735 23450 1803 23506
rect 1859 23450 1927 23506
rect 1983 23450 2051 23506
rect 2107 23450 2117 23506
rect 305 23382 2117 23450
rect 305 23326 315 23382
rect 371 23326 439 23382
rect 495 23326 563 23382
rect 619 23326 687 23382
rect 743 23326 811 23382
rect 867 23326 935 23382
rect 991 23326 1059 23382
rect 1115 23326 1183 23382
rect 1239 23326 1307 23382
rect 1363 23326 1431 23382
rect 1487 23326 1555 23382
rect 1611 23326 1679 23382
rect 1735 23326 1803 23382
rect 1859 23326 1927 23382
rect 1983 23326 2051 23382
rect 2107 23326 2117 23382
rect 305 23258 2117 23326
rect 305 23202 315 23258
rect 371 23202 439 23258
rect 495 23202 563 23258
rect 619 23202 687 23258
rect 743 23202 811 23258
rect 867 23202 935 23258
rect 991 23202 1059 23258
rect 1115 23202 1183 23258
rect 1239 23202 1307 23258
rect 1363 23202 1431 23258
rect 1487 23202 1555 23258
rect 1611 23202 1679 23258
rect 1735 23202 1803 23258
rect 1859 23202 1927 23258
rect 1983 23202 2051 23258
rect 2107 23202 2117 23258
rect 305 23134 2117 23202
rect 305 23078 315 23134
rect 371 23078 439 23134
rect 495 23078 563 23134
rect 619 23078 687 23134
rect 743 23078 811 23134
rect 867 23078 935 23134
rect 991 23078 1059 23134
rect 1115 23078 1183 23134
rect 1239 23078 1307 23134
rect 1363 23078 1431 23134
rect 1487 23078 1555 23134
rect 1611 23078 1679 23134
rect 1735 23078 1803 23134
rect 1859 23078 1927 23134
rect 1983 23078 2051 23134
rect 2107 23078 2117 23134
rect 305 23010 2117 23078
rect 305 22954 315 23010
rect 371 22954 439 23010
rect 495 22954 563 23010
rect 619 22954 687 23010
rect 743 22954 811 23010
rect 867 22954 935 23010
rect 991 22954 1059 23010
rect 1115 22954 1183 23010
rect 1239 22954 1307 23010
rect 1363 22954 1431 23010
rect 1487 22954 1555 23010
rect 1611 22954 1679 23010
rect 1735 22954 1803 23010
rect 1859 22954 1927 23010
rect 1983 22954 2051 23010
rect 2107 22954 2117 23010
rect 305 22886 2117 22954
rect 305 22830 315 22886
rect 371 22830 439 22886
rect 495 22830 563 22886
rect 619 22830 687 22886
rect 743 22830 811 22886
rect 867 22830 935 22886
rect 991 22830 1059 22886
rect 1115 22830 1183 22886
rect 1239 22830 1307 22886
rect 1363 22830 1431 22886
rect 1487 22830 1555 22886
rect 1611 22830 1679 22886
rect 1735 22830 1803 22886
rect 1859 22830 1927 22886
rect 1983 22830 2051 22886
rect 2107 22830 2117 22886
rect 305 22762 2117 22830
rect 305 22706 315 22762
rect 371 22706 439 22762
rect 495 22706 563 22762
rect 619 22706 687 22762
rect 743 22706 811 22762
rect 867 22706 935 22762
rect 991 22706 1059 22762
rect 1115 22706 1183 22762
rect 1239 22706 1307 22762
rect 1363 22706 1431 22762
rect 1487 22706 1555 22762
rect 1611 22706 1679 22762
rect 1735 22706 1803 22762
rect 1859 22706 1927 22762
rect 1983 22706 2051 22762
rect 2107 22706 2117 22762
rect 305 22638 2117 22706
rect 305 22582 315 22638
rect 371 22582 439 22638
rect 495 22582 563 22638
rect 619 22582 687 22638
rect 743 22582 811 22638
rect 867 22582 935 22638
rect 991 22582 1059 22638
rect 1115 22582 1183 22638
rect 1239 22582 1307 22638
rect 1363 22582 1431 22638
rect 1487 22582 1555 22638
rect 1611 22582 1679 22638
rect 1735 22582 1803 22638
rect 1859 22582 1927 22638
rect 1983 22582 2051 22638
rect 2107 22582 2117 22638
rect 305 22514 2117 22582
rect 305 22458 315 22514
rect 371 22458 439 22514
rect 495 22458 563 22514
rect 619 22458 687 22514
rect 743 22458 811 22514
rect 867 22458 935 22514
rect 991 22458 1059 22514
rect 1115 22458 1183 22514
rect 1239 22458 1307 22514
rect 1363 22458 1431 22514
rect 1487 22458 1555 22514
rect 1611 22458 1679 22514
rect 1735 22458 1803 22514
rect 1859 22458 1927 22514
rect 1983 22458 2051 22514
rect 2107 22458 2117 22514
rect 305 22390 2117 22458
rect 305 22334 315 22390
rect 371 22334 439 22390
rect 495 22334 563 22390
rect 619 22334 687 22390
rect 743 22334 811 22390
rect 867 22334 935 22390
rect 991 22334 1059 22390
rect 1115 22334 1183 22390
rect 1239 22334 1307 22390
rect 1363 22334 1431 22390
rect 1487 22334 1555 22390
rect 1611 22334 1679 22390
rect 1735 22334 1803 22390
rect 1859 22334 1927 22390
rect 1983 22334 2051 22390
rect 2107 22334 2117 22390
rect 305 22266 2117 22334
rect 305 22210 315 22266
rect 371 22210 439 22266
rect 495 22210 563 22266
rect 619 22210 687 22266
rect 743 22210 811 22266
rect 867 22210 935 22266
rect 991 22210 1059 22266
rect 1115 22210 1183 22266
rect 1239 22210 1307 22266
rect 1363 22210 1431 22266
rect 1487 22210 1555 22266
rect 1611 22210 1679 22266
rect 1735 22210 1803 22266
rect 1859 22210 1927 22266
rect 1983 22210 2051 22266
rect 2107 22210 2117 22266
rect 305 22142 2117 22210
rect 305 22086 315 22142
rect 371 22086 439 22142
rect 495 22086 563 22142
rect 619 22086 687 22142
rect 743 22086 811 22142
rect 867 22086 935 22142
rect 991 22086 1059 22142
rect 1115 22086 1183 22142
rect 1239 22086 1307 22142
rect 1363 22086 1431 22142
rect 1487 22086 1555 22142
rect 1611 22086 1679 22142
rect 1735 22086 1803 22142
rect 1859 22086 1927 22142
rect 1983 22086 2051 22142
rect 2107 22086 2117 22142
rect 305 22018 2117 22086
rect 305 21962 315 22018
rect 371 21962 439 22018
rect 495 21962 563 22018
rect 619 21962 687 22018
rect 743 21962 811 22018
rect 867 21962 935 22018
rect 991 21962 1059 22018
rect 1115 21962 1183 22018
rect 1239 21962 1307 22018
rect 1363 21962 1431 22018
rect 1487 21962 1555 22018
rect 1611 21962 1679 22018
rect 1735 21962 1803 22018
rect 1859 21962 1927 22018
rect 1983 21962 2051 22018
rect 2107 21962 2117 22018
rect 305 21894 2117 21962
rect 305 21838 315 21894
rect 371 21838 439 21894
rect 495 21838 563 21894
rect 619 21838 687 21894
rect 743 21838 811 21894
rect 867 21838 935 21894
rect 991 21838 1059 21894
rect 1115 21838 1183 21894
rect 1239 21838 1307 21894
rect 1363 21838 1431 21894
rect 1487 21838 1555 21894
rect 1611 21838 1679 21894
rect 1735 21838 1803 21894
rect 1859 21838 1927 21894
rect 1983 21838 2051 21894
rect 2107 21838 2117 21894
rect 305 21770 2117 21838
rect 305 21714 315 21770
rect 371 21714 439 21770
rect 495 21714 563 21770
rect 619 21714 687 21770
rect 743 21714 811 21770
rect 867 21714 935 21770
rect 991 21714 1059 21770
rect 1115 21714 1183 21770
rect 1239 21714 1307 21770
rect 1363 21714 1431 21770
rect 1487 21714 1555 21770
rect 1611 21714 1679 21770
rect 1735 21714 1803 21770
rect 1859 21714 1927 21770
rect 1983 21714 2051 21770
rect 2107 21714 2117 21770
rect 305 21646 2117 21714
rect 305 21590 315 21646
rect 371 21590 439 21646
rect 495 21590 563 21646
rect 619 21590 687 21646
rect 743 21590 811 21646
rect 867 21590 935 21646
rect 991 21590 1059 21646
rect 1115 21590 1183 21646
rect 1239 21590 1307 21646
rect 1363 21590 1431 21646
rect 1487 21590 1555 21646
rect 1611 21590 1679 21646
rect 1735 21590 1803 21646
rect 1859 21590 1927 21646
rect 1983 21590 2051 21646
rect 2107 21590 2117 21646
rect 305 21522 2117 21590
rect 305 21466 315 21522
rect 371 21466 439 21522
rect 495 21466 563 21522
rect 619 21466 687 21522
rect 743 21466 811 21522
rect 867 21466 935 21522
rect 991 21466 1059 21522
rect 1115 21466 1183 21522
rect 1239 21466 1307 21522
rect 1363 21466 1431 21522
rect 1487 21466 1555 21522
rect 1611 21466 1679 21522
rect 1735 21466 1803 21522
rect 1859 21466 1927 21522
rect 1983 21466 2051 21522
rect 2107 21466 2117 21522
rect 305 21398 2117 21466
rect 305 21342 315 21398
rect 371 21342 439 21398
rect 495 21342 563 21398
rect 619 21342 687 21398
rect 743 21342 811 21398
rect 867 21342 935 21398
rect 991 21342 1059 21398
rect 1115 21342 1183 21398
rect 1239 21342 1307 21398
rect 1363 21342 1431 21398
rect 1487 21342 1555 21398
rect 1611 21342 1679 21398
rect 1735 21342 1803 21398
rect 1859 21342 1927 21398
rect 1983 21342 2051 21398
rect 2107 21342 2117 21398
rect 305 21274 2117 21342
rect 305 21218 315 21274
rect 371 21218 439 21274
rect 495 21218 563 21274
rect 619 21218 687 21274
rect 743 21218 811 21274
rect 867 21218 935 21274
rect 991 21218 1059 21274
rect 1115 21218 1183 21274
rect 1239 21218 1307 21274
rect 1363 21218 1431 21274
rect 1487 21218 1555 21274
rect 1611 21218 1679 21274
rect 1735 21218 1803 21274
rect 1859 21218 1927 21274
rect 1983 21218 2051 21274
rect 2107 21218 2117 21274
rect 305 21150 2117 21218
rect 305 21094 315 21150
rect 371 21094 439 21150
rect 495 21094 563 21150
rect 619 21094 687 21150
rect 743 21094 811 21150
rect 867 21094 935 21150
rect 991 21094 1059 21150
rect 1115 21094 1183 21150
rect 1239 21094 1307 21150
rect 1363 21094 1431 21150
rect 1487 21094 1555 21150
rect 1611 21094 1679 21150
rect 1735 21094 1803 21150
rect 1859 21094 1927 21150
rect 1983 21094 2051 21150
rect 2107 21094 2117 21150
rect 305 21026 2117 21094
rect 305 20970 315 21026
rect 371 20970 439 21026
rect 495 20970 563 21026
rect 619 20970 687 21026
rect 743 20970 811 21026
rect 867 20970 935 21026
rect 991 20970 1059 21026
rect 1115 20970 1183 21026
rect 1239 20970 1307 21026
rect 1363 20970 1431 21026
rect 1487 20970 1555 21026
rect 1611 20970 1679 21026
rect 1735 20970 1803 21026
rect 1859 20970 1927 21026
rect 1983 20970 2051 21026
rect 2107 20970 2117 21026
rect 305 20902 2117 20970
rect 305 20846 315 20902
rect 371 20846 439 20902
rect 495 20846 563 20902
rect 619 20846 687 20902
rect 743 20846 811 20902
rect 867 20846 935 20902
rect 991 20846 1059 20902
rect 1115 20846 1183 20902
rect 1239 20846 1307 20902
rect 1363 20846 1431 20902
rect 1487 20846 1555 20902
rect 1611 20846 1679 20902
rect 1735 20846 1803 20902
rect 1859 20846 1927 20902
rect 1983 20846 2051 20902
rect 2107 20846 2117 20902
rect 305 20836 2117 20846
rect 2798 23754 4734 23764
rect 2798 23698 2808 23754
rect 2864 23698 2932 23754
rect 2988 23698 3056 23754
rect 3112 23698 3180 23754
rect 3236 23698 3304 23754
rect 3360 23698 3428 23754
rect 3484 23698 3552 23754
rect 3608 23698 3676 23754
rect 3732 23698 3800 23754
rect 3856 23698 3924 23754
rect 3980 23698 4048 23754
rect 4104 23698 4172 23754
rect 4228 23698 4296 23754
rect 4352 23698 4420 23754
rect 4476 23698 4544 23754
rect 4600 23698 4668 23754
rect 4724 23698 4734 23754
rect 2798 23630 4734 23698
rect 2798 23574 2808 23630
rect 2864 23574 2932 23630
rect 2988 23574 3056 23630
rect 3112 23574 3180 23630
rect 3236 23574 3304 23630
rect 3360 23574 3428 23630
rect 3484 23574 3552 23630
rect 3608 23574 3676 23630
rect 3732 23574 3800 23630
rect 3856 23574 3924 23630
rect 3980 23574 4048 23630
rect 4104 23574 4172 23630
rect 4228 23574 4296 23630
rect 4352 23574 4420 23630
rect 4476 23574 4544 23630
rect 4600 23574 4668 23630
rect 4724 23574 4734 23630
rect 2798 23506 4734 23574
rect 2798 23450 2808 23506
rect 2864 23450 2932 23506
rect 2988 23450 3056 23506
rect 3112 23450 3180 23506
rect 3236 23450 3304 23506
rect 3360 23450 3428 23506
rect 3484 23450 3552 23506
rect 3608 23450 3676 23506
rect 3732 23450 3800 23506
rect 3856 23450 3924 23506
rect 3980 23450 4048 23506
rect 4104 23450 4172 23506
rect 4228 23450 4296 23506
rect 4352 23450 4420 23506
rect 4476 23450 4544 23506
rect 4600 23450 4668 23506
rect 4724 23450 4734 23506
rect 2798 23382 4734 23450
rect 2798 23326 2808 23382
rect 2864 23326 2932 23382
rect 2988 23326 3056 23382
rect 3112 23326 3180 23382
rect 3236 23326 3304 23382
rect 3360 23326 3428 23382
rect 3484 23326 3552 23382
rect 3608 23326 3676 23382
rect 3732 23326 3800 23382
rect 3856 23326 3924 23382
rect 3980 23326 4048 23382
rect 4104 23326 4172 23382
rect 4228 23326 4296 23382
rect 4352 23326 4420 23382
rect 4476 23326 4544 23382
rect 4600 23326 4668 23382
rect 4724 23326 4734 23382
rect 2798 23258 4734 23326
rect 2798 23202 2808 23258
rect 2864 23202 2932 23258
rect 2988 23202 3056 23258
rect 3112 23202 3180 23258
rect 3236 23202 3304 23258
rect 3360 23202 3428 23258
rect 3484 23202 3552 23258
rect 3608 23202 3676 23258
rect 3732 23202 3800 23258
rect 3856 23202 3924 23258
rect 3980 23202 4048 23258
rect 4104 23202 4172 23258
rect 4228 23202 4296 23258
rect 4352 23202 4420 23258
rect 4476 23202 4544 23258
rect 4600 23202 4668 23258
rect 4724 23202 4734 23258
rect 2798 23134 4734 23202
rect 2798 23078 2808 23134
rect 2864 23078 2932 23134
rect 2988 23078 3056 23134
rect 3112 23078 3180 23134
rect 3236 23078 3304 23134
rect 3360 23078 3428 23134
rect 3484 23078 3552 23134
rect 3608 23078 3676 23134
rect 3732 23078 3800 23134
rect 3856 23078 3924 23134
rect 3980 23078 4048 23134
rect 4104 23078 4172 23134
rect 4228 23078 4296 23134
rect 4352 23078 4420 23134
rect 4476 23078 4544 23134
rect 4600 23078 4668 23134
rect 4724 23078 4734 23134
rect 2798 23010 4734 23078
rect 2798 22954 2808 23010
rect 2864 22954 2932 23010
rect 2988 22954 3056 23010
rect 3112 22954 3180 23010
rect 3236 22954 3304 23010
rect 3360 22954 3428 23010
rect 3484 22954 3552 23010
rect 3608 22954 3676 23010
rect 3732 22954 3800 23010
rect 3856 22954 3924 23010
rect 3980 22954 4048 23010
rect 4104 22954 4172 23010
rect 4228 22954 4296 23010
rect 4352 22954 4420 23010
rect 4476 22954 4544 23010
rect 4600 22954 4668 23010
rect 4724 22954 4734 23010
rect 2798 22886 4734 22954
rect 2798 22830 2808 22886
rect 2864 22830 2932 22886
rect 2988 22830 3056 22886
rect 3112 22830 3180 22886
rect 3236 22830 3304 22886
rect 3360 22830 3428 22886
rect 3484 22830 3552 22886
rect 3608 22830 3676 22886
rect 3732 22830 3800 22886
rect 3856 22830 3924 22886
rect 3980 22830 4048 22886
rect 4104 22830 4172 22886
rect 4228 22830 4296 22886
rect 4352 22830 4420 22886
rect 4476 22830 4544 22886
rect 4600 22830 4668 22886
rect 4724 22830 4734 22886
rect 2798 22762 4734 22830
rect 2798 22706 2808 22762
rect 2864 22706 2932 22762
rect 2988 22706 3056 22762
rect 3112 22706 3180 22762
rect 3236 22706 3304 22762
rect 3360 22706 3428 22762
rect 3484 22706 3552 22762
rect 3608 22706 3676 22762
rect 3732 22706 3800 22762
rect 3856 22706 3924 22762
rect 3980 22706 4048 22762
rect 4104 22706 4172 22762
rect 4228 22706 4296 22762
rect 4352 22706 4420 22762
rect 4476 22706 4544 22762
rect 4600 22706 4668 22762
rect 4724 22706 4734 22762
rect 2798 22638 4734 22706
rect 2798 22582 2808 22638
rect 2864 22582 2932 22638
rect 2988 22582 3056 22638
rect 3112 22582 3180 22638
rect 3236 22582 3304 22638
rect 3360 22582 3428 22638
rect 3484 22582 3552 22638
rect 3608 22582 3676 22638
rect 3732 22582 3800 22638
rect 3856 22582 3924 22638
rect 3980 22582 4048 22638
rect 4104 22582 4172 22638
rect 4228 22582 4296 22638
rect 4352 22582 4420 22638
rect 4476 22582 4544 22638
rect 4600 22582 4668 22638
rect 4724 22582 4734 22638
rect 2798 22514 4734 22582
rect 2798 22458 2808 22514
rect 2864 22458 2932 22514
rect 2988 22458 3056 22514
rect 3112 22458 3180 22514
rect 3236 22458 3304 22514
rect 3360 22458 3428 22514
rect 3484 22458 3552 22514
rect 3608 22458 3676 22514
rect 3732 22458 3800 22514
rect 3856 22458 3924 22514
rect 3980 22458 4048 22514
rect 4104 22458 4172 22514
rect 4228 22458 4296 22514
rect 4352 22458 4420 22514
rect 4476 22458 4544 22514
rect 4600 22458 4668 22514
rect 4724 22458 4734 22514
rect 2798 22390 4734 22458
rect 2798 22334 2808 22390
rect 2864 22334 2932 22390
rect 2988 22334 3056 22390
rect 3112 22334 3180 22390
rect 3236 22334 3304 22390
rect 3360 22334 3428 22390
rect 3484 22334 3552 22390
rect 3608 22334 3676 22390
rect 3732 22334 3800 22390
rect 3856 22334 3924 22390
rect 3980 22334 4048 22390
rect 4104 22334 4172 22390
rect 4228 22334 4296 22390
rect 4352 22334 4420 22390
rect 4476 22334 4544 22390
rect 4600 22334 4668 22390
rect 4724 22334 4734 22390
rect 2798 22266 4734 22334
rect 2798 22210 2808 22266
rect 2864 22210 2932 22266
rect 2988 22210 3056 22266
rect 3112 22210 3180 22266
rect 3236 22210 3304 22266
rect 3360 22210 3428 22266
rect 3484 22210 3552 22266
rect 3608 22210 3676 22266
rect 3732 22210 3800 22266
rect 3856 22210 3924 22266
rect 3980 22210 4048 22266
rect 4104 22210 4172 22266
rect 4228 22210 4296 22266
rect 4352 22210 4420 22266
rect 4476 22210 4544 22266
rect 4600 22210 4668 22266
rect 4724 22210 4734 22266
rect 2798 22142 4734 22210
rect 2798 22086 2808 22142
rect 2864 22086 2932 22142
rect 2988 22086 3056 22142
rect 3112 22086 3180 22142
rect 3236 22086 3304 22142
rect 3360 22086 3428 22142
rect 3484 22086 3552 22142
rect 3608 22086 3676 22142
rect 3732 22086 3800 22142
rect 3856 22086 3924 22142
rect 3980 22086 4048 22142
rect 4104 22086 4172 22142
rect 4228 22086 4296 22142
rect 4352 22086 4420 22142
rect 4476 22086 4544 22142
rect 4600 22086 4668 22142
rect 4724 22086 4734 22142
rect 2798 22018 4734 22086
rect 2798 21962 2808 22018
rect 2864 21962 2932 22018
rect 2988 21962 3056 22018
rect 3112 21962 3180 22018
rect 3236 21962 3304 22018
rect 3360 21962 3428 22018
rect 3484 21962 3552 22018
rect 3608 21962 3676 22018
rect 3732 21962 3800 22018
rect 3856 21962 3924 22018
rect 3980 21962 4048 22018
rect 4104 21962 4172 22018
rect 4228 21962 4296 22018
rect 4352 21962 4420 22018
rect 4476 21962 4544 22018
rect 4600 21962 4668 22018
rect 4724 21962 4734 22018
rect 2798 21894 4734 21962
rect 2798 21838 2808 21894
rect 2864 21838 2932 21894
rect 2988 21838 3056 21894
rect 3112 21838 3180 21894
rect 3236 21838 3304 21894
rect 3360 21838 3428 21894
rect 3484 21838 3552 21894
rect 3608 21838 3676 21894
rect 3732 21838 3800 21894
rect 3856 21838 3924 21894
rect 3980 21838 4048 21894
rect 4104 21838 4172 21894
rect 4228 21838 4296 21894
rect 4352 21838 4420 21894
rect 4476 21838 4544 21894
rect 4600 21838 4668 21894
rect 4724 21838 4734 21894
rect 2798 21770 4734 21838
rect 2798 21714 2808 21770
rect 2864 21714 2932 21770
rect 2988 21714 3056 21770
rect 3112 21714 3180 21770
rect 3236 21714 3304 21770
rect 3360 21714 3428 21770
rect 3484 21714 3552 21770
rect 3608 21714 3676 21770
rect 3732 21714 3800 21770
rect 3856 21714 3924 21770
rect 3980 21714 4048 21770
rect 4104 21714 4172 21770
rect 4228 21714 4296 21770
rect 4352 21714 4420 21770
rect 4476 21714 4544 21770
rect 4600 21714 4668 21770
rect 4724 21714 4734 21770
rect 2798 21646 4734 21714
rect 2798 21590 2808 21646
rect 2864 21590 2932 21646
rect 2988 21590 3056 21646
rect 3112 21590 3180 21646
rect 3236 21590 3304 21646
rect 3360 21590 3428 21646
rect 3484 21590 3552 21646
rect 3608 21590 3676 21646
rect 3732 21590 3800 21646
rect 3856 21590 3924 21646
rect 3980 21590 4048 21646
rect 4104 21590 4172 21646
rect 4228 21590 4296 21646
rect 4352 21590 4420 21646
rect 4476 21590 4544 21646
rect 4600 21590 4668 21646
rect 4724 21590 4734 21646
rect 2798 21522 4734 21590
rect 2798 21466 2808 21522
rect 2864 21466 2932 21522
rect 2988 21466 3056 21522
rect 3112 21466 3180 21522
rect 3236 21466 3304 21522
rect 3360 21466 3428 21522
rect 3484 21466 3552 21522
rect 3608 21466 3676 21522
rect 3732 21466 3800 21522
rect 3856 21466 3924 21522
rect 3980 21466 4048 21522
rect 4104 21466 4172 21522
rect 4228 21466 4296 21522
rect 4352 21466 4420 21522
rect 4476 21466 4544 21522
rect 4600 21466 4668 21522
rect 4724 21466 4734 21522
rect 2798 21398 4734 21466
rect 2798 21342 2808 21398
rect 2864 21342 2932 21398
rect 2988 21342 3056 21398
rect 3112 21342 3180 21398
rect 3236 21342 3304 21398
rect 3360 21342 3428 21398
rect 3484 21342 3552 21398
rect 3608 21342 3676 21398
rect 3732 21342 3800 21398
rect 3856 21342 3924 21398
rect 3980 21342 4048 21398
rect 4104 21342 4172 21398
rect 4228 21342 4296 21398
rect 4352 21342 4420 21398
rect 4476 21342 4544 21398
rect 4600 21342 4668 21398
rect 4724 21342 4734 21398
rect 2798 21274 4734 21342
rect 2798 21218 2808 21274
rect 2864 21218 2932 21274
rect 2988 21218 3056 21274
rect 3112 21218 3180 21274
rect 3236 21218 3304 21274
rect 3360 21218 3428 21274
rect 3484 21218 3552 21274
rect 3608 21218 3676 21274
rect 3732 21218 3800 21274
rect 3856 21218 3924 21274
rect 3980 21218 4048 21274
rect 4104 21218 4172 21274
rect 4228 21218 4296 21274
rect 4352 21218 4420 21274
rect 4476 21218 4544 21274
rect 4600 21218 4668 21274
rect 4724 21218 4734 21274
rect 2798 21150 4734 21218
rect 2798 21094 2808 21150
rect 2864 21094 2932 21150
rect 2988 21094 3056 21150
rect 3112 21094 3180 21150
rect 3236 21094 3304 21150
rect 3360 21094 3428 21150
rect 3484 21094 3552 21150
rect 3608 21094 3676 21150
rect 3732 21094 3800 21150
rect 3856 21094 3924 21150
rect 3980 21094 4048 21150
rect 4104 21094 4172 21150
rect 4228 21094 4296 21150
rect 4352 21094 4420 21150
rect 4476 21094 4544 21150
rect 4600 21094 4668 21150
rect 4724 21094 4734 21150
rect 2798 21026 4734 21094
rect 2798 20970 2808 21026
rect 2864 20970 2932 21026
rect 2988 20970 3056 21026
rect 3112 20970 3180 21026
rect 3236 20970 3304 21026
rect 3360 20970 3428 21026
rect 3484 20970 3552 21026
rect 3608 20970 3676 21026
rect 3732 20970 3800 21026
rect 3856 20970 3924 21026
rect 3980 20970 4048 21026
rect 4104 20970 4172 21026
rect 4228 20970 4296 21026
rect 4352 20970 4420 21026
rect 4476 20970 4544 21026
rect 4600 20970 4668 21026
rect 4724 20970 4734 21026
rect 2798 20902 4734 20970
rect 2798 20846 2808 20902
rect 2864 20846 2932 20902
rect 2988 20846 3056 20902
rect 3112 20846 3180 20902
rect 3236 20846 3304 20902
rect 3360 20846 3428 20902
rect 3484 20846 3552 20902
rect 3608 20846 3676 20902
rect 3732 20846 3800 20902
rect 3856 20846 3924 20902
rect 3980 20846 4048 20902
rect 4104 20846 4172 20902
rect 4228 20846 4296 20902
rect 4352 20846 4420 20902
rect 4476 20846 4544 20902
rect 4600 20846 4668 20902
rect 4724 20846 4734 20902
rect 2798 20836 4734 20846
rect 5168 23754 7104 23764
rect 5168 23698 5178 23754
rect 5234 23698 5302 23754
rect 5358 23698 5426 23754
rect 5482 23698 5550 23754
rect 5606 23698 5674 23754
rect 5730 23698 5798 23754
rect 5854 23698 5922 23754
rect 5978 23698 6046 23754
rect 6102 23698 6170 23754
rect 6226 23698 6294 23754
rect 6350 23698 6418 23754
rect 6474 23698 6542 23754
rect 6598 23698 6666 23754
rect 6722 23698 6790 23754
rect 6846 23698 6914 23754
rect 6970 23698 7038 23754
rect 7094 23698 7104 23754
rect 5168 23630 7104 23698
rect 5168 23574 5178 23630
rect 5234 23574 5302 23630
rect 5358 23574 5426 23630
rect 5482 23574 5550 23630
rect 5606 23574 5674 23630
rect 5730 23574 5798 23630
rect 5854 23574 5922 23630
rect 5978 23574 6046 23630
rect 6102 23574 6170 23630
rect 6226 23574 6294 23630
rect 6350 23574 6418 23630
rect 6474 23574 6542 23630
rect 6598 23574 6666 23630
rect 6722 23574 6790 23630
rect 6846 23574 6914 23630
rect 6970 23574 7038 23630
rect 7094 23574 7104 23630
rect 5168 23506 7104 23574
rect 5168 23450 5178 23506
rect 5234 23450 5302 23506
rect 5358 23450 5426 23506
rect 5482 23450 5550 23506
rect 5606 23450 5674 23506
rect 5730 23450 5798 23506
rect 5854 23450 5922 23506
rect 5978 23450 6046 23506
rect 6102 23450 6170 23506
rect 6226 23450 6294 23506
rect 6350 23450 6418 23506
rect 6474 23450 6542 23506
rect 6598 23450 6666 23506
rect 6722 23450 6790 23506
rect 6846 23450 6914 23506
rect 6970 23450 7038 23506
rect 7094 23450 7104 23506
rect 5168 23382 7104 23450
rect 5168 23326 5178 23382
rect 5234 23326 5302 23382
rect 5358 23326 5426 23382
rect 5482 23326 5550 23382
rect 5606 23326 5674 23382
rect 5730 23326 5798 23382
rect 5854 23326 5922 23382
rect 5978 23326 6046 23382
rect 6102 23326 6170 23382
rect 6226 23326 6294 23382
rect 6350 23326 6418 23382
rect 6474 23326 6542 23382
rect 6598 23326 6666 23382
rect 6722 23326 6790 23382
rect 6846 23326 6914 23382
rect 6970 23326 7038 23382
rect 7094 23326 7104 23382
rect 5168 23258 7104 23326
rect 5168 23202 5178 23258
rect 5234 23202 5302 23258
rect 5358 23202 5426 23258
rect 5482 23202 5550 23258
rect 5606 23202 5674 23258
rect 5730 23202 5798 23258
rect 5854 23202 5922 23258
rect 5978 23202 6046 23258
rect 6102 23202 6170 23258
rect 6226 23202 6294 23258
rect 6350 23202 6418 23258
rect 6474 23202 6542 23258
rect 6598 23202 6666 23258
rect 6722 23202 6790 23258
rect 6846 23202 6914 23258
rect 6970 23202 7038 23258
rect 7094 23202 7104 23258
rect 5168 23134 7104 23202
rect 5168 23078 5178 23134
rect 5234 23078 5302 23134
rect 5358 23078 5426 23134
rect 5482 23078 5550 23134
rect 5606 23078 5674 23134
rect 5730 23078 5798 23134
rect 5854 23078 5922 23134
rect 5978 23078 6046 23134
rect 6102 23078 6170 23134
rect 6226 23078 6294 23134
rect 6350 23078 6418 23134
rect 6474 23078 6542 23134
rect 6598 23078 6666 23134
rect 6722 23078 6790 23134
rect 6846 23078 6914 23134
rect 6970 23078 7038 23134
rect 7094 23078 7104 23134
rect 5168 23010 7104 23078
rect 5168 22954 5178 23010
rect 5234 22954 5302 23010
rect 5358 22954 5426 23010
rect 5482 22954 5550 23010
rect 5606 22954 5674 23010
rect 5730 22954 5798 23010
rect 5854 22954 5922 23010
rect 5978 22954 6046 23010
rect 6102 22954 6170 23010
rect 6226 22954 6294 23010
rect 6350 22954 6418 23010
rect 6474 22954 6542 23010
rect 6598 22954 6666 23010
rect 6722 22954 6790 23010
rect 6846 22954 6914 23010
rect 6970 22954 7038 23010
rect 7094 22954 7104 23010
rect 5168 22886 7104 22954
rect 5168 22830 5178 22886
rect 5234 22830 5302 22886
rect 5358 22830 5426 22886
rect 5482 22830 5550 22886
rect 5606 22830 5674 22886
rect 5730 22830 5798 22886
rect 5854 22830 5922 22886
rect 5978 22830 6046 22886
rect 6102 22830 6170 22886
rect 6226 22830 6294 22886
rect 6350 22830 6418 22886
rect 6474 22830 6542 22886
rect 6598 22830 6666 22886
rect 6722 22830 6790 22886
rect 6846 22830 6914 22886
rect 6970 22830 7038 22886
rect 7094 22830 7104 22886
rect 5168 22762 7104 22830
rect 5168 22706 5178 22762
rect 5234 22706 5302 22762
rect 5358 22706 5426 22762
rect 5482 22706 5550 22762
rect 5606 22706 5674 22762
rect 5730 22706 5798 22762
rect 5854 22706 5922 22762
rect 5978 22706 6046 22762
rect 6102 22706 6170 22762
rect 6226 22706 6294 22762
rect 6350 22706 6418 22762
rect 6474 22706 6542 22762
rect 6598 22706 6666 22762
rect 6722 22706 6790 22762
rect 6846 22706 6914 22762
rect 6970 22706 7038 22762
rect 7094 22706 7104 22762
rect 5168 22638 7104 22706
rect 5168 22582 5178 22638
rect 5234 22582 5302 22638
rect 5358 22582 5426 22638
rect 5482 22582 5550 22638
rect 5606 22582 5674 22638
rect 5730 22582 5798 22638
rect 5854 22582 5922 22638
rect 5978 22582 6046 22638
rect 6102 22582 6170 22638
rect 6226 22582 6294 22638
rect 6350 22582 6418 22638
rect 6474 22582 6542 22638
rect 6598 22582 6666 22638
rect 6722 22582 6790 22638
rect 6846 22582 6914 22638
rect 6970 22582 7038 22638
rect 7094 22582 7104 22638
rect 5168 22514 7104 22582
rect 5168 22458 5178 22514
rect 5234 22458 5302 22514
rect 5358 22458 5426 22514
rect 5482 22458 5550 22514
rect 5606 22458 5674 22514
rect 5730 22458 5798 22514
rect 5854 22458 5922 22514
rect 5978 22458 6046 22514
rect 6102 22458 6170 22514
rect 6226 22458 6294 22514
rect 6350 22458 6418 22514
rect 6474 22458 6542 22514
rect 6598 22458 6666 22514
rect 6722 22458 6790 22514
rect 6846 22458 6914 22514
rect 6970 22458 7038 22514
rect 7094 22458 7104 22514
rect 5168 22390 7104 22458
rect 5168 22334 5178 22390
rect 5234 22334 5302 22390
rect 5358 22334 5426 22390
rect 5482 22334 5550 22390
rect 5606 22334 5674 22390
rect 5730 22334 5798 22390
rect 5854 22334 5922 22390
rect 5978 22334 6046 22390
rect 6102 22334 6170 22390
rect 6226 22334 6294 22390
rect 6350 22334 6418 22390
rect 6474 22334 6542 22390
rect 6598 22334 6666 22390
rect 6722 22334 6790 22390
rect 6846 22334 6914 22390
rect 6970 22334 7038 22390
rect 7094 22334 7104 22390
rect 5168 22266 7104 22334
rect 5168 22210 5178 22266
rect 5234 22210 5302 22266
rect 5358 22210 5426 22266
rect 5482 22210 5550 22266
rect 5606 22210 5674 22266
rect 5730 22210 5798 22266
rect 5854 22210 5922 22266
rect 5978 22210 6046 22266
rect 6102 22210 6170 22266
rect 6226 22210 6294 22266
rect 6350 22210 6418 22266
rect 6474 22210 6542 22266
rect 6598 22210 6666 22266
rect 6722 22210 6790 22266
rect 6846 22210 6914 22266
rect 6970 22210 7038 22266
rect 7094 22210 7104 22266
rect 5168 22142 7104 22210
rect 5168 22086 5178 22142
rect 5234 22086 5302 22142
rect 5358 22086 5426 22142
rect 5482 22086 5550 22142
rect 5606 22086 5674 22142
rect 5730 22086 5798 22142
rect 5854 22086 5922 22142
rect 5978 22086 6046 22142
rect 6102 22086 6170 22142
rect 6226 22086 6294 22142
rect 6350 22086 6418 22142
rect 6474 22086 6542 22142
rect 6598 22086 6666 22142
rect 6722 22086 6790 22142
rect 6846 22086 6914 22142
rect 6970 22086 7038 22142
rect 7094 22086 7104 22142
rect 5168 22018 7104 22086
rect 5168 21962 5178 22018
rect 5234 21962 5302 22018
rect 5358 21962 5426 22018
rect 5482 21962 5550 22018
rect 5606 21962 5674 22018
rect 5730 21962 5798 22018
rect 5854 21962 5922 22018
rect 5978 21962 6046 22018
rect 6102 21962 6170 22018
rect 6226 21962 6294 22018
rect 6350 21962 6418 22018
rect 6474 21962 6542 22018
rect 6598 21962 6666 22018
rect 6722 21962 6790 22018
rect 6846 21962 6914 22018
rect 6970 21962 7038 22018
rect 7094 21962 7104 22018
rect 5168 21894 7104 21962
rect 5168 21838 5178 21894
rect 5234 21838 5302 21894
rect 5358 21838 5426 21894
rect 5482 21838 5550 21894
rect 5606 21838 5674 21894
rect 5730 21838 5798 21894
rect 5854 21838 5922 21894
rect 5978 21838 6046 21894
rect 6102 21838 6170 21894
rect 6226 21838 6294 21894
rect 6350 21838 6418 21894
rect 6474 21838 6542 21894
rect 6598 21838 6666 21894
rect 6722 21838 6790 21894
rect 6846 21838 6914 21894
rect 6970 21838 7038 21894
rect 7094 21838 7104 21894
rect 5168 21770 7104 21838
rect 5168 21714 5178 21770
rect 5234 21714 5302 21770
rect 5358 21714 5426 21770
rect 5482 21714 5550 21770
rect 5606 21714 5674 21770
rect 5730 21714 5798 21770
rect 5854 21714 5922 21770
rect 5978 21714 6046 21770
rect 6102 21714 6170 21770
rect 6226 21714 6294 21770
rect 6350 21714 6418 21770
rect 6474 21714 6542 21770
rect 6598 21714 6666 21770
rect 6722 21714 6790 21770
rect 6846 21714 6914 21770
rect 6970 21714 7038 21770
rect 7094 21714 7104 21770
rect 5168 21646 7104 21714
rect 5168 21590 5178 21646
rect 5234 21590 5302 21646
rect 5358 21590 5426 21646
rect 5482 21590 5550 21646
rect 5606 21590 5674 21646
rect 5730 21590 5798 21646
rect 5854 21590 5922 21646
rect 5978 21590 6046 21646
rect 6102 21590 6170 21646
rect 6226 21590 6294 21646
rect 6350 21590 6418 21646
rect 6474 21590 6542 21646
rect 6598 21590 6666 21646
rect 6722 21590 6790 21646
rect 6846 21590 6914 21646
rect 6970 21590 7038 21646
rect 7094 21590 7104 21646
rect 5168 21522 7104 21590
rect 5168 21466 5178 21522
rect 5234 21466 5302 21522
rect 5358 21466 5426 21522
rect 5482 21466 5550 21522
rect 5606 21466 5674 21522
rect 5730 21466 5798 21522
rect 5854 21466 5922 21522
rect 5978 21466 6046 21522
rect 6102 21466 6170 21522
rect 6226 21466 6294 21522
rect 6350 21466 6418 21522
rect 6474 21466 6542 21522
rect 6598 21466 6666 21522
rect 6722 21466 6790 21522
rect 6846 21466 6914 21522
rect 6970 21466 7038 21522
rect 7094 21466 7104 21522
rect 5168 21398 7104 21466
rect 5168 21342 5178 21398
rect 5234 21342 5302 21398
rect 5358 21342 5426 21398
rect 5482 21342 5550 21398
rect 5606 21342 5674 21398
rect 5730 21342 5798 21398
rect 5854 21342 5922 21398
rect 5978 21342 6046 21398
rect 6102 21342 6170 21398
rect 6226 21342 6294 21398
rect 6350 21342 6418 21398
rect 6474 21342 6542 21398
rect 6598 21342 6666 21398
rect 6722 21342 6790 21398
rect 6846 21342 6914 21398
rect 6970 21342 7038 21398
rect 7094 21342 7104 21398
rect 5168 21274 7104 21342
rect 5168 21218 5178 21274
rect 5234 21218 5302 21274
rect 5358 21218 5426 21274
rect 5482 21218 5550 21274
rect 5606 21218 5674 21274
rect 5730 21218 5798 21274
rect 5854 21218 5922 21274
rect 5978 21218 6046 21274
rect 6102 21218 6170 21274
rect 6226 21218 6294 21274
rect 6350 21218 6418 21274
rect 6474 21218 6542 21274
rect 6598 21218 6666 21274
rect 6722 21218 6790 21274
rect 6846 21218 6914 21274
rect 6970 21218 7038 21274
rect 7094 21218 7104 21274
rect 5168 21150 7104 21218
rect 5168 21094 5178 21150
rect 5234 21094 5302 21150
rect 5358 21094 5426 21150
rect 5482 21094 5550 21150
rect 5606 21094 5674 21150
rect 5730 21094 5798 21150
rect 5854 21094 5922 21150
rect 5978 21094 6046 21150
rect 6102 21094 6170 21150
rect 6226 21094 6294 21150
rect 6350 21094 6418 21150
rect 6474 21094 6542 21150
rect 6598 21094 6666 21150
rect 6722 21094 6790 21150
rect 6846 21094 6914 21150
rect 6970 21094 7038 21150
rect 7094 21094 7104 21150
rect 5168 21026 7104 21094
rect 5168 20970 5178 21026
rect 5234 20970 5302 21026
rect 5358 20970 5426 21026
rect 5482 20970 5550 21026
rect 5606 20970 5674 21026
rect 5730 20970 5798 21026
rect 5854 20970 5922 21026
rect 5978 20970 6046 21026
rect 6102 20970 6170 21026
rect 6226 20970 6294 21026
rect 6350 20970 6418 21026
rect 6474 20970 6542 21026
rect 6598 20970 6666 21026
rect 6722 20970 6790 21026
rect 6846 20970 6914 21026
rect 6970 20970 7038 21026
rect 7094 20970 7104 21026
rect 5168 20902 7104 20970
rect 5168 20846 5178 20902
rect 5234 20846 5302 20902
rect 5358 20846 5426 20902
rect 5482 20846 5550 20902
rect 5606 20846 5674 20902
rect 5730 20846 5798 20902
rect 5854 20846 5922 20902
rect 5978 20846 6046 20902
rect 6102 20846 6170 20902
rect 6226 20846 6294 20902
rect 6350 20846 6418 20902
rect 6474 20846 6542 20902
rect 6598 20846 6666 20902
rect 6722 20846 6790 20902
rect 6846 20846 6914 20902
rect 6970 20846 7038 20902
rect 7094 20846 7104 20902
rect 5168 20836 7104 20846
rect 7874 23754 9810 23764
rect 7874 23698 7884 23754
rect 7940 23698 8008 23754
rect 8064 23698 8132 23754
rect 8188 23698 8256 23754
rect 8312 23698 8380 23754
rect 8436 23698 8504 23754
rect 8560 23698 8628 23754
rect 8684 23698 8752 23754
rect 8808 23698 8876 23754
rect 8932 23698 9000 23754
rect 9056 23698 9124 23754
rect 9180 23698 9248 23754
rect 9304 23698 9372 23754
rect 9428 23698 9496 23754
rect 9552 23698 9620 23754
rect 9676 23698 9744 23754
rect 9800 23698 9810 23754
rect 7874 23630 9810 23698
rect 7874 23574 7884 23630
rect 7940 23574 8008 23630
rect 8064 23574 8132 23630
rect 8188 23574 8256 23630
rect 8312 23574 8380 23630
rect 8436 23574 8504 23630
rect 8560 23574 8628 23630
rect 8684 23574 8752 23630
rect 8808 23574 8876 23630
rect 8932 23574 9000 23630
rect 9056 23574 9124 23630
rect 9180 23574 9248 23630
rect 9304 23574 9372 23630
rect 9428 23574 9496 23630
rect 9552 23574 9620 23630
rect 9676 23574 9744 23630
rect 9800 23574 9810 23630
rect 7874 23506 9810 23574
rect 7874 23450 7884 23506
rect 7940 23450 8008 23506
rect 8064 23450 8132 23506
rect 8188 23450 8256 23506
rect 8312 23450 8380 23506
rect 8436 23450 8504 23506
rect 8560 23450 8628 23506
rect 8684 23450 8752 23506
rect 8808 23450 8876 23506
rect 8932 23450 9000 23506
rect 9056 23450 9124 23506
rect 9180 23450 9248 23506
rect 9304 23450 9372 23506
rect 9428 23450 9496 23506
rect 9552 23450 9620 23506
rect 9676 23450 9744 23506
rect 9800 23450 9810 23506
rect 7874 23382 9810 23450
rect 7874 23326 7884 23382
rect 7940 23326 8008 23382
rect 8064 23326 8132 23382
rect 8188 23326 8256 23382
rect 8312 23326 8380 23382
rect 8436 23326 8504 23382
rect 8560 23326 8628 23382
rect 8684 23326 8752 23382
rect 8808 23326 8876 23382
rect 8932 23326 9000 23382
rect 9056 23326 9124 23382
rect 9180 23326 9248 23382
rect 9304 23326 9372 23382
rect 9428 23326 9496 23382
rect 9552 23326 9620 23382
rect 9676 23326 9744 23382
rect 9800 23326 9810 23382
rect 7874 23258 9810 23326
rect 7874 23202 7884 23258
rect 7940 23202 8008 23258
rect 8064 23202 8132 23258
rect 8188 23202 8256 23258
rect 8312 23202 8380 23258
rect 8436 23202 8504 23258
rect 8560 23202 8628 23258
rect 8684 23202 8752 23258
rect 8808 23202 8876 23258
rect 8932 23202 9000 23258
rect 9056 23202 9124 23258
rect 9180 23202 9248 23258
rect 9304 23202 9372 23258
rect 9428 23202 9496 23258
rect 9552 23202 9620 23258
rect 9676 23202 9744 23258
rect 9800 23202 9810 23258
rect 7874 23134 9810 23202
rect 7874 23078 7884 23134
rect 7940 23078 8008 23134
rect 8064 23078 8132 23134
rect 8188 23078 8256 23134
rect 8312 23078 8380 23134
rect 8436 23078 8504 23134
rect 8560 23078 8628 23134
rect 8684 23078 8752 23134
rect 8808 23078 8876 23134
rect 8932 23078 9000 23134
rect 9056 23078 9124 23134
rect 9180 23078 9248 23134
rect 9304 23078 9372 23134
rect 9428 23078 9496 23134
rect 9552 23078 9620 23134
rect 9676 23078 9744 23134
rect 9800 23078 9810 23134
rect 7874 23010 9810 23078
rect 7874 22954 7884 23010
rect 7940 22954 8008 23010
rect 8064 22954 8132 23010
rect 8188 22954 8256 23010
rect 8312 22954 8380 23010
rect 8436 22954 8504 23010
rect 8560 22954 8628 23010
rect 8684 22954 8752 23010
rect 8808 22954 8876 23010
rect 8932 22954 9000 23010
rect 9056 22954 9124 23010
rect 9180 22954 9248 23010
rect 9304 22954 9372 23010
rect 9428 22954 9496 23010
rect 9552 22954 9620 23010
rect 9676 22954 9744 23010
rect 9800 22954 9810 23010
rect 7874 22886 9810 22954
rect 7874 22830 7884 22886
rect 7940 22830 8008 22886
rect 8064 22830 8132 22886
rect 8188 22830 8256 22886
rect 8312 22830 8380 22886
rect 8436 22830 8504 22886
rect 8560 22830 8628 22886
rect 8684 22830 8752 22886
rect 8808 22830 8876 22886
rect 8932 22830 9000 22886
rect 9056 22830 9124 22886
rect 9180 22830 9248 22886
rect 9304 22830 9372 22886
rect 9428 22830 9496 22886
rect 9552 22830 9620 22886
rect 9676 22830 9744 22886
rect 9800 22830 9810 22886
rect 7874 22762 9810 22830
rect 7874 22706 7884 22762
rect 7940 22706 8008 22762
rect 8064 22706 8132 22762
rect 8188 22706 8256 22762
rect 8312 22706 8380 22762
rect 8436 22706 8504 22762
rect 8560 22706 8628 22762
rect 8684 22706 8752 22762
rect 8808 22706 8876 22762
rect 8932 22706 9000 22762
rect 9056 22706 9124 22762
rect 9180 22706 9248 22762
rect 9304 22706 9372 22762
rect 9428 22706 9496 22762
rect 9552 22706 9620 22762
rect 9676 22706 9744 22762
rect 9800 22706 9810 22762
rect 7874 22638 9810 22706
rect 7874 22582 7884 22638
rect 7940 22582 8008 22638
rect 8064 22582 8132 22638
rect 8188 22582 8256 22638
rect 8312 22582 8380 22638
rect 8436 22582 8504 22638
rect 8560 22582 8628 22638
rect 8684 22582 8752 22638
rect 8808 22582 8876 22638
rect 8932 22582 9000 22638
rect 9056 22582 9124 22638
rect 9180 22582 9248 22638
rect 9304 22582 9372 22638
rect 9428 22582 9496 22638
rect 9552 22582 9620 22638
rect 9676 22582 9744 22638
rect 9800 22582 9810 22638
rect 7874 22514 9810 22582
rect 7874 22458 7884 22514
rect 7940 22458 8008 22514
rect 8064 22458 8132 22514
rect 8188 22458 8256 22514
rect 8312 22458 8380 22514
rect 8436 22458 8504 22514
rect 8560 22458 8628 22514
rect 8684 22458 8752 22514
rect 8808 22458 8876 22514
rect 8932 22458 9000 22514
rect 9056 22458 9124 22514
rect 9180 22458 9248 22514
rect 9304 22458 9372 22514
rect 9428 22458 9496 22514
rect 9552 22458 9620 22514
rect 9676 22458 9744 22514
rect 9800 22458 9810 22514
rect 7874 22390 9810 22458
rect 7874 22334 7884 22390
rect 7940 22334 8008 22390
rect 8064 22334 8132 22390
rect 8188 22334 8256 22390
rect 8312 22334 8380 22390
rect 8436 22334 8504 22390
rect 8560 22334 8628 22390
rect 8684 22334 8752 22390
rect 8808 22334 8876 22390
rect 8932 22334 9000 22390
rect 9056 22334 9124 22390
rect 9180 22334 9248 22390
rect 9304 22334 9372 22390
rect 9428 22334 9496 22390
rect 9552 22334 9620 22390
rect 9676 22334 9744 22390
rect 9800 22334 9810 22390
rect 7874 22266 9810 22334
rect 7874 22210 7884 22266
rect 7940 22210 8008 22266
rect 8064 22210 8132 22266
rect 8188 22210 8256 22266
rect 8312 22210 8380 22266
rect 8436 22210 8504 22266
rect 8560 22210 8628 22266
rect 8684 22210 8752 22266
rect 8808 22210 8876 22266
rect 8932 22210 9000 22266
rect 9056 22210 9124 22266
rect 9180 22210 9248 22266
rect 9304 22210 9372 22266
rect 9428 22210 9496 22266
rect 9552 22210 9620 22266
rect 9676 22210 9744 22266
rect 9800 22210 9810 22266
rect 7874 22142 9810 22210
rect 7874 22086 7884 22142
rect 7940 22086 8008 22142
rect 8064 22086 8132 22142
rect 8188 22086 8256 22142
rect 8312 22086 8380 22142
rect 8436 22086 8504 22142
rect 8560 22086 8628 22142
rect 8684 22086 8752 22142
rect 8808 22086 8876 22142
rect 8932 22086 9000 22142
rect 9056 22086 9124 22142
rect 9180 22086 9248 22142
rect 9304 22086 9372 22142
rect 9428 22086 9496 22142
rect 9552 22086 9620 22142
rect 9676 22086 9744 22142
rect 9800 22086 9810 22142
rect 7874 22018 9810 22086
rect 7874 21962 7884 22018
rect 7940 21962 8008 22018
rect 8064 21962 8132 22018
rect 8188 21962 8256 22018
rect 8312 21962 8380 22018
rect 8436 21962 8504 22018
rect 8560 21962 8628 22018
rect 8684 21962 8752 22018
rect 8808 21962 8876 22018
rect 8932 21962 9000 22018
rect 9056 21962 9124 22018
rect 9180 21962 9248 22018
rect 9304 21962 9372 22018
rect 9428 21962 9496 22018
rect 9552 21962 9620 22018
rect 9676 21962 9744 22018
rect 9800 21962 9810 22018
rect 7874 21894 9810 21962
rect 7874 21838 7884 21894
rect 7940 21838 8008 21894
rect 8064 21838 8132 21894
rect 8188 21838 8256 21894
rect 8312 21838 8380 21894
rect 8436 21838 8504 21894
rect 8560 21838 8628 21894
rect 8684 21838 8752 21894
rect 8808 21838 8876 21894
rect 8932 21838 9000 21894
rect 9056 21838 9124 21894
rect 9180 21838 9248 21894
rect 9304 21838 9372 21894
rect 9428 21838 9496 21894
rect 9552 21838 9620 21894
rect 9676 21838 9744 21894
rect 9800 21838 9810 21894
rect 7874 21770 9810 21838
rect 7874 21714 7884 21770
rect 7940 21714 8008 21770
rect 8064 21714 8132 21770
rect 8188 21714 8256 21770
rect 8312 21714 8380 21770
rect 8436 21714 8504 21770
rect 8560 21714 8628 21770
rect 8684 21714 8752 21770
rect 8808 21714 8876 21770
rect 8932 21714 9000 21770
rect 9056 21714 9124 21770
rect 9180 21714 9248 21770
rect 9304 21714 9372 21770
rect 9428 21714 9496 21770
rect 9552 21714 9620 21770
rect 9676 21714 9744 21770
rect 9800 21714 9810 21770
rect 7874 21646 9810 21714
rect 7874 21590 7884 21646
rect 7940 21590 8008 21646
rect 8064 21590 8132 21646
rect 8188 21590 8256 21646
rect 8312 21590 8380 21646
rect 8436 21590 8504 21646
rect 8560 21590 8628 21646
rect 8684 21590 8752 21646
rect 8808 21590 8876 21646
rect 8932 21590 9000 21646
rect 9056 21590 9124 21646
rect 9180 21590 9248 21646
rect 9304 21590 9372 21646
rect 9428 21590 9496 21646
rect 9552 21590 9620 21646
rect 9676 21590 9744 21646
rect 9800 21590 9810 21646
rect 7874 21522 9810 21590
rect 7874 21466 7884 21522
rect 7940 21466 8008 21522
rect 8064 21466 8132 21522
rect 8188 21466 8256 21522
rect 8312 21466 8380 21522
rect 8436 21466 8504 21522
rect 8560 21466 8628 21522
rect 8684 21466 8752 21522
rect 8808 21466 8876 21522
rect 8932 21466 9000 21522
rect 9056 21466 9124 21522
rect 9180 21466 9248 21522
rect 9304 21466 9372 21522
rect 9428 21466 9496 21522
rect 9552 21466 9620 21522
rect 9676 21466 9744 21522
rect 9800 21466 9810 21522
rect 7874 21398 9810 21466
rect 7874 21342 7884 21398
rect 7940 21342 8008 21398
rect 8064 21342 8132 21398
rect 8188 21342 8256 21398
rect 8312 21342 8380 21398
rect 8436 21342 8504 21398
rect 8560 21342 8628 21398
rect 8684 21342 8752 21398
rect 8808 21342 8876 21398
rect 8932 21342 9000 21398
rect 9056 21342 9124 21398
rect 9180 21342 9248 21398
rect 9304 21342 9372 21398
rect 9428 21342 9496 21398
rect 9552 21342 9620 21398
rect 9676 21342 9744 21398
rect 9800 21342 9810 21398
rect 7874 21274 9810 21342
rect 7874 21218 7884 21274
rect 7940 21218 8008 21274
rect 8064 21218 8132 21274
rect 8188 21218 8256 21274
rect 8312 21218 8380 21274
rect 8436 21218 8504 21274
rect 8560 21218 8628 21274
rect 8684 21218 8752 21274
rect 8808 21218 8876 21274
rect 8932 21218 9000 21274
rect 9056 21218 9124 21274
rect 9180 21218 9248 21274
rect 9304 21218 9372 21274
rect 9428 21218 9496 21274
rect 9552 21218 9620 21274
rect 9676 21218 9744 21274
rect 9800 21218 9810 21274
rect 7874 21150 9810 21218
rect 7874 21094 7884 21150
rect 7940 21094 8008 21150
rect 8064 21094 8132 21150
rect 8188 21094 8256 21150
rect 8312 21094 8380 21150
rect 8436 21094 8504 21150
rect 8560 21094 8628 21150
rect 8684 21094 8752 21150
rect 8808 21094 8876 21150
rect 8932 21094 9000 21150
rect 9056 21094 9124 21150
rect 9180 21094 9248 21150
rect 9304 21094 9372 21150
rect 9428 21094 9496 21150
rect 9552 21094 9620 21150
rect 9676 21094 9744 21150
rect 9800 21094 9810 21150
rect 7874 21026 9810 21094
rect 7874 20970 7884 21026
rect 7940 20970 8008 21026
rect 8064 20970 8132 21026
rect 8188 20970 8256 21026
rect 8312 20970 8380 21026
rect 8436 20970 8504 21026
rect 8560 20970 8628 21026
rect 8684 20970 8752 21026
rect 8808 20970 8876 21026
rect 8932 20970 9000 21026
rect 9056 20970 9124 21026
rect 9180 20970 9248 21026
rect 9304 20970 9372 21026
rect 9428 20970 9496 21026
rect 9552 20970 9620 21026
rect 9676 20970 9744 21026
rect 9800 20970 9810 21026
rect 7874 20902 9810 20970
rect 7874 20846 7884 20902
rect 7940 20846 8008 20902
rect 8064 20846 8132 20902
rect 8188 20846 8256 20902
rect 8312 20846 8380 20902
rect 8436 20846 8504 20902
rect 8560 20846 8628 20902
rect 8684 20846 8752 20902
rect 8808 20846 8876 20902
rect 8932 20846 9000 20902
rect 9056 20846 9124 20902
rect 9180 20846 9248 20902
rect 9304 20846 9372 20902
rect 9428 20846 9496 20902
rect 9552 20846 9620 20902
rect 9676 20846 9744 20902
rect 9800 20846 9810 20902
rect 7874 20836 9810 20846
rect 10244 23754 12180 23764
rect 10244 23698 10254 23754
rect 10310 23698 10378 23754
rect 10434 23698 10502 23754
rect 10558 23698 10626 23754
rect 10682 23698 10750 23754
rect 10806 23698 10874 23754
rect 10930 23698 10998 23754
rect 11054 23698 11122 23754
rect 11178 23698 11246 23754
rect 11302 23698 11370 23754
rect 11426 23698 11494 23754
rect 11550 23698 11618 23754
rect 11674 23698 11742 23754
rect 11798 23698 11866 23754
rect 11922 23698 11990 23754
rect 12046 23698 12114 23754
rect 12170 23698 12180 23754
rect 10244 23630 12180 23698
rect 10244 23574 10254 23630
rect 10310 23574 10378 23630
rect 10434 23574 10502 23630
rect 10558 23574 10626 23630
rect 10682 23574 10750 23630
rect 10806 23574 10874 23630
rect 10930 23574 10998 23630
rect 11054 23574 11122 23630
rect 11178 23574 11246 23630
rect 11302 23574 11370 23630
rect 11426 23574 11494 23630
rect 11550 23574 11618 23630
rect 11674 23574 11742 23630
rect 11798 23574 11866 23630
rect 11922 23574 11990 23630
rect 12046 23574 12114 23630
rect 12170 23574 12180 23630
rect 10244 23506 12180 23574
rect 10244 23450 10254 23506
rect 10310 23450 10378 23506
rect 10434 23450 10502 23506
rect 10558 23450 10626 23506
rect 10682 23450 10750 23506
rect 10806 23450 10874 23506
rect 10930 23450 10998 23506
rect 11054 23450 11122 23506
rect 11178 23450 11246 23506
rect 11302 23450 11370 23506
rect 11426 23450 11494 23506
rect 11550 23450 11618 23506
rect 11674 23450 11742 23506
rect 11798 23450 11866 23506
rect 11922 23450 11990 23506
rect 12046 23450 12114 23506
rect 12170 23450 12180 23506
rect 10244 23382 12180 23450
rect 10244 23326 10254 23382
rect 10310 23326 10378 23382
rect 10434 23326 10502 23382
rect 10558 23326 10626 23382
rect 10682 23326 10750 23382
rect 10806 23326 10874 23382
rect 10930 23326 10998 23382
rect 11054 23326 11122 23382
rect 11178 23326 11246 23382
rect 11302 23326 11370 23382
rect 11426 23326 11494 23382
rect 11550 23326 11618 23382
rect 11674 23326 11742 23382
rect 11798 23326 11866 23382
rect 11922 23326 11990 23382
rect 12046 23326 12114 23382
rect 12170 23326 12180 23382
rect 10244 23258 12180 23326
rect 10244 23202 10254 23258
rect 10310 23202 10378 23258
rect 10434 23202 10502 23258
rect 10558 23202 10626 23258
rect 10682 23202 10750 23258
rect 10806 23202 10874 23258
rect 10930 23202 10998 23258
rect 11054 23202 11122 23258
rect 11178 23202 11246 23258
rect 11302 23202 11370 23258
rect 11426 23202 11494 23258
rect 11550 23202 11618 23258
rect 11674 23202 11742 23258
rect 11798 23202 11866 23258
rect 11922 23202 11990 23258
rect 12046 23202 12114 23258
rect 12170 23202 12180 23258
rect 10244 23134 12180 23202
rect 10244 23078 10254 23134
rect 10310 23078 10378 23134
rect 10434 23078 10502 23134
rect 10558 23078 10626 23134
rect 10682 23078 10750 23134
rect 10806 23078 10874 23134
rect 10930 23078 10998 23134
rect 11054 23078 11122 23134
rect 11178 23078 11246 23134
rect 11302 23078 11370 23134
rect 11426 23078 11494 23134
rect 11550 23078 11618 23134
rect 11674 23078 11742 23134
rect 11798 23078 11866 23134
rect 11922 23078 11990 23134
rect 12046 23078 12114 23134
rect 12170 23078 12180 23134
rect 10244 23010 12180 23078
rect 10244 22954 10254 23010
rect 10310 22954 10378 23010
rect 10434 22954 10502 23010
rect 10558 22954 10626 23010
rect 10682 22954 10750 23010
rect 10806 22954 10874 23010
rect 10930 22954 10998 23010
rect 11054 22954 11122 23010
rect 11178 22954 11246 23010
rect 11302 22954 11370 23010
rect 11426 22954 11494 23010
rect 11550 22954 11618 23010
rect 11674 22954 11742 23010
rect 11798 22954 11866 23010
rect 11922 22954 11990 23010
rect 12046 22954 12114 23010
rect 12170 22954 12180 23010
rect 10244 22886 12180 22954
rect 10244 22830 10254 22886
rect 10310 22830 10378 22886
rect 10434 22830 10502 22886
rect 10558 22830 10626 22886
rect 10682 22830 10750 22886
rect 10806 22830 10874 22886
rect 10930 22830 10998 22886
rect 11054 22830 11122 22886
rect 11178 22830 11246 22886
rect 11302 22830 11370 22886
rect 11426 22830 11494 22886
rect 11550 22830 11618 22886
rect 11674 22830 11742 22886
rect 11798 22830 11866 22886
rect 11922 22830 11990 22886
rect 12046 22830 12114 22886
rect 12170 22830 12180 22886
rect 10244 22762 12180 22830
rect 10244 22706 10254 22762
rect 10310 22706 10378 22762
rect 10434 22706 10502 22762
rect 10558 22706 10626 22762
rect 10682 22706 10750 22762
rect 10806 22706 10874 22762
rect 10930 22706 10998 22762
rect 11054 22706 11122 22762
rect 11178 22706 11246 22762
rect 11302 22706 11370 22762
rect 11426 22706 11494 22762
rect 11550 22706 11618 22762
rect 11674 22706 11742 22762
rect 11798 22706 11866 22762
rect 11922 22706 11990 22762
rect 12046 22706 12114 22762
rect 12170 22706 12180 22762
rect 10244 22638 12180 22706
rect 10244 22582 10254 22638
rect 10310 22582 10378 22638
rect 10434 22582 10502 22638
rect 10558 22582 10626 22638
rect 10682 22582 10750 22638
rect 10806 22582 10874 22638
rect 10930 22582 10998 22638
rect 11054 22582 11122 22638
rect 11178 22582 11246 22638
rect 11302 22582 11370 22638
rect 11426 22582 11494 22638
rect 11550 22582 11618 22638
rect 11674 22582 11742 22638
rect 11798 22582 11866 22638
rect 11922 22582 11990 22638
rect 12046 22582 12114 22638
rect 12170 22582 12180 22638
rect 10244 22514 12180 22582
rect 10244 22458 10254 22514
rect 10310 22458 10378 22514
rect 10434 22458 10502 22514
rect 10558 22458 10626 22514
rect 10682 22458 10750 22514
rect 10806 22458 10874 22514
rect 10930 22458 10998 22514
rect 11054 22458 11122 22514
rect 11178 22458 11246 22514
rect 11302 22458 11370 22514
rect 11426 22458 11494 22514
rect 11550 22458 11618 22514
rect 11674 22458 11742 22514
rect 11798 22458 11866 22514
rect 11922 22458 11990 22514
rect 12046 22458 12114 22514
rect 12170 22458 12180 22514
rect 10244 22390 12180 22458
rect 10244 22334 10254 22390
rect 10310 22334 10378 22390
rect 10434 22334 10502 22390
rect 10558 22334 10626 22390
rect 10682 22334 10750 22390
rect 10806 22334 10874 22390
rect 10930 22334 10998 22390
rect 11054 22334 11122 22390
rect 11178 22334 11246 22390
rect 11302 22334 11370 22390
rect 11426 22334 11494 22390
rect 11550 22334 11618 22390
rect 11674 22334 11742 22390
rect 11798 22334 11866 22390
rect 11922 22334 11990 22390
rect 12046 22334 12114 22390
rect 12170 22334 12180 22390
rect 10244 22266 12180 22334
rect 10244 22210 10254 22266
rect 10310 22210 10378 22266
rect 10434 22210 10502 22266
rect 10558 22210 10626 22266
rect 10682 22210 10750 22266
rect 10806 22210 10874 22266
rect 10930 22210 10998 22266
rect 11054 22210 11122 22266
rect 11178 22210 11246 22266
rect 11302 22210 11370 22266
rect 11426 22210 11494 22266
rect 11550 22210 11618 22266
rect 11674 22210 11742 22266
rect 11798 22210 11866 22266
rect 11922 22210 11990 22266
rect 12046 22210 12114 22266
rect 12170 22210 12180 22266
rect 10244 22142 12180 22210
rect 10244 22086 10254 22142
rect 10310 22086 10378 22142
rect 10434 22086 10502 22142
rect 10558 22086 10626 22142
rect 10682 22086 10750 22142
rect 10806 22086 10874 22142
rect 10930 22086 10998 22142
rect 11054 22086 11122 22142
rect 11178 22086 11246 22142
rect 11302 22086 11370 22142
rect 11426 22086 11494 22142
rect 11550 22086 11618 22142
rect 11674 22086 11742 22142
rect 11798 22086 11866 22142
rect 11922 22086 11990 22142
rect 12046 22086 12114 22142
rect 12170 22086 12180 22142
rect 10244 22018 12180 22086
rect 10244 21962 10254 22018
rect 10310 21962 10378 22018
rect 10434 21962 10502 22018
rect 10558 21962 10626 22018
rect 10682 21962 10750 22018
rect 10806 21962 10874 22018
rect 10930 21962 10998 22018
rect 11054 21962 11122 22018
rect 11178 21962 11246 22018
rect 11302 21962 11370 22018
rect 11426 21962 11494 22018
rect 11550 21962 11618 22018
rect 11674 21962 11742 22018
rect 11798 21962 11866 22018
rect 11922 21962 11990 22018
rect 12046 21962 12114 22018
rect 12170 21962 12180 22018
rect 10244 21894 12180 21962
rect 10244 21838 10254 21894
rect 10310 21838 10378 21894
rect 10434 21838 10502 21894
rect 10558 21838 10626 21894
rect 10682 21838 10750 21894
rect 10806 21838 10874 21894
rect 10930 21838 10998 21894
rect 11054 21838 11122 21894
rect 11178 21838 11246 21894
rect 11302 21838 11370 21894
rect 11426 21838 11494 21894
rect 11550 21838 11618 21894
rect 11674 21838 11742 21894
rect 11798 21838 11866 21894
rect 11922 21838 11990 21894
rect 12046 21838 12114 21894
rect 12170 21838 12180 21894
rect 10244 21770 12180 21838
rect 10244 21714 10254 21770
rect 10310 21714 10378 21770
rect 10434 21714 10502 21770
rect 10558 21714 10626 21770
rect 10682 21714 10750 21770
rect 10806 21714 10874 21770
rect 10930 21714 10998 21770
rect 11054 21714 11122 21770
rect 11178 21714 11246 21770
rect 11302 21714 11370 21770
rect 11426 21714 11494 21770
rect 11550 21714 11618 21770
rect 11674 21714 11742 21770
rect 11798 21714 11866 21770
rect 11922 21714 11990 21770
rect 12046 21714 12114 21770
rect 12170 21714 12180 21770
rect 10244 21646 12180 21714
rect 10244 21590 10254 21646
rect 10310 21590 10378 21646
rect 10434 21590 10502 21646
rect 10558 21590 10626 21646
rect 10682 21590 10750 21646
rect 10806 21590 10874 21646
rect 10930 21590 10998 21646
rect 11054 21590 11122 21646
rect 11178 21590 11246 21646
rect 11302 21590 11370 21646
rect 11426 21590 11494 21646
rect 11550 21590 11618 21646
rect 11674 21590 11742 21646
rect 11798 21590 11866 21646
rect 11922 21590 11990 21646
rect 12046 21590 12114 21646
rect 12170 21590 12180 21646
rect 10244 21522 12180 21590
rect 10244 21466 10254 21522
rect 10310 21466 10378 21522
rect 10434 21466 10502 21522
rect 10558 21466 10626 21522
rect 10682 21466 10750 21522
rect 10806 21466 10874 21522
rect 10930 21466 10998 21522
rect 11054 21466 11122 21522
rect 11178 21466 11246 21522
rect 11302 21466 11370 21522
rect 11426 21466 11494 21522
rect 11550 21466 11618 21522
rect 11674 21466 11742 21522
rect 11798 21466 11866 21522
rect 11922 21466 11990 21522
rect 12046 21466 12114 21522
rect 12170 21466 12180 21522
rect 10244 21398 12180 21466
rect 10244 21342 10254 21398
rect 10310 21342 10378 21398
rect 10434 21342 10502 21398
rect 10558 21342 10626 21398
rect 10682 21342 10750 21398
rect 10806 21342 10874 21398
rect 10930 21342 10998 21398
rect 11054 21342 11122 21398
rect 11178 21342 11246 21398
rect 11302 21342 11370 21398
rect 11426 21342 11494 21398
rect 11550 21342 11618 21398
rect 11674 21342 11742 21398
rect 11798 21342 11866 21398
rect 11922 21342 11990 21398
rect 12046 21342 12114 21398
rect 12170 21342 12180 21398
rect 10244 21274 12180 21342
rect 10244 21218 10254 21274
rect 10310 21218 10378 21274
rect 10434 21218 10502 21274
rect 10558 21218 10626 21274
rect 10682 21218 10750 21274
rect 10806 21218 10874 21274
rect 10930 21218 10998 21274
rect 11054 21218 11122 21274
rect 11178 21218 11246 21274
rect 11302 21218 11370 21274
rect 11426 21218 11494 21274
rect 11550 21218 11618 21274
rect 11674 21218 11742 21274
rect 11798 21218 11866 21274
rect 11922 21218 11990 21274
rect 12046 21218 12114 21274
rect 12170 21218 12180 21274
rect 10244 21150 12180 21218
rect 10244 21094 10254 21150
rect 10310 21094 10378 21150
rect 10434 21094 10502 21150
rect 10558 21094 10626 21150
rect 10682 21094 10750 21150
rect 10806 21094 10874 21150
rect 10930 21094 10998 21150
rect 11054 21094 11122 21150
rect 11178 21094 11246 21150
rect 11302 21094 11370 21150
rect 11426 21094 11494 21150
rect 11550 21094 11618 21150
rect 11674 21094 11742 21150
rect 11798 21094 11866 21150
rect 11922 21094 11990 21150
rect 12046 21094 12114 21150
rect 12170 21094 12180 21150
rect 10244 21026 12180 21094
rect 10244 20970 10254 21026
rect 10310 20970 10378 21026
rect 10434 20970 10502 21026
rect 10558 20970 10626 21026
rect 10682 20970 10750 21026
rect 10806 20970 10874 21026
rect 10930 20970 10998 21026
rect 11054 20970 11122 21026
rect 11178 20970 11246 21026
rect 11302 20970 11370 21026
rect 11426 20970 11494 21026
rect 11550 20970 11618 21026
rect 11674 20970 11742 21026
rect 11798 20970 11866 21026
rect 11922 20970 11990 21026
rect 12046 20970 12114 21026
rect 12170 20970 12180 21026
rect 10244 20902 12180 20970
rect 10244 20846 10254 20902
rect 10310 20846 10378 20902
rect 10434 20846 10502 20902
rect 10558 20846 10626 20902
rect 10682 20846 10750 20902
rect 10806 20846 10874 20902
rect 10930 20846 10998 20902
rect 11054 20846 11122 20902
rect 11178 20846 11246 20902
rect 11302 20846 11370 20902
rect 11426 20846 11494 20902
rect 11550 20846 11618 20902
rect 11674 20846 11742 20902
rect 11798 20846 11866 20902
rect 11922 20846 11990 20902
rect 12046 20846 12114 20902
rect 12170 20846 12180 20902
rect 10244 20836 12180 20846
rect 12861 23754 14673 23764
rect 12861 23698 12871 23754
rect 12927 23698 12995 23754
rect 13051 23698 13119 23754
rect 13175 23698 13243 23754
rect 13299 23698 13367 23754
rect 13423 23698 13491 23754
rect 13547 23698 13615 23754
rect 13671 23698 13739 23754
rect 13795 23698 13863 23754
rect 13919 23698 13987 23754
rect 14043 23698 14111 23754
rect 14167 23698 14235 23754
rect 14291 23698 14359 23754
rect 14415 23698 14483 23754
rect 14539 23698 14607 23754
rect 14663 23698 14673 23754
rect 12861 23630 14673 23698
rect 12861 23574 12871 23630
rect 12927 23574 12995 23630
rect 13051 23574 13119 23630
rect 13175 23574 13243 23630
rect 13299 23574 13367 23630
rect 13423 23574 13491 23630
rect 13547 23574 13615 23630
rect 13671 23574 13739 23630
rect 13795 23574 13863 23630
rect 13919 23574 13987 23630
rect 14043 23574 14111 23630
rect 14167 23574 14235 23630
rect 14291 23574 14359 23630
rect 14415 23574 14483 23630
rect 14539 23574 14607 23630
rect 14663 23574 14673 23630
rect 12861 23506 14673 23574
rect 12861 23450 12871 23506
rect 12927 23450 12995 23506
rect 13051 23450 13119 23506
rect 13175 23450 13243 23506
rect 13299 23450 13367 23506
rect 13423 23450 13491 23506
rect 13547 23450 13615 23506
rect 13671 23450 13739 23506
rect 13795 23450 13863 23506
rect 13919 23450 13987 23506
rect 14043 23450 14111 23506
rect 14167 23450 14235 23506
rect 14291 23450 14359 23506
rect 14415 23450 14483 23506
rect 14539 23450 14607 23506
rect 14663 23450 14673 23506
rect 12861 23382 14673 23450
rect 12861 23326 12871 23382
rect 12927 23326 12995 23382
rect 13051 23326 13119 23382
rect 13175 23326 13243 23382
rect 13299 23326 13367 23382
rect 13423 23326 13491 23382
rect 13547 23326 13615 23382
rect 13671 23326 13739 23382
rect 13795 23326 13863 23382
rect 13919 23326 13987 23382
rect 14043 23326 14111 23382
rect 14167 23326 14235 23382
rect 14291 23326 14359 23382
rect 14415 23326 14483 23382
rect 14539 23326 14607 23382
rect 14663 23326 14673 23382
rect 12861 23258 14673 23326
rect 12861 23202 12871 23258
rect 12927 23202 12995 23258
rect 13051 23202 13119 23258
rect 13175 23202 13243 23258
rect 13299 23202 13367 23258
rect 13423 23202 13491 23258
rect 13547 23202 13615 23258
rect 13671 23202 13739 23258
rect 13795 23202 13863 23258
rect 13919 23202 13987 23258
rect 14043 23202 14111 23258
rect 14167 23202 14235 23258
rect 14291 23202 14359 23258
rect 14415 23202 14483 23258
rect 14539 23202 14607 23258
rect 14663 23202 14673 23258
rect 12861 23134 14673 23202
rect 12861 23078 12871 23134
rect 12927 23078 12995 23134
rect 13051 23078 13119 23134
rect 13175 23078 13243 23134
rect 13299 23078 13367 23134
rect 13423 23078 13491 23134
rect 13547 23078 13615 23134
rect 13671 23078 13739 23134
rect 13795 23078 13863 23134
rect 13919 23078 13987 23134
rect 14043 23078 14111 23134
rect 14167 23078 14235 23134
rect 14291 23078 14359 23134
rect 14415 23078 14483 23134
rect 14539 23078 14607 23134
rect 14663 23078 14673 23134
rect 12861 23010 14673 23078
rect 12861 22954 12871 23010
rect 12927 22954 12995 23010
rect 13051 22954 13119 23010
rect 13175 22954 13243 23010
rect 13299 22954 13367 23010
rect 13423 22954 13491 23010
rect 13547 22954 13615 23010
rect 13671 22954 13739 23010
rect 13795 22954 13863 23010
rect 13919 22954 13987 23010
rect 14043 22954 14111 23010
rect 14167 22954 14235 23010
rect 14291 22954 14359 23010
rect 14415 22954 14483 23010
rect 14539 22954 14607 23010
rect 14663 22954 14673 23010
rect 12861 22886 14673 22954
rect 12861 22830 12871 22886
rect 12927 22830 12995 22886
rect 13051 22830 13119 22886
rect 13175 22830 13243 22886
rect 13299 22830 13367 22886
rect 13423 22830 13491 22886
rect 13547 22830 13615 22886
rect 13671 22830 13739 22886
rect 13795 22830 13863 22886
rect 13919 22830 13987 22886
rect 14043 22830 14111 22886
rect 14167 22830 14235 22886
rect 14291 22830 14359 22886
rect 14415 22830 14483 22886
rect 14539 22830 14607 22886
rect 14663 22830 14673 22886
rect 12861 22762 14673 22830
rect 12861 22706 12871 22762
rect 12927 22706 12995 22762
rect 13051 22706 13119 22762
rect 13175 22706 13243 22762
rect 13299 22706 13367 22762
rect 13423 22706 13491 22762
rect 13547 22706 13615 22762
rect 13671 22706 13739 22762
rect 13795 22706 13863 22762
rect 13919 22706 13987 22762
rect 14043 22706 14111 22762
rect 14167 22706 14235 22762
rect 14291 22706 14359 22762
rect 14415 22706 14483 22762
rect 14539 22706 14607 22762
rect 14663 22706 14673 22762
rect 12861 22638 14673 22706
rect 12861 22582 12871 22638
rect 12927 22582 12995 22638
rect 13051 22582 13119 22638
rect 13175 22582 13243 22638
rect 13299 22582 13367 22638
rect 13423 22582 13491 22638
rect 13547 22582 13615 22638
rect 13671 22582 13739 22638
rect 13795 22582 13863 22638
rect 13919 22582 13987 22638
rect 14043 22582 14111 22638
rect 14167 22582 14235 22638
rect 14291 22582 14359 22638
rect 14415 22582 14483 22638
rect 14539 22582 14607 22638
rect 14663 22582 14673 22638
rect 12861 22514 14673 22582
rect 12861 22458 12871 22514
rect 12927 22458 12995 22514
rect 13051 22458 13119 22514
rect 13175 22458 13243 22514
rect 13299 22458 13367 22514
rect 13423 22458 13491 22514
rect 13547 22458 13615 22514
rect 13671 22458 13739 22514
rect 13795 22458 13863 22514
rect 13919 22458 13987 22514
rect 14043 22458 14111 22514
rect 14167 22458 14235 22514
rect 14291 22458 14359 22514
rect 14415 22458 14483 22514
rect 14539 22458 14607 22514
rect 14663 22458 14673 22514
rect 12861 22390 14673 22458
rect 12861 22334 12871 22390
rect 12927 22334 12995 22390
rect 13051 22334 13119 22390
rect 13175 22334 13243 22390
rect 13299 22334 13367 22390
rect 13423 22334 13491 22390
rect 13547 22334 13615 22390
rect 13671 22334 13739 22390
rect 13795 22334 13863 22390
rect 13919 22334 13987 22390
rect 14043 22334 14111 22390
rect 14167 22334 14235 22390
rect 14291 22334 14359 22390
rect 14415 22334 14483 22390
rect 14539 22334 14607 22390
rect 14663 22334 14673 22390
rect 12861 22266 14673 22334
rect 12861 22210 12871 22266
rect 12927 22210 12995 22266
rect 13051 22210 13119 22266
rect 13175 22210 13243 22266
rect 13299 22210 13367 22266
rect 13423 22210 13491 22266
rect 13547 22210 13615 22266
rect 13671 22210 13739 22266
rect 13795 22210 13863 22266
rect 13919 22210 13987 22266
rect 14043 22210 14111 22266
rect 14167 22210 14235 22266
rect 14291 22210 14359 22266
rect 14415 22210 14483 22266
rect 14539 22210 14607 22266
rect 14663 22210 14673 22266
rect 12861 22142 14673 22210
rect 12861 22086 12871 22142
rect 12927 22086 12995 22142
rect 13051 22086 13119 22142
rect 13175 22086 13243 22142
rect 13299 22086 13367 22142
rect 13423 22086 13491 22142
rect 13547 22086 13615 22142
rect 13671 22086 13739 22142
rect 13795 22086 13863 22142
rect 13919 22086 13987 22142
rect 14043 22086 14111 22142
rect 14167 22086 14235 22142
rect 14291 22086 14359 22142
rect 14415 22086 14483 22142
rect 14539 22086 14607 22142
rect 14663 22086 14673 22142
rect 12861 22018 14673 22086
rect 12861 21962 12871 22018
rect 12927 21962 12995 22018
rect 13051 21962 13119 22018
rect 13175 21962 13243 22018
rect 13299 21962 13367 22018
rect 13423 21962 13491 22018
rect 13547 21962 13615 22018
rect 13671 21962 13739 22018
rect 13795 21962 13863 22018
rect 13919 21962 13987 22018
rect 14043 21962 14111 22018
rect 14167 21962 14235 22018
rect 14291 21962 14359 22018
rect 14415 21962 14483 22018
rect 14539 21962 14607 22018
rect 14663 21962 14673 22018
rect 12861 21894 14673 21962
rect 12861 21838 12871 21894
rect 12927 21838 12995 21894
rect 13051 21838 13119 21894
rect 13175 21838 13243 21894
rect 13299 21838 13367 21894
rect 13423 21838 13491 21894
rect 13547 21838 13615 21894
rect 13671 21838 13739 21894
rect 13795 21838 13863 21894
rect 13919 21838 13987 21894
rect 14043 21838 14111 21894
rect 14167 21838 14235 21894
rect 14291 21838 14359 21894
rect 14415 21838 14483 21894
rect 14539 21838 14607 21894
rect 14663 21838 14673 21894
rect 12861 21770 14673 21838
rect 12861 21714 12871 21770
rect 12927 21714 12995 21770
rect 13051 21714 13119 21770
rect 13175 21714 13243 21770
rect 13299 21714 13367 21770
rect 13423 21714 13491 21770
rect 13547 21714 13615 21770
rect 13671 21714 13739 21770
rect 13795 21714 13863 21770
rect 13919 21714 13987 21770
rect 14043 21714 14111 21770
rect 14167 21714 14235 21770
rect 14291 21714 14359 21770
rect 14415 21714 14483 21770
rect 14539 21714 14607 21770
rect 14663 21714 14673 21770
rect 12861 21646 14673 21714
rect 12861 21590 12871 21646
rect 12927 21590 12995 21646
rect 13051 21590 13119 21646
rect 13175 21590 13243 21646
rect 13299 21590 13367 21646
rect 13423 21590 13491 21646
rect 13547 21590 13615 21646
rect 13671 21590 13739 21646
rect 13795 21590 13863 21646
rect 13919 21590 13987 21646
rect 14043 21590 14111 21646
rect 14167 21590 14235 21646
rect 14291 21590 14359 21646
rect 14415 21590 14483 21646
rect 14539 21590 14607 21646
rect 14663 21590 14673 21646
rect 12861 21522 14673 21590
rect 12861 21466 12871 21522
rect 12927 21466 12995 21522
rect 13051 21466 13119 21522
rect 13175 21466 13243 21522
rect 13299 21466 13367 21522
rect 13423 21466 13491 21522
rect 13547 21466 13615 21522
rect 13671 21466 13739 21522
rect 13795 21466 13863 21522
rect 13919 21466 13987 21522
rect 14043 21466 14111 21522
rect 14167 21466 14235 21522
rect 14291 21466 14359 21522
rect 14415 21466 14483 21522
rect 14539 21466 14607 21522
rect 14663 21466 14673 21522
rect 12861 21398 14673 21466
rect 12861 21342 12871 21398
rect 12927 21342 12995 21398
rect 13051 21342 13119 21398
rect 13175 21342 13243 21398
rect 13299 21342 13367 21398
rect 13423 21342 13491 21398
rect 13547 21342 13615 21398
rect 13671 21342 13739 21398
rect 13795 21342 13863 21398
rect 13919 21342 13987 21398
rect 14043 21342 14111 21398
rect 14167 21342 14235 21398
rect 14291 21342 14359 21398
rect 14415 21342 14483 21398
rect 14539 21342 14607 21398
rect 14663 21342 14673 21398
rect 12861 21274 14673 21342
rect 12861 21218 12871 21274
rect 12927 21218 12995 21274
rect 13051 21218 13119 21274
rect 13175 21218 13243 21274
rect 13299 21218 13367 21274
rect 13423 21218 13491 21274
rect 13547 21218 13615 21274
rect 13671 21218 13739 21274
rect 13795 21218 13863 21274
rect 13919 21218 13987 21274
rect 14043 21218 14111 21274
rect 14167 21218 14235 21274
rect 14291 21218 14359 21274
rect 14415 21218 14483 21274
rect 14539 21218 14607 21274
rect 14663 21218 14673 21274
rect 12861 21150 14673 21218
rect 12861 21094 12871 21150
rect 12927 21094 12995 21150
rect 13051 21094 13119 21150
rect 13175 21094 13243 21150
rect 13299 21094 13367 21150
rect 13423 21094 13491 21150
rect 13547 21094 13615 21150
rect 13671 21094 13739 21150
rect 13795 21094 13863 21150
rect 13919 21094 13987 21150
rect 14043 21094 14111 21150
rect 14167 21094 14235 21150
rect 14291 21094 14359 21150
rect 14415 21094 14483 21150
rect 14539 21094 14607 21150
rect 14663 21094 14673 21150
rect 12861 21026 14673 21094
rect 12861 20970 12871 21026
rect 12927 20970 12995 21026
rect 13051 20970 13119 21026
rect 13175 20970 13243 21026
rect 13299 20970 13367 21026
rect 13423 20970 13491 21026
rect 13547 20970 13615 21026
rect 13671 20970 13739 21026
rect 13795 20970 13863 21026
rect 13919 20970 13987 21026
rect 14043 20970 14111 21026
rect 14167 20970 14235 21026
rect 14291 20970 14359 21026
rect 14415 20970 14483 21026
rect 14539 20970 14607 21026
rect 14663 20970 14673 21026
rect 12861 20902 14673 20970
rect 12861 20846 12871 20902
rect 12927 20846 12995 20902
rect 13051 20846 13119 20902
rect 13175 20846 13243 20902
rect 13299 20846 13367 20902
rect 13423 20846 13491 20902
rect 13547 20846 13615 20902
rect 13671 20846 13739 20902
rect 13795 20846 13863 20902
rect 13919 20846 13987 20902
rect 14043 20846 14111 20902
rect 14167 20846 14235 20902
rect 14291 20846 14359 20902
rect 14415 20846 14483 20902
rect 14539 20846 14607 20902
rect 14663 20846 14673 20902
rect 12861 20836 14673 20846
rect 305 20554 2117 20564
rect 305 20498 315 20554
rect 371 20498 439 20554
rect 495 20498 563 20554
rect 619 20498 687 20554
rect 743 20498 811 20554
rect 867 20498 935 20554
rect 991 20498 1059 20554
rect 1115 20498 1183 20554
rect 1239 20498 1307 20554
rect 1363 20498 1431 20554
rect 1487 20498 1555 20554
rect 1611 20498 1679 20554
rect 1735 20498 1803 20554
rect 1859 20498 1927 20554
rect 1983 20498 2051 20554
rect 2107 20498 2117 20554
rect 305 20430 2117 20498
rect 305 20374 315 20430
rect 371 20374 439 20430
rect 495 20374 563 20430
rect 619 20374 687 20430
rect 743 20374 811 20430
rect 867 20374 935 20430
rect 991 20374 1059 20430
rect 1115 20374 1183 20430
rect 1239 20374 1307 20430
rect 1363 20374 1431 20430
rect 1487 20374 1555 20430
rect 1611 20374 1679 20430
rect 1735 20374 1803 20430
rect 1859 20374 1927 20430
rect 1983 20374 2051 20430
rect 2107 20374 2117 20430
rect 305 20306 2117 20374
rect 305 20250 315 20306
rect 371 20250 439 20306
rect 495 20250 563 20306
rect 619 20250 687 20306
rect 743 20250 811 20306
rect 867 20250 935 20306
rect 991 20250 1059 20306
rect 1115 20250 1183 20306
rect 1239 20250 1307 20306
rect 1363 20250 1431 20306
rect 1487 20250 1555 20306
rect 1611 20250 1679 20306
rect 1735 20250 1803 20306
rect 1859 20250 1927 20306
rect 1983 20250 2051 20306
rect 2107 20250 2117 20306
rect 305 20182 2117 20250
rect 305 20126 315 20182
rect 371 20126 439 20182
rect 495 20126 563 20182
rect 619 20126 687 20182
rect 743 20126 811 20182
rect 867 20126 935 20182
rect 991 20126 1059 20182
rect 1115 20126 1183 20182
rect 1239 20126 1307 20182
rect 1363 20126 1431 20182
rect 1487 20126 1555 20182
rect 1611 20126 1679 20182
rect 1735 20126 1803 20182
rect 1859 20126 1927 20182
rect 1983 20126 2051 20182
rect 2107 20126 2117 20182
rect 305 20058 2117 20126
rect 305 20002 315 20058
rect 371 20002 439 20058
rect 495 20002 563 20058
rect 619 20002 687 20058
rect 743 20002 811 20058
rect 867 20002 935 20058
rect 991 20002 1059 20058
rect 1115 20002 1183 20058
rect 1239 20002 1307 20058
rect 1363 20002 1431 20058
rect 1487 20002 1555 20058
rect 1611 20002 1679 20058
rect 1735 20002 1803 20058
rect 1859 20002 1927 20058
rect 1983 20002 2051 20058
rect 2107 20002 2117 20058
rect 305 19934 2117 20002
rect 305 19878 315 19934
rect 371 19878 439 19934
rect 495 19878 563 19934
rect 619 19878 687 19934
rect 743 19878 811 19934
rect 867 19878 935 19934
rect 991 19878 1059 19934
rect 1115 19878 1183 19934
rect 1239 19878 1307 19934
rect 1363 19878 1431 19934
rect 1487 19878 1555 19934
rect 1611 19878 1679 19934
rect 1735 19878 1803 19934
rect 1859 19878 1927 19934
rect 1983 19878 2051 19934
rect 2107 19878 2117 19934
rect 305 19810 2117 19878
rect 305 19754 315 19810
rect 371 19754 439 19810
rect 495 19754 563 19810
rect 619 19754 687 19810
rect 743 19754 811 19810
rect 867 19754 935 19810
rect 991 19754 1059 19810
rect 1115 19754 1183 19810
rect 1239 19754 1307 19810
rect 1363 19754 1431 19810
rect 1487 19754 1555 19810
rect 1611 19754 1679 19810
rect 1735 19754 1803 19810
rect 1859 19754 1927 19810
rect 1983 19754 2051 19810
rect 2107 19754 2117 19810
rect 305 19686 2117 19754
rect 305 19630 315 19686
rect 371 19630 439 19686
rect 495 19630 563 19686
rect 619 19630 687 19686
rect 743 19630 811 19686
rect 867 19630 935 19686
rect 991 19630 1059 19686
rect 1115 19630 1183 19686
rect 1239 19630 1307 19686
rect 1363 19630 1431 19686
rect 1487 19630 1555 19686
rect 1611 19630 1679 19686
rect 1735 19630 1803 19686
rect 1859 19630 1927 19686
rect 1983 19630 2051 19686
rect 2107 19630 2117 19686
rect 305 19562 2117 19630
rect 305 19506 315 19562
rect 371 19506 439 19562
rect 495 19506 563 19562
rect 619 19506 687 19562
rect 743 19506 811 19562
rect 867 19506 935 19562
rect 991 19506 1059 19562
rect 1115 19506 1183 19562
rect 1239 19506 1307 19562
rect 1363 19506 1431 19562
rect 1487 19506 1555 19562
rect 1611 19506 1679 19562
rect 1735 19506 1803 19562
rect 1859 19506 1927 19562
rect 1983 19506 2051 19562
rect 2107 19506 2117 19562
rect 305 19438 2117 19506
rect 305 19382 315 19438
rect 371 19382 439 19438
rect 495 19382 563 19438
rect 619 19382 687 19438
rect 743 19382 811 19438
rect 867 19382 935 19438
rect 991 19382 1059 19438
rect 1115 19382 1183 19438
rect 1239 19382 1307 19438
rect 1363 19382 1431 19438
rect 1487 19382 1555 19438
rect 1611 19382 1679 19438
rect 1735 19382 1803 19438
rect 1859 19382 1927 19438
rect 1983 19382 2051 19438
rect 2107 19382 2117 19438
rect 305 19314 2117 19382
rect 305 19258 315 19314
rect 371 19258 439 19314
rect 495 19258 563 19314
rect 619 19258 687 19314
rect 743 19258 811 19314
rect 867 19258 935 19314
rect 991 19258 1059 19314
rect 1115 19258 1183 19314
rect 1239 19258 1307 19314
rect 1363 19258 1431 19314
rect 1487 19258 1555 19314
rect 1611 19258 1679 19314
rect 1735 19258 1803 19314
rect 1859 19258 1927 19314
rect 1983 19258 2051 19314
rect 2107 19258 2117 19314
rect 305 19190 2117 19258
rect 305 19134 315 19190
rect 371 19134 439 19190
rect 495 19134 563 19190
rect 619 19134 687 19190
rect 743 19134 811 19190
rect 867 19134 935 19190
rect 991 19134 1059 19190
rect 1115 19134 1183 19190
rect 1239 19134 1307 19190
rect 1363 19134 1431 19190
rect 1487 19134 1555 19190
rect 1611 19134 1679 19190
rect 1735 19134 1803 19190
rect 1859 19134 1927 19190
rect 1983 19134 2051 19190
rect 2107 19134 2117 19190
rect 305 19066 2117 19134
rect 305 19010 315 19066
rect 371 19010 439 19066
rect 495 19010 563 19066
rect 619 19010 687 19066
rect 743 19010 811 19066
rect 867 19010 935 19066
rect 991 19010 1059 19066
rect 1115 19010 1183 19066
rect 1239 19010 1307 19066
rect 1363 19010 1431 19066
rect 1487 19010 1555 19066
rect 1611 19010 1679 19066
rect 1735 19010 1803 19066
rect 1859 19010 1927 19066
rect 1983 19010 2051 19066
rect 2107 19010 2117 19066
rect 305 18942 2117 19010
rect 305 18886 315 18942
rect 371 18886 439 18942
rect 495 18886 563 18942
rect 619 18886 687 18942
rect 743 18886 811 18942
rect 867 18886 935 18942
rect 991 18886 1059 18942
rect 1115 18886 1183 18942
rect 1239 18886 1307 18942
rect 1363 18886 1431 18942
rect 1487 18886 1555 18942
rect 1611 18886 1679 18942
rect 1735 18886 1803 18942
rect 1859 18886 1927 18942
rect 1983 18886 2051 18942
rect 2107 18886 2117 18942
rect 305 18818 2117 18886
rect 305 18762 315 18818
rect 371 18762 439 18818
rect 495 18762 563 18818
rect 619 18762 687 18818
rect 743 18762 811 18818
rect 867 18762 935 18818
rect 991 18762 1059 18818
rect 1115 18762 1183 18818
rect 1239 18762 1307 18818
rect 1363 18762 1431 18818
rect 1487 18762 1555 18818
rect 1611 18762 1679 18818
rect 1735 18762 1803 18818
rect 1859 18762 1927 18818
rect 1983 18762 2051 18818
rect 2107 18762 2117 18818
rect 305 18694 2117 18762
rect 305 18638 315 18694
rect 371 18638 439 18694
rect 495 18638 563 18694
rect 619 18638 687 18694
rect 743 18638 811 18694
rect 867 18638 935 18694
rect 991 18638 1059 18694
rect 1115 18638 1183 18694
rect 1239 18638 1307 18694
rect 1363 18638 1431 18694
rect 1487 18638 1555 18694
rect 1611 18638 1679 18694
rect 1735 18638 1803 18694
rect 1859 18638 1927 18694
rect 1983 18638 2051 18694
rect 2107 18638 2117 18694
rect 305 18570 2117 18638
rect 305 18514 315 18570
rect 371 18514 439 18570
rect 495 18514 563 18570
rect 619 18514 687 18570
rect 743 18514 811 18570
rect 867 18514 935 18570
rect 991 18514 1059 18570
rect 1115 18514 1183 18570
rect 1239 18514 1307 18570
rect 1363 18514 1431 18570
rect 1487 18514 1555 18570
rect 1611 18514 1679 18570
rect 1735 18514 1803 18570
rect 1859 18514 1927 18570
rect 1983 18514 2051 18570
rect 2107 18514 2117 18570
rect 305 18446 2117 18514
rect 305 18390 315 18446
rect 371 18390 439 18446
rect 495 18390 563 18446
rect 619 18390 687 18446
rect 743 18390 811 18446
rect 867 18390 935 18446
rect 991 18390 1059 18446
rect 1115 18390 1183 18446
rect 1239 18390 1307 18446
rect 1363 18390 1431 18446
rect 1487 18390 1555 18446
rect 1611 18390 1679 18446
rect 1735 18390 1803 18446
rect 1859 18390 1927 18446
rect 1983 18390 2051 18446
rect 2107 18390 2117 18446
rect 305 18322 2117 18390
rect 305 18266 315 18322
rect 371 18266 439 18322
rect 495 18266 563 18322
rect 619 18266 687 18322
rect 743 18266 811 18322
rect 867 18266 935 18322
rect 991 18266 1059 18322
rect 1115 18266 1183 18322
rect 1239 18266 1307 18322
rect 1363 18266 1431 18322
rect 1487 18266 1555 18322
rect 1611 18266 1679 18322
rect 1735 18266 1803 18322
rect 1859 18266 1927 18322
rect 1983 18266 2051 18322
rect 2107 18266 2117 18322
rect 305 18198 2117 18266
rect 305 18142 315 18198
rect 371 18142 439 18198
rect 495 18142 563 18198
rect 619 18142 687 18198
rect 743 18142 811 18198
rect 867 18142 935 18198
rect 991 18142 1059 18198
rect 1115 18142 1183 18198
rect 1239 18142 1307 18198
rect 1363 18142 1431 18198
rect 1487 18142 1555 18198
rect 1611 18142 1679 18198
rect 1735 18142 1803 18198
rect 1859 18142 1927 18198
rect 1983 18142 2051 18198
rect 2107 18142 2117 18198
rect 305 18074 2117 18142
rect 305 18018 315 18074
rect 371 18018 439 18074
rect 495 18018 563 18074
rect 619 18018 687 18074
rect 743 18018 811 18074
rect 867 18018 935 18074
rect 991 18018 1059 18074
rect 1115 18018 1183 18074
rect 1239 18018 1307 18074
rect 1363 18018 1431 18074
rect 1487 18018 1555 18074
rect 1611 18018 1679 18074
rect 1735 18018 1803 18074
rect 1859 18018 1927 18074
rect 1983 18018 2051 18074
rect 2107 18018 2117 18074
rect 305 17950 2117 18018
rect 305 17894 315 17950
rect 371 17894 439 17950
rect 495 17894 563 17950
rect 619 17894 687 17950
rect 743 17894 811 17950
rect 867 17894 935 17950
rect 991 17894 1059 17950
rect 1115 17894 1183 17950
rect 1239 17894 1307 17950
rect 1363 17894 1431 17950
rect 1487 17894 1555 17950
rect 1611 17894 1679 17950
rect 1735 17894 1803 17950
rect 1859 17894 1927 17950
rect 1983 17894 2051 17950
rect 2107 17894 2117 17950
rect 305 17826 2117 17894
rect 305 17770 315 17826
rect 371 17770 439 17826
rect 495 17770 563 17826
rect 619 17770 687 17826
rect 743 17770 811 17826
rect 867 17770 935 17826
rect 991 17770 1059 17826
rect 1115 17770 1183 17826
rect 1239 17770 1307 17826
rect 1363 17770 1431 17826
rect 1487 17770 1555 17826
rect 1611 17770 1679 17826
rect 1735 17770 1803 17826
rect 1859 17770 1927 17826
rect 1983 17770 2051 17826
rect 2107 17770 2117 17826
rect 305 17702 2117 17770
rect 305 17646 315 17702
rect 371 17646 439 17702
rect 495 17646 563 17702
rect 619 17646 687 17702
rect 743 17646 811 17702
rect 867 17646 935 17702
rect 991 17646 1059 17702
rect 1115 17646 1183 17702
rect 1239 17646 1307 17702
rect 1363 17646 1431 17702
rect 1487 17646 1555 17702
rect 1611 17646 1679 17702
rect 1735 17646 1803 17702
rect 1859 17646 1927 17702
rect 1983 17646 2051 17702
rect 2107 17646 2117 17702
rect 305 17636 2117 17646
rect 2798 20554 4734 20564
rect 2798 20498 2808 20554
rect 2864 20498 2932 20554
rect 2988 20498 3056 20554
rect 3112 20498 3180 20554
rect 3236 20498 3304 20554
rect 3360 20498 3428 20554
rect 3484 20498 3552 20554
rect 3608 20498 3676 20554
rect 3732 20498 3800 20554
rect 3856 20498 3924 20554
rect 3980 20498 4048 20554
rect 4104 20498 4172 20554
rect 4228 20498 4296 20554
rect 4352 20498 4420 20554
rect 4476 20498 4544 20554
rect 4600 20498 4668 20554
rect 4724 20498 4734 20554
rect 2798 20430 4734 20498
rect 2798 20374 2808 20430
rect 2864 20374 2932 20430
rect 2988 20374 3056 20430
rect 3112 20374 3180 20430
rect 3236 20374 3304 20430
rect 3360 20374 3428 20430
rect 3484 20374 3552 20430
rect 3608 20374 3676 20430
rect 3732 20374 3800 20430
rect 3856 20374 3924 20430
rect 3980 20374 4048 20430
rect 4104 20374 4172 20430
rect 4228 20374 4296 20430
rect 4352 20374 4420 20430
rect 4476 20374 4544 20430
rect 4600 20374 4668 20430
rect 4724 20374 4734 20430
rect 2798 20306 4734 20374
rect 2798 20250 2808 20306
rect 2864 20250 2932 20306
rect 2988 20250 3056 20306
rect 3112 20250 3180 20306
rect 3236 20250 3304 20306
rect 3360 20250 3428 20306
rect 3484 20250 3552 20306
rect 3608 20250 3676 20306
rect 3732 20250 3800 20306
rect 3856 20250 3924 20306
rect 3980 20250 4048 20306
rect 4104 20250 4172 20306
rect 4228 20250 4296 20306
rect 4352 20250 4420 20306
rect 4476 20250 4544 20306
rect 4600 20250 4668 20306
rect 4724 20250 4734 20306
rect 2798 20182 4734 20250
rect 2798 20126 2808 20182
rect 2864 20126 2932 20182
rect 2988 20126 3056 20182
rect 3112 20126 3180 20182
rect 3236 20126 3304 20182
rect 3360 20126 3428 20182
rect 3484 20126 3552 20182
rect 3608 20126 3676 20182
rect 3732 20126 3800 20182
rect 3856 20126 3924 20182
rect 3980 20126 4048 20182
rect 4104 20126 4172 20182
rect 4228 20126 4296 20182
rect 4352 20126 4420 20182
rect 4476 20126 4544 20182
rect 4600 20126 4668 20182
rect 4724 20126 4734 20182
rect 2798 20058 4734 20126
rect 2798 20002 2808 20058
rect 2864 20002 2932 20058
rect 2988 20002 3056 20058
rect 3112 20002 3180 20058
rect 3236 20002 3304 20058
rect 3360 20002 3428 20058
rect 3484 20002 3552 20058
rect 3608 20002 3676 20058
rect 3732 20002 3800 20058
rect 3856 20002 3924 20058
rect 3980 20002 4048 20058
rect 4104 20002 4172 20058
rect 4228 20002 4296 20058
rect 4352 20002 4420 20058
rect 4476 20002 4544 20058
rect 4600 20002 4668 20058
rect 4724 20002 4734 20058
rect 2798 19934 4734 20002
rect 2798 19878 2808 19934
rect 2864 19878 2932 19934
rect 2988 19878 3056 19934
rect 3112 19878 3180 19934
rect 3236 19878 3304 19934
rect 3360 19878 3428 19934
rect 3484 19878 3552 19934
rect 3608 19878 3676 19934
rect 3732 19878 3800 19934
rect 3856 19878 3924 19934
rect 3980 19878 4048 19934
rect 4104 19878 4172 19934
rect 4228 19878 4296 19934
rect 4352 19878 4420 19934
rect 4476 19878 4544 19934
rect 4600 19878 4668 19934
rect 4724 19878 4734 19934
rect 2798 19810 4734 19878
rect 2798 19754 2808 19810
rect 2864 19754 2932 19810
rect 2988 19754 3056 19810
rect 3112 19754 3180 19810
rect 3236 19754 3304 19810
rect 3360 19754 3428 19810
rect 3484 19754 3552 19810
rect 3608 19754 3676 19810
rect 3732 19754 3800 19810
rect 3856 19754 3924 19810
rect 3980 19754 4048 19810
rect 4104 19754 4172 19810
rect 4228 19754 4296 19810
rect 4352 19754 4420 19810
rect 4476 19754 4544 19810
rect 4600 19754 4668 19810
rect 4724 19754 4734 19810
rect 2798 19686 4734 19754
rect 2798 19630 2808 19686
rect 2864 19630 2932 19686
rect 2988 19630 3056 19686
rect 3112 19630 3180 19686
rect 3236 19630 3304 19686
rect 3360 19630 3428 19686
rect 3484 19630 3552 19686
rect 3608 19630 3676 19686
rect 3732 19630 3800 19686
rect 3856 19630 3924 19686
rect 3980 19630 4048 19686
rect 4104 19630 4172 19686
rect 4228 19630 4296 19686
rect 4352 19630 4420 19686
rect 4476 19630 4544 19686
rect 4600 19630 4668 19686
rect 4724 19630 4734 19686
rect 2798 19562 4734 19630
rect 2798 19506 2808 19562
rect 2864 19506 2932 19562
rect 2988 19506 3056 19562
rect 3112 19506 3180 19562
rect 3236 19506 3304 19562
rect 3360 19506 3428 19562
rect 3484 19506 3552 19562
rect 3608 19506 3676 19562
rect 3732 19506 3800 19562
rect 3856 19506 3924 19562
rect 3980 19506 4048 19562
rect 4104 19506 4172 19562
rect 4228 19506 4296 19562
rect 4352 19506 4420 19562
rect 4476 19506 4544 19562
rect 4600 19506 4668 19562
rect 4724 19506 4734 19562
rect 2798 19438 4734 19506
rect 2798 19382 2808 19438
rect 2864 19382 2932 19438
rect 2988 19382 3056 19438
rect 3112 19382 3180 19438
rect 3236 19382 3304 19438
rect 3360 19382 3428 19438
rect 3484 19382 3552 19438
rect 3608 19382 3676 19438
rect 3732 19382 3800 19438
rect 3856 19382 3924 19438
rect 3980 19382 4048 19438
rect 4104 19382 4172 19438
rect 4228 19382 4296 19438
rect 4352 19382 4420 19438
rect 4476 19382 4544 19438
rect 4600 19382 4668 19438
rect 4724 19382 4734 19438
rect 2798 19314 4734 19382
rect 2798 19258 2808 19314
rect 2864 19258 2932 19314
rect 2988 19258 3056 19314
rect 3112 19258 3180 19314
rect 3236 19258 3304 19314
rect 3360 19258 3428 19314
rect 3484 19258 3552 19314
rect 3608 19258 3676 19314
rect 3732 19258 3800 19314
rect 3856 19258 3924 19314
rect 3980 19258 4048 19314
rect 4104 19258 4172 19314
rect 4228 19258 4296 19314
rect 4352 19258 4420 19314
rect 4476 19258 4544 19314
rect 4600 19258 4668 19314
rect 4724 19258 4734 19314
rect 2798 19190 4734 19258
rect 2798 19134 2808 19190
rect 2864 19134 2932 19190
rect 2988 19134 3056 19190
rect 3112 19134 3180 19190
rect 3236 19134 3304 19190
rect 3360 19134 3428 19190
rect 3484 19134 3552 19190
rect 3608 19134 3676 19190
rect 3732 19134 3800 19190
rect 3856 19134 3924 19190
rect 3980 19134 4048 19190
rect 4104 19134 4172 19190
rect 4228 19134 4296 19190
rect 4352 19134 4420 19190
rect 4476 19134 4544 19190
rect 4600 19134 4668 19190
rect 4724 19134 4734 19190
rect 2798 19066 4734 19134
rect 2798 19010 2808 19066
rect 2864 19010 2932 19066
rect 2988 19010 3056 19066
rect 3112 19010 3180 19066
rect 3236 19010 3304 19066
rect 3360 19010 3428 19066
rect 3484 19010 3552 19066
rect 3608 19010 3676 19066
rect 3732 19010 3800 19066
rect 3856 19010 3924 19066
rect 3980 19010 4048 19066
rect 4104 19010 4172 19066
rect 4228 19010 4296 19066
rect 4352 19010 4420 19066
rect 4476 19010 4544 19066
rect 4600 19010 4668 19066
rect 4724 19010 4734 19066
rect 2798 18942 4734 19010
rect 2798 18886 2808 18942
rect 2864 18886 2932 18942
rect 2988 18886 3056 18942
rect 3112 18886 3180 18942
rect 3236 18886 3304 18942
rect 3360 18886 3428 18942
rect 3484 18886 3552 18942
rect 3608 18886 3676 18942
rect 3732 18886 3800 18942
rect 3856 18886 3924 18942
rect 3980 18886 4048 18942
rect 4104 18886 4172 18942
rect 4228 18886 4296 18942
rect 4352 18886 4420 18942
rect 4476 18886 4544 18942
rect 4600 18886 4668 18942
rect 4724 18886 4734 18942
rect 2798 18818 4734 18886
rect 2798 18762 2808 18818
rect 2864 18762 2932 18818
rect 2988 18762 3056 18818
rect 3112 18762 3180 18818
rect 3236 18762 3304 18818
rect 3360 18762 3428 18818
rect 3484 18762 3552 18818
rect 3608 18762 3676 18818
rect 3732 18762 3800 18818
rect 3856 18762 3924 18818
rect 3980 18762 4048 18818
rect 4104 18762 4172 18818
rect 4228 18762 4296 18818
rect 4352 18762 4420 18818
rect 4476 18762 4544 18818
rect 4600 18762 4668 18818
rect 4724 18762 4734 18818
rect 2798 18694 4734 18762
rect 2798 18638 2808 18694
rect 2864 18638 2932 18694
rect 2988 18638 3056 18694
rect 3112 18638 3180 18694
rect 3236 18638 3304 18694
rect 3360 18638 3428 18694
rect 3484 18638 3552 18694
rect 3608 18638 3676 18694
rect 3732 18638 3800 18694
rect 3856 18638 3924 18694
rect 3980 18638 4048 18694
rect 4104 18638 4172 18694
rect 4228 18638 4296 18694
rect 4352 18638 4420 18694
rect 4476 18638 4544 18694
rect 4600 18638 4668 18694
rect 4724 18638 4734 18694
rect 2798 18570 4734 18638
rect 2798 18514 2808 18570
rect 2864 18514 2932 18570
rect 2988 18514 3056 18570
rect 3112 18514 3180 18570
rect 3236 18514 3304 18570
rect 3360 18514 3428 18570
rect 3484 18514 3552 18570
rect 3608 18514 3676 18570
rect 3732 18514 3800 18570
rect 3856 18514 3924 18570
rect 3980 18514 4048 18570
rect 4104 18514 4172 18570
rect 4228 18514 4296 18570
rect 4352 18514 4420 18570
rect 4476 18514 4544 18570
rect 4600 18514 4668 18570
rect 4724 18514 4734 18570
rect 2798 18446 4734 18514
rect 2798 18390 2808 18446
rect 2864 18390 2932 18446
rect 2988 18390 3056 18446
rect 3112 18390 3180 18446
rect 3236 18390 3304 18446
rect 3360 18390 3428 18446
rect 3484 18390 3552 18446
rect 3608 18390 3676 18446
rect 3732 18390 3800 18446
rect 3856 18390 3924 18446
rect 3980 18390 4048 18446
rect 4104 18390 4172 18446
rect 4228 18390 4296 18446
rect 4352 18390 4420 18446
rect 4476 18390 4544 18446
rect 4600 18390 4668 18446
rect 4724 18390 4734 18446
rect 2798 18322 4734 18390
rect 2798 18266 2808 18322
rect 2864 18266 2932 18322
rect 2988 18266 3056 18322
rect 3112 18266 3180 18322
rect 3236 18266 3304 18322
rect 3360 18266 3428 18322
rect 3484 18266 3552 18322
rect 3608 18266 3676 18322
rect 3732 18266 3800 18322
rect 3856 18266 3924 18322
rect 3980 18266 4048 18322
rect 4104 18266 4172 18322
rect 4228 18266 4296 18322
rect 4352 18266 4420 18322
rect 4476 18266 4544 18322
rect 4600 18266 4668 18322
rect 4724 18266 4734 18322
rect 2798 18198 4734 18266
rect 2798 18142 2808 18198
rect 2864 18142 2932 18198
rect 2988 18142 3056 18198
rect 3112 18142 3180 18198
rect 3236 18142 3304 18198
rect 3360 18142 3428 18198
rect 3484 18142 3552 18198
rect 3608 18142 3676 18198
rect 3732 18142 3800 18198
rect 3856 18142 3924 18198
rect 3980 18142 4048 18198
rect 4104 18142 4172 18198
rect 4228 18142 4296 18198
rect 4352 18142 4420 18198
rect 4476 18142 4544 18198
rect 4600 18142 4668 18198
rect 4724 18142 4734 18198
rect 2798 18074 4734 18142
rect 2798 18018 2808 18074
rect 2864 18018 2932 18074
rect 2988 18018 3056 18074
rect 3112 18018 3180 18074
rect 3236 18018 3304 18074
rect 3360 18018 3428 18074
rect 3484 18018 3552 18074
rect 3608 18018 3676 18074
rect 3732 18018 3800 18074
rect 3856 18018 3924 18074
rect 3980 18018 4048 18074
rect 4104 18018 4172 18074
rect 4228 18018 4296 18074
rect 4352 18018 4420 18074
rect 4476 18018 4544 18074
rect 4600 18018 4668 18074
rect 4724 18018 4734 18074
rect 2798 17950 4734 18018
rect 2798 17894 2808 17950
rect 2864 17894 2932 17950
rect 2988 17894 3056 17950
rect 3112 17894 3180 17950
rect 3236 17894 3304 17950
rect 3360 17894 3428 17950
rect 3484 17894 3552 17950
rect 3608 17894 3676 17950
rect 3732 17894 3800 17950
rect 3856 17894 3924 17950
rect 3980 17894 4048 17950
rect 4104 17894 4172 17950
rect 4228 17894 4296 17950
rect 4352 17894 4420 17950
rect 4476 17894 4544 17950
rect 4600 17894 4668 17950
rect 4724 17894 4734 17950
rect 2798 17826 4734 17894
rect 2798 17770 2808 17826
rect 2864 17770 2932 17826
rect 2988 17770 3056 17826
rect 3112 17770 3180 17826
rect 3236 17770 3304 17826
rect 3360 17770 3428 17826
rect 3484 17770 3552 17826
rect 3608 17770 3676 17826
rect 3732 17770 3800 17826
rect 3856 17770 3924 17826
rect 3980 17770 4048 17826
rect 4104 17770 4172 17826
rect 4228 17770 4296 17826
rect 4352 17770 4420 17826
rect 4476 17770 4544 17826
rect 4600 17770 4668 17826
rect 4724 17770 4734 17826
rect 2798 17702 4734 17770
rect 2798 17646 2808 17702
rect 2864 17646 2932 17702
rect 2988 17646 3056 17702
rect 3112 17646 3180 17702
rect 3236 17646 3304 17702
rect 3360 17646 3428 17702
rect 3484 17646 3552 17702
rect 3608 17646 3676 17702
rect 3732 17646 3800 17702
rect 3856 17646 3924 17702
rect 3980 17646 4048 17702
rect 4104 17646 4172 17702
rect 4228 17646 4296 17702
rect 4352 17646 4420 17702
rect 4476 17646 4544 17702
rect 4600 17646 4668 17702
rect 4724 17646 4734 17702
rect 2798 17636 4734 17646
rect 5168 20554 7104 20564
rect 5168 20498 5178 20554
rect 5234 20498 5302 20554
rect 5358 20498 5426 20554
rect 5482 20498 5550 20554
rect 5606 20498 5674 20554
rect 5730 20498 5798 20554
rect 5854 20498 5922 20554
rect 5978 20498 6046 20554
rect 6102 20498 6170 20554
rect 6226 20498 6294 20554
rect 6350 20498 6418 20554
rect 6474 20498 6542 20554
rect 6598 20498 6666 20554
rect 6722 20498 6790 20554
rect 6846 20498 6914 20554
rect 6970 20498 7038 20554
rect 7094 20498 7104 20554
rect 5168 20430 7104 20498
rect 5168 20374 5178 20430
rect 5234 20374 5302 20430
rect 5358 20374 5426 20430
rect 5482 20374 5550 20430
rect 5606 20374 5674 20430
rect 5730 20374 5798 20430
rect 5854 20374 5922 20430
rect 5978 20374 6046 20430
rect 6102 20374 6170 20430
rect 6226 20374 6294 20430
rect 6350 20374 6418 20430
rect 6474 20374 6542 20430
rect 6598 20374 6666 20430
rect 6722 20374 6790 20430
rect 6846 20374 6914 20430
rect 6970 20374 7038 20430
rect 7094 20374 7104 20430
rect 5168 20306 7104 20374
rect 5168 20250 5178 20306
rect 5234 20250 5302 20306
rect 5358 20250 5426 20306
rect 5482 20250 5550 20306
rect 5606 20250 5674 20306
rect 5730 20250 5798 20306
rect 5854 20250 5922 20306
rect 5978 20250 6046 20306
rect 6102 20250 6170 20306
rect 6226 20250 6294 20306
rect 6350 20250 6418 20306
rect 6474 20250 6542 20306
rect 6598 20250 6666 20306
rect 6722 20250 6790 20306
rect 6846 20250 6914 20306
rect 6970 20250 7038 20306
rect 7094 20250 7104 20306
rect 5168 20182 7104 20250
rect 5168 20126 5178 20182
rect 5234 20126 5302 20182
rect 5358 20126 5426 20182
rect 5482 20126 5550 20182
rect 5606 20126 5674 20182
rect 5730 20126 5798 20182
rect 5854 20126 5922 20182
rect 5978 20126 6046 20182
rect 6102 20126 6170 20182
rect 6226 20126 6294 20182
rect 6350 20126 6418 20182
rect 6474 20126 6542 20182
rect 6598 20126 6666 20182
rect 6722 20126 6790 20182
rect 6846 20126 6914 20182
rect 6970 20126 7038 20182
rect 7094 20126 7104 20182
rect 5168 20058 7104 20126
rect 5168 20002 5178 20058
rect 5234 20002 5302 20058
rect 5358 20002 5426 20058
rect 5482 20002 5550 20058
rect 5606 20002 5674 20058
rect 5730 20002 5798 20058
rect 5854 20002 5922 20058
rect 5978 20002 6046 20058
rect 6102 20002 6170 20058
rect 6226 20002 6294 20058
rect 6350 20002 6418 20058
rect 6474 20002 6542 20058
rect 6598 20002 6666 20058
rect 6722 20002 6790 20058
rect 6846 20002 6914 20058
rect 6970 20002 7038 20058
rect 7094 20002 7104 20058
rect 5168 19934 7104 20002
rect 5168 19878 5178 19934
rect 5234 19878 5302 19934
rect 5358 19878 5426 19934
rect 5482 19878 5550 19934
rect 5606 19878 5674 19934
rect 5730 19878 5798 19934
rect 5854 19878 5922 19934
rect 5978 19878 6046 19934
rect 6102 19878 6170 19934
rect 6226 19878 6294 19934
rect 6350 19878 6418 19934
rect 6474 19878 6542 19934
rect 6598 19878 6666 19934
rect 6722 19878 6790 19934
rect 6846 19878 6914 19934
rect 6970 19878 7038 19934
rect 7094 19878 7104 19934
rect 5168 19810 7104 19878
rect 5168 19754 5178 19810
rect 5234 19754 5302 19810
rect 5358 19754 5426 19810
rect 5482 19754 5550 19810
rect 5606 19754 5674 19810
rect 5730 19754 5798 19810
rect 5854 19754 5922 19810
rect 5978 19754 6046 19810
rect 6102 19754 6170 19810
rect 6226 19754 6294 19810
rect 6350 19754 6418 19810
rect 6474 19754 6542 19810
rect 6598 19754 6666 19810
rect 6722 19754 6790 19810
rect 6846 19754 6914 19810
rect 6970 19754 7038 19810
rect 7094 19754 7104 19810
rect 5168 19686 7104 19754
rect 5168 19630 5178 19686
rect 5234 19630 5302 19686
rect 5358 19630 5426 19686
rect 5482 19630 5550 19686
rect 5606 19630 5674 19686
rect 5730 19630 5798 19686
rect 5854 19630 5922 19686
rect 5978 19630 6046 19686
rect 6102 19630 6170 19686
rect 6226 19630 6294 19686
rect 6350 19630 6418 19686
rect 6474 19630 6542 19686
rect 6598 19630 6666 19686
rect 6722 19630 6790 19686
rect 6846 19630 6914 19686
rect 6970 19630 7038 19686
rect 7094 19630 7104 19686
rect 5168 19562 7104 19630
rect 5168 19506 5178 19562
rect 5234 19506 5302 19562
rect 5358 19506 5426 19562
rect 5482 19506 5550 19562
rect 5606 19506 5674 19562
rect 5730 19506 5798 19562
rect 5854 19506 5922 19562
rect 5978 19506 6046 19562
rect 6102 19506 6170 19562
rect 6226 19506 6294 19562
rect 6350 19506 6418 19562
rect 6474 19506 6542 19562
rect 6598 19506 6666 19562
rect 6722 19506 6790 19562
rect 6846 19506 6914 19562
rect 6970 19506 7038 19562
rect 7094 19506 7104 19562
rect 5168 19438 7104 19506
rect 5168 19382 5178 19438
rect 5234 19382 5302 19438
rect 5358 19382 5426 19438
rect 5482 19382 5550 19438
rect 5606 19382 5674 19438
rect 5730 19382 5798 19438
rect 5854 19382 5922 19438
rect 5978 19382 6046 19438
rect 6102 19382 6170 19438
rect 6226 19382 6294 19438
rect 6350 19382 6418 19438
rect 6474 19382 6542 19438
rect 6598 19382 6666 19438
rect 6722 19382 6790 19438
rect 6846 19382 6914 19438
rect 6970 19382 7038 19438
rect 7094 19382 7104 19438
rect 5168 19314 7104 19382
rect 5168 19258 5178 19314
rect 5234 19258 5302 19314
rect 5358 19258 5426 19314
rect 5482 19258 5550 19314
rect 5606 19258 5674 19314
rect 5730 19258 5798 19314
rect 5854 19258 5922 19314
rect 5978 19258 6046 19314
rect 6102 19258 6170 19314
rect 6226 19258 6294 19314
rect 6350 19258 6418 19314
rect 6474 19258 6542 19314
rect 6598 19258 6666 19314
rect 6722 19258 6790 19314
rect 6846 19258 6914 19314
rect 6970 19258 7038 19314
rect 7094 19258 7104 19314
rect 5168 19190 7104 19258
rect 5168 19134 5178 19190
rect 5234 19134 5302 19190
rect 5358 19134 5426 19190
rect 5482 19134 5550 19190
rect 5606 19134 5674 19190
rect 5730 19134 5798 19190
rect 5854 19134 5922 19190
rect 5978 19134 6046 19190
rect 6102 19134 6170 19190
rect 6226 19134 6294 19190
rect 6350 19134 6418 19190
rect 6474 19134 6542 19190
rect 6598 19134 6666 19190
rect 6722 19134 6790 19190
rect 6846 19134 6914 19190
rect 6970 19134 7038 19190
rect 7094 19134 7104 19190
rect 5168 19066 7104 19134
rect 5168 19010 5178 19066
rect 5234 19010 5302 19066
rect 5358 19010 5426 19066
rect 5482 19010 5550 19066
rect 5606 19010 5674 19066
rect 5730 19010 5798 19066
rect 5854 19010 5922 19066
rect 5978 19010 6046 19066
rect 6102 19010 6170 19066
rect 6226 19010 6294 19066
rect 6350 19010 6418 19066
rect 6474 19010 6542 19066
rect 6598 19010 6666 19066
rect 6722 19010 6790 19066
rect 6846 19010 6914 19066
rect 6970 19010 7038 19066
rect 7094 19010 7104 19066
rect 5168 18942 7104 19010
rect 5168 18886 5178 18942
rect 5234 18886 5302 18942
rect 5358 18886 5426 18942
rect 5482 18886 5550 18942
rect 5606 18886 5674 18942
rect 5730 18886 5798 18942
rect 5854 18886 5922 18942
rect 5978 18886 6046 18942
rect 6102 18886 6170 18942
rect 6226 18886 6294 18942
rect 6350 18886 6418 18942
rect 6474 18886 6542 18942
rect 6598 18886 6666 18942
rect 6722 18886 6790 18942
rect 6846 18886 6914 18942
rect 6970 18886 7038 18942
rect 7094 18886 7104 18942
rect 5168 18818 7104 18886
rect 5168 18762 5178 18818
rect 5234 18762 5302 18818
rect 5358 18762 5426 18818
rect 5482 18762 5550 18818
rect 5606 18762 5674 18818
rect 5730 18762 5798 18818
rect 5854 18762 5922 18818
rect 5978 18762 6046 18818
rect 6102 18762 6170 18818
rect 6226 18762 6294 18818
rect 6350 18762 6418 18818
rect 6474 18762 6542 18818
rect 6598 18762 6666 18818
rect 6722 18762 6790 18818
rect 6846 18762 6914 18818
rect 6970 18762 7038 18818
rect 7094 18762 7104 18818
rect 5168 18694 7104 18762
rect 5168 18638 5178 18694
rect 5234 18638 5302 18694
rect 5358 18638 5426 18694
rect 5482 18638 5550 18694
rect 5606 18638 5674 18694
rect 5730 18638 5798 18694
rect 5854 18638 5922 18694
rect 5978 18638 6046 18694
rect 6102 18638 6170 18694
rect 6226 18638 6294 18694
rect 6350 18638 6418 18694
rect 6474 18638 6542 18694
rect 6598 18638 6666 18694
rect 6722 18638 6790 18694
rect 6846 18638 6914 18694
rect 6970 18638 7038 18694
rect 7094 18638 7104 18694
rect 5168 18570 7104 18638
rect 5168 18514 5178 18570
rect 5234 18514 5302 18570
rect 5358 18514 5426 18570
rect 5482 18514 5550 18570
rect 5606 18514 5674 18570
rect 5730 18514 5798 18570
rect 5854 18514 5922 18570
rect 5978 18514 6046 18570
rect 6102 18514 6170 18570
rect 6226 18514 6294 18570
rect 6350 18514 6418 18570
rect 6474 18514 6542 18570
rect 6598 18514 6666 18570
rect 6722 18514 6790 18570
rect 6846 18514 6914 18570
rect 6970 18514 7038 18570
rect 7094 18514 7104 18570
rect 5168 18446 7104 18514
rect 5168 18390 5178 18446
rect 5234 18390 5302 18446
rect 5358 18390 5426 18446
rect 5482 18390 5550 18446
rect 5606 18390 5674 18446
rect 5730 18390 5798 18446
rect 5854 18390 5922 18446
rect 5978 18390 6046 18446
rect 6102 18390 6170 18446
rect 6226 18390 6294 18446
rect 6350 18390 6418 18446
rect 6474 18390 6542 18446
rect 6598 18390 6666 18446
rect 6722 18390 6790 18446
rect 6846 18390 6914 18446
rect 6970 18390 7038 18446
rect 7094 18390 7104 18446
rect 5168 18322 7104 18390
rect 5168 18266 5178 18322
rect 5234 18266 5302 18322
rect 5358 18266 5426 18322
rect 5482 18266 5550 18322
rect 5606 18266 5674 18322
rect 5730 18266 5798 18322
rect 5854 18266 5922 18322
rect 5978 18266 6046 18322
rect 6102 18266 6170 18322
rect 6226 18266 6294 18322
rect 6350 18266 6418 18322
rect 6474 18266 6542 18322
rect 6598 18266 6666 18322
rect 6722 18266 6790 18322
rect 6846 18266 6914 18322
rect 6970 18266 7038 18322
rect 7094 18266 7104 18322
rect 5168 18198 7104 18266
rect 5168 18142 5178 18198
rect 5234 18142 5302 18198
rect 5358 18142 5426 18198
rect 5482 18142 5550 18198
rect 5606 18142 5674 18198
rect 5730 18142 5798 18198
rect 5854 18142 5922 18198
rect 5978 18142 6046 18198
rect 6102 18142 6170 18198
rect 6226 18142 6294 18198
rect 6350 18142 6418 18198
rect 6474 18142 6542 18198
rect 6598 18142 6666 18198
rect 6722 18142 6790 18198
rect 6846 18142 6914 18198
rect 6970 18142 7038 18198
rect 7094 18142 7104 18198
rect 5168 18074 7104 18142
rect 5168 18018 5178 18074
rect 5234 18018 5302 18074
rect 5358 18018 5426 18074
rect 5482 18018 5550 18074
rect 5606 18018 5674 18074
rect 5730 18018 5798 18074
rect 5854 18018 5922 18074
rect 5978 18018 6046 18074
rect 6102 18018 6170 18074
rect 6226 18018 6294 18074
rect 6350 18018 6418 18074
rect 6474 18018 6542 18074
rect 6598 18018 6666 18074
rect 6722 18018 6790 18074
rect 6846 18018 6914 18074
rect 6970 18018 7038 18074
rect 7094 18018 7104 18074
rect 5168 17950 7104 18018
rect 5168 17894 5178 17950
rect 5234 17894 5302 17950
rect 5358 17894 5426 17950
rect 5482 17894 5550 17950
rect 5606 17894 5674 17950
rect 5730 17894 5798 17950
rect 5854 17894 5922 17950
rect 5978 17894 6046 17950
rect 6102 17894 6170 17950
rect 6226 17894 6294 17950
rect 6350 17894 6418 17950
rect 6474 17894 6542 17950
rect 6598 17894 6666 17950
rect 6722 17894 6790 17950
rect 6846 17894 6914 17950
rect 6970 17894 7038 17950
rect 7094 17894 7104 17950
rect 5168 17826 7104 17894
rect 5168 17770 5178 17826
rect 5234 17770 5302 17826
rect 5358 17770 5426 17826
rect 5482 17770 5550 17826
rect 5606 17770 5674 17826
rect 5730 17770 5798 17826
rect 5854 17770 5922 17826
rect 5978 17770 6046 17826
rect 6102 17770 6170 17826
rect 6226 17770 6294 17826
rect 6350 17770 6418 17826
rect 6474 17770 6542 17826
rect 6598 17770 6666 17826
rect 6722 17770 6790 17826
rect 6846 17770 6914 17826
rect 6970 17770 7038 17826
rect 7094 17770 7104 17826
rect 5168 17702 7104 17770
rect 5168 17646 5178 17702
rect 5234 17646 5302 17702
rect 5358 17646 5426 17702
rect 5482 17646 5550 17702
rect 5606 17646 5674 17702
rect 5730 17646 5798 17702
rect 5854 17646 5922 17702
rect 5978 17646 6046 17702
rect 6102 17646 6170 17702
rect 6226 17646 6294 17702
rect 6350 17646 6418 17702
rect 6474 17646 6542 17702
rect 6598 17646 6666 17702
rect 6722 17646 6790 17702
rect 6846 17646 6914 17702
rect 6970 17646 7038 17702
rect 7094 17646 7104 17702
rect 5168 17636 7104 17646
rect 7874 20554 9810 20564
rect 7874 20498 7884 20554
rect 7940 20498 8008 20554
rect 8064 20498 8132 20554
rect 8188 20498 8256 20554
rect 8312 20498 8380 20554
rect 8436 20498 8504 20554
rect 8560 20498 8628 20554
rect 8684 20498 8752 20554
rect 8808 20498 8876 20554
rect 8932 20498 9000 20554
rect 9056 20498 9124 20554
rect 9180 20498 9248 20554
rect 9304 20498 9372 20554
rect 9428 20498 9496 20554
rect 9552 20498 9620 20554
rect 9676 20498 9744 20554
rect 9800 20498 9810 20554
rect 7874 20430 9810 20498
rect 7874 20374 7884 20430
rect 7940 20374 8008 20430
rect 8064 20374 8132 20430
rect 8188 20374 8256 20430
rect 8312 20374 8380 20430
rect 8436 20374 8504 20430
rect 8560 20374 8628 20430
rect 8684 20374 8752 20430
rect 8808 20374 8876 20430
rect 8932 20374 9000 20430
rect 9056 20374 9124 20430
rect 9180 20374 9248 20430
rect 9304 20374 9372 20430
rect 9428 20374 9496 20430
rect 9552 20374 9620 20430
rect 9676 20374 9744 20430
rect 9800 20374 9810 20430
rect 7874 20306 9810 20374
rect 7874 20250 7884 20306
rect 7940 20250 8008 20306
rect 8064 20250 8132 20306
rect 8188 20250 8256 20306
rect 8312 20250 8380 20306
rect 8436 20250 8504 20306
rect 8560 20250 8628 20306
rect 8684 20250 8752 20306
rect 8808 20250 8876 20306
rect 8932 20250 9000 20306
rect 9056 20250 9124 20306
rect 9180 20250 9248 20306
rect 9304 20250 9372 20306
rect 9428 20250 9496 20306
rect 9552 20250 9620 20306
rect 9676 20250 9744 20306
rect 9800 20250 9810 20306
rect 7874 20182 9810 20250
rect 7874 20126 7884 20182
rect 7940 20126 8008 20182
rect 8064 20126 8132 20182
rect 8188 20126 8256 20182
rect 8312 20126 8380 20182
rect 8436 20126 8504 20182
rect 8560 20126 8628 20182
rect 8684 20126 8752 20182
rect 8808 20126 8876 20182
rect 8932 20126 9000 20182
rect 9056 20126 9124 20182
rect 9180 20126 9248 20182
rect 9304 20126 9372 20182
rect 9428 20126 9496 20182
rect 9552 20126 9620 20182
rect 9676 20126 9744 20182
rect 9800 20126 9810 20182
rect 7874 20058 9810 20126
rect 7874 20002 7884 20058
rect 7940 20002 8008 20058
rect 8064 20002 8132 20058
rect 8188 20002 8256 20058
rect 8312 20002 8380 20058
rect 8436 20002 8504 20058
rect 8560 20002 8628 20058
rect 8684 20002 8752 20058
rect 8808 20002 8876 20058
rect 8932 20002 9000 20058
rect 9056 20002 9124 20058
rect 9180 20002 9248 20058
rect 9304 20002 9372 20058
rect 9428 20002 9496 20058
rect 9552 20002 9620 20058
rect 9676 20002 9744 20058
rect 9800 20002 9810 20058
rect 7874 19934 9810 20002
rect 7874 19878 7884 19934
rect 7940 19878 8008 19934
rect 8064 19878 8132 19934
rect 8188 19878 8256 19934
rect 8312 19878 8380 19934
rect 8436 19878 8504 19934
rect 8560 19878 8628 19934
rect 8684 19878 8752 19934
rect 8808 19878 8876 19934
rect 8932 19878 9000 19934
rect 9056 19878 9124 19934
rect 9180 19878 9248 19934
rect 9304 19878 9372 19934
rect 9428 19878 9496 19934
rect 9552 19878 9620 19934
rect 9676 19878 9744 19934
rect 9800 19878 9810 19934
rect 7874 19810 9810 19878
rect 7874 19754 7884 19810
rect 7940 19754 8008 19810
rect 8064 19754 8132 19810
rect 8188 19754 8256 19810
rect 8312 19754 8380 19810
rect 8436 19754 8504 19810
rect 8560 19754 8628 19810
rect 8684 19754 8752 19810
rect 8808 19754 8876 19810
rect 8932 19754 9000 19810
rect 9056 19754 9124 19810
rect 9180 19754 9248 19810
rect 9304 19754 9372 19810
rect 9428 19754 9496 19810
rect 9552 19754 9620 19810
rect 9676 19754 9744 19810
rect 9800 19754 9810 19810
rect 7874 19686 9810 19754
rect 7874 19630 7884 19686
rect 7940 19630 8008 19686
rect 8064 19630 8132 19686
rect 8188 19630 8256 19686
rect 8312 19630 8380 19686
rect 8436 19630 8504 19686
rect 8560 19630 8628 19686
rect 8684 19630 8752 19686
rect 8808 19630 8876 19686
rect 8932 19630 9000 19686
rect 9056 19630 9124 19686
rect 9180 19630 9248 19686
rect 9304 19630 9372 19686
rect 9428 19630 9496 19686
rect 9552 19630 9620 19686
rect 9676 19630 9744 19686
rect 9800 19630 9810 19686
rect 7874 19562 9810 19630
rect 7874 19506 7884 19562
rect 7940 19506 8008 19562
rect 8064 19506 8132 19562
rect 8188 19506 8256 19562
rect 8312 19506 8380 19562
rect 8436 19506 8504 19562
rect 8560 19506 8628 19562
rect 8684 19506 8752 19562
rect 8808 19506 8876 19562
rect 8932 19506 9000 19562
rect 9056 19506 9124 19562
rect 9180 19506 9248 19562
rect 9304 19506 9372 19562
rect 9428 19506 9496 19562
rect 9552 19506 9620 19562
rect 9676 19506 9744 19562
rect 9800 19506 9810 19562
rect 7874 19438 9810 19506
rect 7874 19382 7884 19438
rect 7940 19382 8008 19438
rect 8064 19382 8132 19438
rect 8188 19382 8256 19438
rect 8312 19382 8380 19438
rect 8436 19382 8504 19438
rect 8560 19382 8628 19438
rect 8684 19382 8752 19438
rect 8808 19382 8876 19438
rect 8932 19382 9000 19438
rect 9056 19382 9124 19438
rect 9180 19382 9248 19438
rect 9304 19382 9372 19438
rect 9428 19382 9496 19438
rect 9552 19382 9620 19438
rect 9676 19382 9744 19438
rect 9800 19382 9810 19438
rect 7874 19314 9810 19382
rect 7874 19258 7884 19314
rect 7940 19258 8008 19314
rect 8064 19258 8132 19314
rect 8188 19258 8256 19314
rect 8312 19258 8380 19314
rect 8436 19258 8504 19314
rect 8560 19258 8628 19314
rect 8684 19258 8752 19314
rect 8808 19258 8876 19314
rect 8932 19258 9000 19314
rect 9056 19258 9124 19314
rect 9180 19258 9248 19314
rect 9304 19258 9372 19314
rect 9428 19258 9496 19314
rect 9552 19258 9620 19314
rect 9676 19258 9744 19314
rect 9800 19258 9810 19314
rect 7874 19190 9810 19258
rect 7874 19134 7884 19190
rect 7940 19134 8008 19190
rect 8064 19134 8132 19190
rect 8188 19134 8256 19190
rect 8312 19134 8380 19190
rect 8436 19134 8504 19190
rect 8560 19134 8628 19190
rect 8684 19134 8752 19190
rect 8808 19134 8876 19190
rect 8932 19134 9000 19190
rect 9056 19134 9124 19190
rect 9180 19134 9248 19190
rect 9304 19134 9372 19190
rect 9428 19134 9496 19190
rect 9552 19134 9620 19190
rect 9676 19134 9744 19190
rect 9800 19134 9810 19190
rect 7874 19066 9810 19134
rect 7874 19010 7884 19066
rect 7940 19010 8008 19066
rect 8064 19010 8132 19066
rect 8188 19010 8256 19066
rect 8312 19010 8380 19066
rect 8436 19010 8504 19066
rect 8560 19010 8628 19066
rect 8684 19010 8752 19066
rect 8808 19010 8876 19066
rect 8932 19010 9000 19066
rect 9056 19010 9124 19066
rect 9180 19010 9248 19066
rect 9304 19010 9372 19066
rect 9428 19010 9496 19066
rect 9552 19010 9620 19066
rect 9676 19010 9744 19066
rect 9800 19010 9810 19066
rect 7874 18942 9810 19010
rect 7874 18886 7884 18942
rect 7940 18886 8008 18942
rect 8064 18886 8132 18942
rect 8188 18886 8256 18942
rect 8312 18886 8380 18942
rect 8436 18886 8504 18942
rect 8560 18886 8628 18942
rect 8684 18886 8752 18942
rect 8808 18886 8876 18942
rect 8932 18886 9000 18942
rect 9056 18886 9124 18942
rect 9180 18886 9248 18942
rect 9304 18886 9372 18942
rect 9428 18886 9496 18942
rect 9552 18886 9620 18942
rect 9676 18886 9744 18942
rect 9800 18886 9810 18942
rect 7874 18818 9810 18886
rect 7874 18762 7884 18818
rect 7940 18762 8008 18818
rect 8064 18762 8132 18818
rect 8188 18762 8256 18818
rect 8312 18762 8380 18818
rect 8436 18762 8504 18818
rect 8560 18762 8628 18818
rect 8684 18762 8752 18818
rect 8808 18762 8876 18818
rect 8932 18762 9000 18818
rect 9056 18762 9124 18818
rect 9180 18762 9248 18818
rect 9304 18762 9372 18818
rect 9428 18762 9496 18818
rect 9552 18762 9620 18818
rect 9676 18762 9744 18818
rect 9800 18762 9810 18818
rect 7874 18694 9810 18762
rect 7874 18638 7884 18694
rect 7940 18638 8008 18694
rect 8064 18638 8132 18694
rect 8188 18638 8256 18694
rect 8312 18638 8380 18694
rect 8436 18638 8504 18694
rect 8560 18638 8628 18694
rect 8684 18638 8752 18694
rect 8808 18638 8876 18694
rect 8932 18638 9000 18694
rect 9056 18638 9124 18694
rect 9180 18638 9248 18694
rect 9304 18638 9372 18694
rect 9428 18638 9496 18694
rect 9552 18638 9620 18694
rect 9676 18638 9744 18694
rect 9800 18638 9810 18694
rect 7874 18570 9810 18638
rect 7874 18514 7884 18570
rect 7940 18514 8008 18570
rect 8064 18514 8132 18570
rect 8188 18514 8256 18570
rect 8312 18514 8380 18570
rect 8436 18514 8504 18570
rect 8560 18514 8628 18570
rect 8684 18514 8752 18570
rect 8808 18514 8876 18570
rect 8932 18514 9000 18570
rect 9056 18514 9124 18570
rect 9180 18514 9248 18570
rect 9304 18514 9372 18570
rect 9428 18514 9496 18570
rect 9552 18514 9620 18570
rect 9676 18514 9744 18570
rect 9800 18514 9810 18570
rect 7874 18446 9810 18514
rect 7874 18390 7884 18446
rect 7940 18390 8008 18446
rect 8064 18390 8132 18446
rect 8188 18390 8256 18446
rect 8312 18390 8380 18446
rect 8436 18390 8504 18446
rect 8560 18390 8628 18446
rect 8684 18390 8752 18446
rect 8808 18390 8876 18446
rect 8932 18390 9000 18446
rect 9056 18390 9124 18446
rect 9180 18390 9248 18446
rect 9304 18390 9372 18446
rect 9428 18390 9496 18446
rect 9552 18390 9620 18446
rect 9676 18390 9744 18446
rect 9800 18390 9810 18446
rect 7874 18322 9810 18390
rect 7874 18266 7884 18322
rect 7940 18266 8008 18322
rect 8064 18266 8132 18322
rect 8188 18266 8256 18322
rect 8312 18266 8380 18322
rect 8436 18266 8504 18322
rect 8560 18266 8628 18322
rect 8684 18266 8752 18322
rect 8808 18266 8876 18322
rect 8932 18266 9000 18322
rect 9056 18266 9124 18322
rect 9180 18266 9248 18322
rect 9304 18266 9372 18322
rect 9428 18266 9496 18322
rect 9552 18266 9620 18322
rect 9676 18266 9744 18322
rect 9800 18266 9810 18322
rect 7874 18198 9810 18266
rect 7874 18142 7884 18198
rect 7940 18142 8008 18198
rect 8064 18142 8132 18198
rect 8188 18142 8256 18198
rect 8312 18142 8380 18198
rect 8436 18142 8504 18198
rect 8560 18142 8628 18198
rect 8684 18142 8752 18198
rect 8808 18142 8876 18198
rect 8932 18142 9000 18198
rect 9056 18142 9124 18198
rect 9180 18142 9248 18198
rect 9304 18142 9372 18198
rect 9428 18142 9496 18198
rect 9552 18142 9620 18198
rect 9676 18142 9744 18198
rect 9800 18142 9810 18198
rect 7874 18074 9810 18142
rect 7874 18018 7884 18074
rect 7940 18018 8008 18074
rect 8064 18018 8132 18074
rect 8188 18018 8256 18074
rect 8312 18018 8380 18074
rect 8436 18018 8504 18074
rect 8560 18018 8628 18074
rect 8684 18018 8752 18074
rect 8808 18018 8876 18074
rect 8932 18018 9000 18074
rect 9056 18018 9124 18074
rect 9180 18018 9248 18074
rect 9304 18018 9372 18074
rect 9428 18018 9496 18074
rect 9552 18018 9620 18074
rect 9676 18018 9744 18074
rect 9800 18018 9810 18074
rect 7874 17950 9810 18018
rect 7874 17894 7884 17950
rect 7940 17894 8008 17950
rect 8064 17894 8132 17950
rect 8188 17894 8256 17950
rect 8312 17894 8380 17950
rect 8436 17894 8504 17950
rect 8560 17894 8628 17950
rect 8684 17894 8752 17950
rect 8808 17894 8876 17950
rect 8932 17894 9000 17950
rect 9056 17894 9124 17950
rect 9180 17894 9248 17950
rect 9304 17894 9372 17950
rect 9428 17894 9496 17950
rect 9552 17894 9620 17950
rect 9676 17894 9744 17950
rect 9800 17894 9810 17950
rect 7874 17826 9810 17894
rect 7874 17770 7884 17826
rect 7940 17770 8008 17826
rect 8064 17770 8132 17826
rect 8188 17770 8256 17826
rect 8312 17770 8380 17826
rect 8436 17770 8504 17826
rect 8560 17770 8628 17826
rect 8684 17770 8752 17826
rect 8808 17770 8876 17826
rect 8932 17770 9000 17826
rect 9056 17770 9124 17826
rect 9180 17770 9248 17826
rect 9304 17770 9372 17826
rect 9428 17770 9496 17826
rect 9552 17770 9620 17826
rect 9676 17770 9744 17826
rect 9800 17770 9810 17826
rect 7874 17702 9810 17770
rect 7874 17646 7884 17702
rect 7940 17646 8008 17702
rect 8064 17646 8132 17702
rect 8188 17646 8256 17702
rect 8312 17646 8380 17702
rect 8436 17646 8504 17702
rect 8560 17646 8628 17702
rect 8684 17646 8752 17702
rect 8808 17646 8876 17702
rect 8932 17646 9000 17702
rect 9056 17646 9124 17702
rect 9180 17646 9248 17702
rect 9304 17646 9372 17702
rect 9428 17646 9496 17702
rect 9552 17646 9620 17702
rect 9676 17646 9744 17702
rect 9800 17646 9810 17702
rect 7874 17636 9810 17646
rect 10244 20554 12180 20564
rect 10244 20498 10254 20554
rect 10310 20498 10378 20554
rect 10434 20498 10502 20554
rect 10558 20498 10626 20554
rect 10682 20498 10750 20554
rect 10806 20498 10874 20554
rect 10930 20498 10998 20554
rect 11054 20498 11122 20554
rect 11178 20498 11246 20554
rect 11302 20498 11370 20554
rect 11426 20498 11494 20554
rect 11550 20498 11618 20554
rect 11674 20498 11742 20554
rect 11798 20498 11866 20554
rect 11922 20498 11990 20554
rect 12046 20498 12114 20554
rect 12170 20498 12180 20554
rect 10244 20430 12180 20498
rect 10244 20374 10254 20430
rect 10310 20374 10378 20430
rect 10434 20374 10502 20430
rect 10558 20374 10626 20430
rect 10682 20374 10750 20430
rect 10806 20374 10874 20430
rect 10930 20374 10998 20430
rect 11054 20374 11122 20430
rect 11178 20374 11246 20430
rect 11302 20374 11370 20430
rect 11426 20374 11494 20430
rect 11550 20374 11618 20430
rect 11674 20374 11742 20430
rect 11798 20374 11866 20430
rect 11922 20374 11990 20430
rect 12046 20374 12114 20430
rect 12170 20374 12180 20430
rect 10244 20306 12180 20374
rect 10244 20250 10254 20306
rect 10310 20250 10378 20306
rect 10434 20250 10502 20306
rect 10558 20250 10626 20306
rect 10682 20250 10750 20306
rect 10806 20250 10874 20306
rect 10930 20250 10998 20306
rect 11054 20250 11122 20306
rect 11178 20250 11246 20306
rect 11302 20250 11370 20306
rect 11426 20250 11494 20306
rect 11550 20250 11618 20306
rect 11674 20250 11742 20306
rect 11798 20250 11866 20306
rect 11922 20250 11990 20306
rect 12046 20250 12114 20306
rect 12170 20250 12180 20306
rect 10244 20182 12180 20250
rect 10244 20126 10254 20182
rect 10310 20126 10378 20182
rect 10434 20126 10502 20182
rect 10558 20126 10626 20182
rect 10682 20126 10750 20182
rect 10806 20126 10874 20182
rect 10930 20126 10998 20182
rect 11054 20126 11122 20182
rect 11178 20126 11246 20182
rect 11302 20126 11370 20182
rect 11426 20126 11494 20182
rect 11550 20126 11618 20182
rect 11674 20126 11742 20182
rect 11798 20126 11866 20182
rect 11922 20126 11990 20182
rect 12046 20126 12114 20182
rect 12170 20126 12180 20182
rect 10244 20058 12180 20126
rect 10244 20002 10254 20058
rect 10310 20002 10378 20058
rect 10434 20002 10502 20058
rect 10558 20002 10626 20058
rect 10682 20002 10750 20058
rect 10806 20002 10874 20058
rect 10930 20002 10998 20058
rect 11054 20002 11122 20058
rect 11178 20002 11246 20058
rect 11302 20002 11370 20058
rect 11426 20002 11494 20058
rect 11550 20002 11618 20058
rect 11674 20002 11742 20058
rect 11798 20002 11866 20058
rect 11922 20002 11990 20058
rect 12046 20002 12114 20058
rect 12170 20002 12180 20058
rect 10244 19934 12180 20002
rect 10244 19878 10254 19934
rect 10310 19878 10378 19934
rect 10434 19878 10502 19934
rect 10558 19878 10626 19934
rect 10682 19878 10750 19934
rect 10806 19878 10874 19934
rect 10930 19878 10998 19934
rect 11054 19878 11122 19934
rect 11178 19878 11246 19934
rect 11302 19878 11370 19934
rect 11426 19878 11494 19934
rect 11550 19878 11618 19934
rect 11674 19878 11742 19934
rect 11798 19878 11866 19934
rect 11922 19878 11990 19934
rect 12046 19878 12114 19934
rect 12170 19878 12180 19934
rect 10244 19810 12180 19878
rect 10244 19754 10254 19810
rect 10310 19754 10378 19810
rect 10434 19754 10502 19810
rect 10558 19754 10626 19810
rect 10682 19754 10750 19810
rect 10806 19754 10874 19810
rect 10930 19754 10998 19810
rect 11054 19754 11122 19810
rect 11178 19754 11246 19810
rect 11302 19754 11370 19810
rect 11426 19754 11494 19810
rect 11550 19754 11618 19810
rect 11674 19754 11742 19810
rect 11798 19754 11866 19810
rect 11922 19754 11990 19810
rect 12046 19754 12114 19810
rect 12170 19754 12180 19810
rect 10244 19686 12180 19754
rect 10244 19630 10254 19686
rect 10310 19630 10378 19686
rect 10434 19630 10502 19686
rect 10558 19630 10626 19686
rect 10682 19630 10750 19686
rect 10806 19630 10874 19686
rect 10930 19630 10998 19686
rect 11054 19630 11122 19686
rect 11178 19630 11246 19686
rect 11302 19630 11370 19686
rect 11426 19630 11494 19686
rect 11550 19630 11618 19686
rect 11674 19630 11742 19686
rect 11798 19630 11866 19686
rect 11922 19630 11990 19686
rect 12046 19630 12114 19686
rect 12170 19630 12180 19686
rect 10244 19562 12180 19630
rect 10244 19506 10254 19562
rect 10310 19506 10378 19562
rect 10434 19506 10502 19562
rect 10558 19506 10626 19562
rect 10682 19506 10750 19562
rect 10806 19506 10874 19562
rect 10930 19506 10998 19562
rect 11054 19506 11122 19562
rect 11178 19506 11246 19562
rect 11302 19506 11370 19562
rect 11426 19506 11494 19562
rect 11550 19506 11618 19562
rect 11674 19506 11742 19562
rect 11798 19506 11866 19562
rect 11922 19506 11990 19562
rect 12046 19506 12114 19562
rect 12170 19506 12180 19562
rect 10244 19438 12180 19506
rect 10244 19382 10254 19438
rect 10310 19382 10378 19438
rect 10434 19382 10502 19438
rect 10558 19382 10626 19438
rect 10682 19382 10750 19438
rect 10806 19382 10874 19438
rect 10930 19382 10998 19438
rect 11054 19382 11122 19438
rect 11178 19382 11246 19438
rect 11302 19382 11370 19438
rect 11426 19382 11494 19438
rect 11550 19382 11618 19438
rect 11674 19382 11742 19438
rect 11798 19382 11866 19438
rect 11922 19382 11990 19438
rect 12046 19382 12114 19438
rect 12170 19382 12180 19438
rect 10244 19314 12180 19382
rect 10244 19258 10254 19314
rect 10310 19258 10378 19314
rect 10434 19258 10502 19314
rect 10558 19258 10626 19314
rect 10682 19258 10750 19314
rect 10806 19258 10874 19314
rect 10930 19258 10998 19314
rect 11054 19258 11122 19314
rect 11178 19258 11246 19314
rect 11302 19258 11370 19314
rect 11426 19258 11494 19314
rect 11550 19258 11618 19314
rect 11674 19258 11742 19314
rect 11798 19258 11866 19314
rect 11922 19258 11990 19314
rect 12046 19258 12114 19314
rect 12170 19258 12180 19314
rect 10244 19190 12180 19258
rect 10244 19134 10254 19190
rect 10310 19134 10378 19190
rect 10434 19134 10502 19190
rect 10558 19134 10626 19190
rect 10682 19134 10750 19190
rect 10806 19134 10874 19190
rect 10930 19134 10998 19190
rect 11054 19134 11122 19190
rect 11178 19134 11246 19190
rect 11302 19134 11370 19190
rect 11426 19134 11494 19190
rect 11550 19134 11618 19190
rect 11674 19134 11742 19190
rect 11798 19134 11866 19190
rect 11922 19134 11990 19190
rect 12046 19134 12114 19190
rect 12170 19134 12180 19190
rect 10244 19066 12180 19134
rect 10244 19010 10254 19066
rect 10310 19010 10378 19066
rect 10434 19010 10502 19066
rect 10558 19010 10626 19066
rect 10682 19010 10750 19066
rect 10806 19010 10874 19066
rect 10930 19010 10998 19066
rect 11054 19010 11122 19066
rect 11178 19010 11246 19066
rect 11302 19010 11370 19066
rect 11426 19010 11494 19066
rect 11550 19010 11618 19066
rect 11674 19010 11742 19066
rect 11798 19010 11866 19066
rect 11922 19010 11990 19066
rect 12046 19010 12114 19066
rect 12170 19010 12180 19066
rect 10244 18942 12180 19010
rect 10244 18886 10254 18942
rect 10310 18886 10378 18942
rect 10434 18886 10502 18942
rect 10558 18886 10626 18942
rect 10682 18886 10750 18942
rect 10806 18886 10874 18942
rect 10930 18886 10998 18942
rect 11054 18886 11122 18942
rect 11178 18886 11246 18942
rect 11302 18886 11370 18942
rect 11426 18886 11494 18942
rect 11550 18886 11618 18942
rect 11674 18886 11742 18942
rect 11798 18886 11866 18942
rect 11922 18886 11990 18942
rect 12046 18886 12114 18942
rect 12170 18886 12180 18942
rect 10244 18818 12180 18886
rect 10244 18762 10254 18818
rect 10310 18762 10378 18818
rect 10434 18762 10502 18818
rect 10558 18762 10626 18818
rect 10682 18762 10750 18818
rect 10806 18762 10874 18818
rect 10930 18762 10998 18818
rect 11054 18762 11122 18818
rect 11178 18762 11246 18818
rect 11302 18762 11370 18818
rect 11426 18762 11494 18818
rect 11550 18762 11618 18818
rect 11674 18762 11742 18818
rect 11798 18762 11866 18818
rect 11922 18762 11990 18818
rect 12046 18762 12114 18818
rect 12170 18762 12180 18818
rect 10244 18694 12180 18762
rect 10244 18638 10254 18694
rect 10310 18638 10378 18694
rect 10434 18638 10502 18694
rect 10558 18638 10626 18694
rect 10682 18638 10750 18694
rect 10806 18638 10874 18694
rect 10930 18638 10998 18694
rect 11054 18638 11122 18694
rect 11178 18638 11246 18694
rect 11302 18638 11370 18694
rect 11426 18638 11494 18694
rect 11550 18638 11618 18694
rect 11674 18638 11742 18694
rect 11798 18638 11866 18694
rect 11922 18638 11990 18694
rect 12046 18638 12114 18694
rect 12170 18638 12180 18694
rect 10244 18570 12180 18638
rect 10244 18514 10254 18570
rect 10310 18514 10378 18570
rect 10434 18514 10502 18570
rect 10558 18514 10626 18570
rect 10682 18514 10750 18570
rect 10806 18514 10874 18570
rect 10930 18514 10998 18570
rect 11054 18514 11122 18570
rect 11178 18514 11246 18570
rect 11302 18514 11370 18570
rect 11426 18514 11494 18570
rect 11550 18514 11618 18570
rect 11674 18514 11742 18570
rect 11798 18514 11866 18570
rect 11922 18514 11990 18570
rect 12046 18514 12114 18570
rect 12170 18514 12180 18570
rect 10244 18446 12180 18514
rect 10244 18390 10254 18446
rect 10310 18390 10378 18446
rect 10434 18390 10502 18446
rect 10558 18390 10626 18446
rect 10682 18390 10750 18446
rect 10806 18390 10874 18446
rect 10930 18390 10998 18446
rect 11054 18390 11122 18446
rect 11178 18390 11246 18446
rect 11302 18390 11370 18446
rect 11426 18390 11494 18446
rect 11550 18390 11618 18446
rect 11674 18390 11742 18446
rect 11798 18390 11866 18446
rect 11922 18390 11990 18446
rect 12046 18390 12114 18446
rect 12170 18390 12180 18446
rect 10244 18322 12180 18390
rect 10244 18266 10254 18322
rect 10310 18266 10378 18322
rect 10434 18266 10502 18322
rect 10558 18266 10626 18322
rect 10682 18266 10750 18322
rect 10806 18266 10874 18322
rect 10930 18266 10998 18322
rect 11054 18266 11122 18322
rect 11178 18266 11246 18322
rect 11302 18266 11370 18322
rect 11426 18266 11494 18322
rect 11550 18266 11618 18322
rect 11674 18266 11742 18322
rect 11798 18266 11866 18322
rect 11922 18266 11990 18322
rect 12046 18266 12114 18322
rect 12170 18266 12180 18322
rect 10244 18198 12180 18266
rect 10244 18142 10254 18198
rect 10310 18142 10378 18198
rect 10434 18142 10502 18198
rect 10558 18142 10626 18198
rect 10682 18142 10750 18198
rect 10806 18142 10874 18198
rect 10930 18142 10998 18198
rect 11054 18142 11122 18198
rect 11178 18142 11246 18198
rect 11302 18142 11370 18198
rect 11426 18142 11494 18198
rect 11550 18142 11618 18198
rect 11674 18142 11742 18198
rect 11798 18142 11866 18198
rect 11922 18142 11990 18198
rect 12046 18142 12114 18198
rect 12170 18142 12180 18198
rect 10244 18074 12180 18142
rect 10244 18018 10254 18074
rect 10310 18018 10378 18074
rect 10434 18018 10502 18074
rect 10558 18018 10626 18074
rect 10682 18018 10750 18074
rect 10806 18018 10874 18074
rect 10930 18018 10998 18074
rect 11054 18018 11122 18074
rect 11178 18018 11246 18074
rect 11302 18018 11370 18074
rect 11426 18018 11494 18074
rect 11550 18018 11618 18074
rect 11674 18018 11742 18074
rect 11798 18018 11866 18074
rect 11922 18018 11990 18074
rect 12046 18018 12114 18074
rect 12170 18018 12180 18074
rect 10244 17950 12180 18018
rect 10244 17894 10254 17950
rect 10310 17894 10378 17950
rect 10434 17894 10502 17950
rect 10558 17894 10626 17950
rect 10682 17894 10750 17950
rect 10806 17894 10874 17950
rect 10930 17894 10998 17950
rect 11054 17894 11122 17950
rect 11178 17894 11246 17950
rect 11302 17894 11370 17950
rect 11426 17894 11494 17950
rect 11550 17894 11618 17950
rect 11674 17894 11742 17950
rect 11798 17894 11866 17950
rect 11922 17894 11990 17950
rect 12046 17894 12114 17950
rect 12170 17894 12180 17950
rect 10244 17826 12180 17894
rect 10244 17770 10254 17826
rect 10310 17770 10378 17826
rect 10434 17770 10502 17826
rect 10558 17770 10626 17826
rect 10682 17770 10750 17826
rect 10806 17770 10874 17826
rect 10930 17770 10998 17826
rect 11054 17770 11122 17826
rect 11178 17770 11246 17826
rect 11302 17770 11370 17826
rect 11426 17770 11494 17826
rect 11550 17770 11618 17826
rect 11674 17770 11742 17826
rect 11798 17770 11866 17826
rect 11922 17770 11990 17826
rect 12046 17770 12114 17826
rect 12170 17770 12180 17826
rect 10244 17702 12180 17770
rect 10244 17646 10254 17702
rect 10310 17646 10378 17702
rect 10434 17646 10502 17702
rect 10558 17646 10626 17702
rect 10682 17646 10750 17702
rect 10806 17646 10874 17702
rect 10930 17646 10998 17702
rect 11054 17646 11122 17702
rect 11178 17646 11246 17702
rect 11302 17646 11370 17702
rect 11426 17646 11494 17702
rect 11550 17646 11618 17702
rect 11674 17646 11742 17702
rect 11798 17646 11866 17702
rect 11922 17646 11990 17702
rect 12046 17646 12114 17702
rect 12170 17646 12180 17702
rect 10244 17636 12180 17646
rect 12861 20554 14673 20564
rect 12861 20498 12871 20554
rect 12927 20498 12995 20554
rect 13051 20498 13119 20554
rect 13175 20498 13243 20554
rect 13299 20498 13367 20554
rect 13423 20498 13491 20554
rect 13547 20498 13615 20554
rect 13671 20498 13739 20554
rect 13795 20498 13863 20554
rect 13919 20498 13987 20554
rect 14043 20498 14111 20554
rect 14167 20498 14235 20554
rect 14291 20498 14359 20554
rect 14415 20498 14483 20554
rect 14539 20498 14607 20554
rect 14663 20498 14673 20554
rect 12861 20430 14673 20498
rect 12861 20374 12871 20430
rect 12927 20374 12995 20430
rect 13051 20374 13119 20430
rect 13175 20374 13243 20430
rect 13299 20374 13367 20430
rect 13423 20374 13491 20430
rect 13547 20374 13615 20430
rect 13671 20374 13739 20430
rect 13795 20374 13863 20430
rect 13919 20374 13987 20430
rect 14043 20374 14111 20430
rect 14167 20374 14235 20430
rect 14291 20374 14359 20430
rect 14415 20374 14483 20430
rect 14539 20374 14607 20430
rect 14663 20374 14673 20430
rect 12861 20306 14673 20374
rect 12861 20250 12871 20306
rect 12927 20250 12995 20306
rect 13051 20250 13119 20306
rect 13175 20250 13243 20306
rect 13299 20250 13367 20306
rect 13423 20250 13491 20306
rect 13547 20250 13615 20306
rect 13671 20250 13739 20306
rect 13795 20250 13863 20306
rect 13919 20250 13987 20306
rect 14043 20250 14111 20306
rect 14167 20250 14235 20306
rect 14291 20250 14359 20306
rect 14415 20250 14483 20306
rect 14539 20250 14607 20306
rect 14663 20250 14673 20306
rect 12861 20182 14673 20250
rect 12861 20126 12871 20182
rect 12927 20126 12995 20182
rect 13051 20126 13119 20182
rect 13175 20126 13243 20182
rect 13299 20126 13367 20182
rect 13423 20126 13491 20182
rect 13547 20126 13615 20182
rect 13671 20126 13739 20182
rect 13795 20126 13863 20182
rect 13919 20126 13987 20182
rect 14043 20126 14111 20182
rect 14167 20126 14235 20182
rect 14291 20126 14359 20182
rect 14415 20126 14483 20182
rect 14539 20126 14607 20182
rect 14663 20126 14673 20182
rect 12861 20058 14673 20126
rect 12861 20002 12871 20058
rect 12927 20002 12995 20058
rect 13051 20002 13119 20058
rect 13175 20002 13243 20058
rect 13299 20002 13367 20058
rect 13423 20002 13491 20058
rect 13547 20002 13615 20058
rect 13671 20002 13739 20058
rect 13795 20002 13863 20058
rect 13919 20002 13987 20058
rect 14043 20002 14111 20058
rect 14167 20002 14235 20058
rect 14291 20002 14359 20058
rect 14415 20002 14483 20058
rect 14539 20002 14607 20058
rect 14663 20002 14673 20058
rect 12861 19934 14673 20002
rect 12861 19878 12871 19934
rect 12927 19878 12995 19934
rect 13051 19878 13119 19934
rect 13175 19878 13243 19934
rect 13299 19878 13367 19934
rect 13423 19878 13491 19934
rect 13547 19878 13615 19934
rect 13671 19878 13739 19934
rect 13795 19878 13863 19934
rect 13919 19878 13987 19934
rect 14043 19878 14111 19934
rect 14167 19878 14235 19934
rect 14291 19878 14359 19934
rect 14415 19878 14483 19934
rect 14539 19878 14607 19934
rect 14663 19878 14673 19934
rect 12861 19810 14673 19878
rect 12861 19754 12871 19810
rect 12927 19754 12995 19810
rect 13051 19754 13119 19810
rect 13175 19754 13243 19810
rect 13299 19754 13367 19810
rect 13423 19754 13491 19810
rect 13547 19754 13615 19810
rect 13671 19754 13739 19810
rect 13795 19754 13863 19810
rect 13919 19754 13987 19810
rect 14043 19754 14111 19810
rect 14167 19754 14235 19810
rect 14291 19754 14359 19810
rect 14415 19754 14483 19810
rect 14539 19754 14607 19810
rect 14663 19754 14673 19810
rect 12861 19686 14673 19754
rect 12861 19630 12871 19686
rect 12927 19630 12995 19686
rect 13051 19630 13119 19686
rect 13175 19630 13243 19686
rect 13299 19630 13367 19686
rect 13423 19630 13491 19686
rect 13547 19630 13615 19686
rect 13671 19630 13739 19686
rect 13795 19630 13863 19686
rect 13919 19630 13987 19686
rect 14043 19630 14111 19686
rect 14167 19630 14235 19686
rect 14291 19630 14359 19686
rect 14415 19630 14483 19686
rect 14539 19630 14607 19686
rect 14663 19630 14673 19686
rect 12861 19562 14673 19630
rect 12861 19506 12871 19562
rect 12927 19506 12995 19562
rect 13051 19506 13119 19562
rect 13175 19506 13243 19562
rect 13299 19506 13367 19562
rect 13423 19506 13491 19562
rect 13547 19506 13615 19562
rect 13671 19506 13739 19562
rect 13795 19506 13863 19562
rect 13919 19506 13987 19562
rect 14043 19506 14111 19562
rect 14167 19506 14235 19562
rect 14291 19506 14359 19562
rect 14415 19506 14483 19562
rect 14539 19506 14607 19562
rect 14663 19506 14673 19562
rect 12861 19438 14673 19506
rect 12861 19382 12871 19438
rect 12927 19382 12995 19438
rect 13051 19382 13119 19438
rect 13175 19382 13243 19438
rect 13299 19382 13367 19438
rect 13423 19382 13491 19438
rect 13547 19382 13615 19438
rect 13671 19382 13739 19438
rect 13795 19382 13863 19438
rect 13919 19382 13987 19438
rect 14043 19382 14111 19438
rect 14167 19382 14235 19438
rect 14291 19382 14359 19438
rect 14415 19382 14483 19438
rect 14539 19382 14607 19438
rect 14663 19382 14673 19438
rect 12861 19314 14673 19382
rect 12861 19258 12871 19314
rect 12927 19258 12995 19314
rect 13051 19258 13119 19314
rect 13175 19258 13243 19314
rect 13299 19258 13367 19314
rect 13423 19258 13491 19314
rect 13547 19258 13615 19314
rect 13671 19258 13739 19314
rect 13795 19258 13863 19314
rect 13919 19258 13987 19314
rect 14043 19258 14111 19314
rect 14167 19258 14235 19314
rect 14291 19258 14359 19314
rect 14415 19258 14483 19314
rect 14539 19258 14607 19314
rect 14663 19258 14673 19314
rect 12861 19190 14673 19258
rect 12861 19134 12871 19190
rect 12927 19134 12995 19190
rect 13051 19134 13119 19190
rect 13175 19134 13243 19190
rect 13299 19134 13367 19190
rect 13423 19134 13491 19190
rect 13547 19134 13615 19190
rect 13671 19134 13739 19190
rect 13795 19134 13863 19190
rect 13919 19134 13987 19190
rect 14043 19134 14111 19190
rect 14167 19134 14235 19190
rect 14291 19134 14359 19190
rect 14415 19134 14483 19190
rect 14539 19134 14607 19190
rect 14663 19134 14673 19190
rect 12861 19066 14673 19134
rect 12861 19010 12871 19066
rect 12927 19010 12995 19066
rect 13051 19010 13119 19066
rect 13175 19010 13243 19066
rect 13299 19010 13367 19066
rect 13423 19010 13491 19066
rect 13547 19010 13615 19066
rect 13671 19010 13739 19066
rect 13795 19010 13863 19066
rect 13919 19010 13987 19066
rect 14043 19010 14111 19066
rect 14167 19010 14235 19066
rect 14291 19010 14359 19066
rect 14415 19010 14483 19066
rect 14539 19010 14607 19066
rect 14663 19010 14673 19066
rect 12861 18942 14673 19010
rect 12861 18886 12871 18942
rect 12927 18886 12995 18942
rect 13051 18886 13119 18942
rect 13175 18886 13243 18942
rect 13299 18886 13367 18942
rect 13423 18886 13491 18942
rect 13547 18886 13615 18942
rect 13671 18886 13739 18942
rect 13795 18886 13863 18942
rect 13919 18886 13987 18942
rect 14043 18886 14111 18942
rect 14167 18886 14235 18942
rect 14291 18886 14359 18942
rect 14415 18886 14483 18942
rect 14539 18886 14607 18942
rect 14663 18886 14673 18942
rect 12861 18818 14673 18886
rect 12861 18762 12871 18818
rect 12927 18762 12995 18818
rect 13051 18762 13119 18818
rect 13175 18762 13243 18818
rect 13299 18762 13367 18818
rect 13423 18762 13491 18818
rect 13547 18762 13615 18818
rect 13671 18762 13739 18818
rect 13795 18762 13863 18818
rect 13919 18762 13987 18818
rect 14043 18762 14111 18818
rect 14167 18762 14235 18818
rect 14291 18762 14359 18818
rect 14415 18762 14483 18818
rect 14539 18762 14607 18818
rect 14663 18762 14673 18818
rect 12861 18694 14673 18762
rect 12861 18638 12871 18694
rect 12927 18638 12995 18694
rect 13051 18638 13119 18694
rect 13175 18638 13243 18694
rect 13299 18638 13367 18694
rect 13423 18638 13491 18694
rect 13547 18638 13615 18694
rect 13671 18638 13739 18694
rect 13795 18638 13863 18694
rect 13919 18638 13987 18694
rect 14043 18638 14111 18694
rect 14167 18638 14235 18694
rect 14291 18638 14359 18694
rect 14415 18638 14483 18694
rect 14539 18638 14607 18694
rect 14663 18638 14673 18694
rect 12861 18570 14673 18638
rect 12861 18514 12871 18570
rect 12927 18514 12995 18570
rect 13051 18514 13119 18570
rect 13175 18514 13243 18570
rect 13299 18514 13367 18570
rect 13423 18514 13491 18570
rect 13547 18514 13615 18570
rect 13671 18514 13739 18570
rect 13795 18514 13863 18570
rect 13919 18514 13987 18570
rect 14043 18514 14111 18570
rect 14167 18514 14235 18570
rect 14291 18514 14359 18570
rect 14415 18514 14483 18570
rect 14539 18514 14607 18570
rect 14663 18514 14673 18570
rect 12861 18446 14673 18514
rect 12861 18390 12871 18446
rect 12927 18390 12995 18446
rect 13051 18390 13119 18446
rect 13175 18390 13243 18446
rect 13299 18390 13367 18446
rect 13423 18390 13491 18446
rect 13547 18390 13615 18446
rect 13671 18390 13739 18446
rect 13795 18390 13863 18446
rect 13919 18390 13987 18446
rect 14043 18390 14111 18446
rect 14167 18390 14235 18446
rect 14291 18390 14359 18446
rect 14415 18390 14483 18446
rect 14539 18390 14607 18446
rect 14663 18390 14673 18446
rect 12861 18322 14673 18390
rect 12861 18266 12871 18322
rect 12927 18266 12995 18322
rect 13051 18266 13119 18322
rect 13175 18266 13243 18322
rect 13299 18266 13367 18322
rect 13423 18266 13491 18322
rect 13547 18266 13615 18322
rect 13671 18266 13739 18322
rect 13795 18266 13863 18322
rect 13919 18266 13987 18322
rect 14043 18266 14111 18322
rect 14167 18266 14235 18322
rect 14291 18266 14359 18322
rect 14415 18266 14483 18322
rect 14539 18266 14607 18322
rect 14663 18266 14673 18322
rect 12861 18198 14673 18266
rect 12861 18142 12871 18198
rect 12927 18142 12995 18198
rect 13051 18142 13119 18198
rect 13175 18142 13243 18198
rect 13299 18142 13367 18198
rect 13423 18142 13491 18198
rect 13547 18142 13615 18198
rect 13671 18142 13739 18198
rect 13795 18142 13863 18198
rect 13919 18142 13987 18198
rect 14043 18142 14111 18198
rect 14167 18142 14235 18198
rect 14291 18142 14359 18198
rect 14415 18142 14483 18198
rect 14539 18142 14607 18198
rect 14663 18142 14673 18198
rect 12861 18074 14673 18142
rect 12861 18018 12871 18074
rect 12927 18018 12995 18074
rect 13051 18018 13119 18074
rect 13175 18018 13243 18074
rect 13299 18018 13367 18074
rect 13423 18018 13491 18074
rect 13547 18018 13615 18074
rect 13671 18018 13739 18074
rect 13795 18018 13863 18074
rect 13919 18018 13987 18074
rect 14043 18018 14111 18074
rect 14167 18018 14235 18074
rect 14291 18018 14359 18074
rect 14415 18018 14483 18074
rect 14539 18018 14607 18074
rect 14663 18018 14673 18074
rect 12861 17950 14673 18018
rect 12861 17894 12871 17950
rect 12927 17894 12995 17950
rect 13051 17894 13119 17950
rect 13175 17894 13243 17950
rect 13299 17894 13367 17950
rect 13423 17894 13491 17950
rect 13547 17894 13615 17950
rect 13671 17894 13739 17950
rect 13795 17894 13863 17950
rect 13919 17894 13987 17950
rect 14043 17894 14111 17950
rect 14167 17894 14235 17950
rect 14291 17894 14359 17950
rect 14415 17894 14483 17950
rect 14539 17894 14607 17950
rect 14663 17894 14673 17950
rect 12861 17826 14673 17894
rect 12861 17770 12871 17826
rect 12927 17770 12995 17826
rect 13051 17770 13119 17826
rect 13175 17770 13243 17826
rect 13299 17770 13367 17826
rect 13423 17770 13491 17826
rect 13547 17770 13615 17826
rect 13671 17770 13739 17826
rect 13795 17770 13863 17826
rect 13919 17770 13987 17826
rect 14043 17770 14111 17826
rect 14167 17770 14235 17826
rect 14291 17770 14359 17826
rect 14415 17770 14483 17826
rect 14539 17770 14607 17826
rect 14663 17770 14673 17826
rect 12861 17702 14673 17770
rect 12861 17646 12871 17702
rect 12927 17646 12995 17702
rect 13051 17646 13119 17702
rect 13175 17646 13243 17702
rect 13299 17646 13367 17702
rect 13423 17646 13491 17702
rect 13547 17646 13615 17702
rect 13671 17646 13739 17702
rect 13795 17646 13863 17702
rect 13919 17646 13987 17702
rect 14043 17646 14111 17702
rect 14167 17646 14235 17702
rect 14291 17646 14359 17702
rect 14415 17646 14483 17702
rect 14539 17646 14607 17702
rect 14663 17646 14673 17702
rect 12861 17636 14673 17646
rect 305 17354 2117 17364
rect 305 17298 315 17354
rect 371 17298 439 17354
rect 495 17298 563 17354
rect 619 17298 687 17354
rect 743 17298 811 17354
rect 867 17298 935 17354
rect 991 17298 1059 17354
rect 1115 17298 1183 17354
rect 1239 17298 1307 17354
rect 1363 17298 1431 17354
rect 1487 17298 1555 17354
rect 1611 17298 1679 17354
rect 1735 17298 1803 17354
rect 1859 17298 1927 17354
rect 1983 17298 2051 17354
rect 2107 17298 2117 17354
rect 305 17230 2117 17298
rect 305 17174 315 17230
rect 371 17174 439 17230
rect 495 17174 563 17230
rect 619 17174 687 17230
rect 743 17174 811 17230
rect 867 17174 935 17230
rect 991 17174 1059 17230
rect 1115 17174 1183 17230
rect 1239 17174 1307 17230
rect 1363 17174 1431 17230
rect 1487 17174 1555 17230
rect 1611 17174 1679 17230
rect 1735 17174 1803 17230
rect 1859 17174 1927 17230
rect 1983 17174 2051 17230
rect 2107 17174 2117 17230
rect 305 17106 2117 17174
rect 305 17050 315 17106
rect 371 17050 439 17106
rect 495 17050 563 17106
rect 619 17050 687 17106
rect 743 17050 811 17106
rect 867 17050 935 17106
rect 991 17050 1059 17106
rect 1115 17050 1183 17106
rect 1239 17050 1307 17106
rect 1363 17050 1431 17106
rect 1487 17050 1555 17106
rect 1611 17050 1679 17106
rect 1735 17050 1803 17106
rect 1859 17050 1927 17106
rect 1983 17050 2051 17106
rect 2107 17050 2117 17106
rect 305 16982 2117 17050
rect 305 16926 315 16982
rect 371 16926 439 16982
rect 495 16926 563 16982
rect 619 16926 687 16982
rect 743 16926 811 16982
rect 867 16926 935 16982
rect 991 16926 1059 16982
rect 1115 16926 1183 16982
rect 1239 16926 1307 16982
rect 1363 16926 1431 16982
rect 1487 16926 1555 16982
rect 1611 16926 1679 16982
rect 1735 16926 1803 16982
rect 1859 16926 1927 16982
rect 1983 16926 2051 16982
rect 2107 16926 2117 16982
rect 305 16858 2117 16926
rect 305 16802 315 16858
rect 371 16802 439 16858
rect 495 16802 563 16858
rect 619 16802 687 16858
rect 743 16802 811 16858
rect 867 16802 935 16858
rect 991 16802 1059 16858
rect 1115 16802 1183 16858
rect 1239 16802 1307 16858
rect 1363 16802 1431 16858
rect 1487 16802 1555 16858
rect 1611 16802 1679 16858
rect 1735 16802 1803 16858
rect 1859 16802 1927 16858
rect 1983 16802 2051 16858
rect 2107 16802 2117 16858
rect 305 16734 2117 16802
rect 305 16678 315 16734
rect 371 16678 439 16734
rect 495 16678 563 16734
rect 619 16678 687 16734
rect 743 16678 811 16734
rect 867 16678 935 16734
rect 991 16678 1059 16734
rect 1115 16678 1183 16734
rect 1239 16678 1307 16734
rect 1363 16678 1431 16734
rect 1487 16678 1555 16734
rect 1611 16678 1679 16734
rect 1735 16678 1803 16734
rect 1859 16678 1927 16734
rect 1983 16678 2051 16734
rect 2107 16678 2117 16734
rect 305 16610 2117 16678
rect 305 16554 315 16610
rect 371 16554 439 16610
rect 495 16554 563 16610
rect 619 16554 687 16610
rect 743 16554 811 16610
rect 867 16554 935 16610
rect 991 16554 1059 16610
rect 1115 16554 1183 16610
rect 1239 16554 1307 16610
rect 1363 16554 1431 16610
rect 1487 16554 1555 16610
rect 1611 16554 1679 16610
rect 1735 16554 1803 16610
rect 1859 16554 1927 16610
rect 1983 16554 2051 16610
rect 2107 16554 2117 16610
rect 305 16486 2117 16554
rect 305 16430 315 16486
rect 371 16430 439 16486
rect 495 16430 563 16486
rect 619 16430 687 16486
rect 743 16430 811 16486
rect 867 16430 935 16486
rect 991 16430 1059 16486
rect 1115 16430 1183 16486
rect 1239 16430 1307 16486
rect 1363 16430 1431 16486
rect 1487 16430 1555 16486
rect 1611 16430 1679 16486
rect 1735 16430 1803 16486
rect 1859 16430 1927 16486
rect 1983 16430 2051 16486
rect 2107 16430 2117 16486
rect 305 16362 2117 16430
rect 305 16306 315 16362
rect 371 16306 439 16362
rect 495 16306 563 16362
rect 619 16306 687 16362
rect 743 16306 811 16362
rect 867 16306 935 16362
rect 991 16306 1059 16362
rect 1115 16306 1183 16362
rect 1239 16306 1307 16362
rect 1363 16306 1431 16362
rect 1487 16306 1555 16362
rect 1611 16306 1679 16362
rect 1735 16306 1803 16362
rect 1859 16306 1927 16362
rect 1983 16306 2051 16362
rect 2107 16306 2117 16362
rect 305 16238 2117 16306
rect 305 16182 315 16238
rect 371 16182 439 16238
rect 495 16182 563 16238
rect 619 16182 687 16238
rect 743 16182 811 16238
rect 867 16182 935 16238
rect 991 16182 1059 16238
rect 1115 16182 1183 16238
rect 1239 16182 1307 16238
rect 1363 16182 1431 16238
rect 1487 16182 1555 16238
rect 1611 16182 1679 16238
rect 1735 16182 1803 16238
rect 1859 16182 1927 16238
rect 1983 16182 2051 16238
rect 2107 16182 2117 16238
rect 305 16114 2117 16182
rect 305 16058 315 16114
rect 371 16058 439 16114
rect 495 16058 563 16114
rect 619 16058 687 16114
rect 743 16058 811 16114
rect 867 16058 935 16114
rect 991 16058 1059 16114
rect 1115 16058 1183 16114
rect 1239 16058 1307 16114
rect 1363 16058 1431 16114
rect 1487 16058 1555 16114
rect 1611 16058 1679 16114
rect 1735 16058 1803 16114
rect 1859 16058 1927 16114
rect 1983 16058 2051 16114
rect 2107 16058 2117 16114
rect 305 15990 2117 16058
rect 305 15934 315 15990
rect 371 15934 439 15990
rect 495 15934 563 15990
rect 619 15934 687 15990
rect 743 15934 811 15990
rect 867 15934 935 15990
rect 991 15934 1059 15990
rect 1115 15934 1183 15990
rect 1239 15934 1307 15990
rect 1363 15934 1431 15990
rect 1487 15934 1555 15990
rect 1611 15934 1679 15990
rect 1735 15934 1803 15990
rect 1859 15934 1927 15990
rect 1983 15934 2051 15990
rect 2107 15934 2117 15990
rect 305 15866 2117 15934
rect 305 15810 315 15866
rect 371 15810 439 15866
rect 495 15810 563 15866
rect 619 15810 687 15866
rect 743 15810 811 15866
rect 867 15810 935 15866
rect 991 15810 1059 15866
rect 1115 15810 1183 15866
rect 1239 15810 1307 15866
rect 1363 15810 1431 15866
rect 1487 15810 1555 15866
rect 1611 15810 1679 15866
rect 1735 15810 1803 15866
rect 1859 15810 1927 15866
rect 1983 15810 2051 15866
rect 2107 15810 2117 15866
rect 305 15742 2117 15810
rect 305 15686 315 15742
rect 371 15686 439 15742
rect 495 15686 563 15742
rect 619 15686 687 15742
rect 743 15686 811 15742
rect 867 15686 935 15742
rect 991 15686 1059 15742
rect 1115 15686 1183 15742
rect 1239 15686 1307 15742
rect 1363 15686 1431 15742
rect 1487 15686 1555 15742
rect 1611 15686 1679 15742
rect 1735 15686 1803 15742
rect 1859 15686 1927 15742
rect 1983 15686 2051 15742
rect 2107 15686 2117 15742
rect 305 15618 2117 15686
rect 305 15562 315 15618
rect 371 15562 439 15618
rect 495 15562 563 15618
rect 619 15562 687 15618
rect 743 15562 811 15618
rect 867 15562 935 15618
rect 991 15562 1059 15618
rect 1115 15562 1183 15618
rect 1239 15562 1307 15618
rect 1363 15562 1431 15618
rect 1487 15562 1555 15618
rect 1611 15562 1679 15618
rect 1735 15562 1803 15618
rect 1859 15562 1927 15618
rect 1983 15562 2051 15618
rect 2107 15562 2117 15618
rect 305 15494 2117 15562
rect 305 15438 315 15494
rect 371 15438 439 15494
rect 495 15438 563 15494
rect 619 15438 687 15494
rect 743 15438 811 15494
rect 867 15438 935 15494
rect 991 15438 1059 15494
rect 1115 15438 1183 15494
rect 1239 15438 1307 15494
rect 1363 15438 1431 15494
rect 1487 15438 1555 15494
rect 1611 15438 1679 15494
rect 1735 15438 1803 15494
rect 1859 15438 1927 15494
rect 1983 15438 2051 15494
rect 2107 15438 2117 15494
rect 305 15370 2117 15438
rect 305 15314 315 15370
rect 371 15314 439 15370
rect 495 15314 563 15370
rect 619 15314 687 15370
rect 743 15314 811 15370
rect 867 15314 935 15370
rect 991 15314 1059 15370
rect 1115 15314 1183 15370
rect 1239 15314 1307 15370
rect 1363 15314 1431 15370
rect 1487 15314 1555 15370
rect 1611 15314 1679 15370
rect 1735 15314 1803 15370
rect 1859 15314 1927 15370
rect 1983 15314 2051 15370
rect 2107 15314 2117 15370
rect 305 15246 2117 15314
rect 305 15190 315 15246
rect 371 15190 439 15246
rect 495 15190 563 15246
rect 619 15190 687 15246
rect 743 15190 811 15246
rect 867 15190 935 15246
rect 991 15190 1059 15246
rect 1115 15190 1183 15246
rect 1239 15190 1307 15246
rect 1363 15190 1431 15246
rect 1487 15190 1555 15246
rect 1611 15190 1679 15246
rect 1735 15190 1803 15246
rect 1859 15190 1927 15246
rect 1983 15190 2051 15246
rect 2107 15190 2117 15246
rect 305 15122 2117 15190
rect 305 15066 315 15122
rect 371 15066 439 15122
rect 495 15066 563 15122
rect 619 15066 687 15122
rect 743 15066 811 15122
rect 867 15066 935 15122
rect 991 15066 1059 15122
rect 1115 15066 1183 15122
rect 1239 15066 1307 15122
rect 1363 15066 1431 15122
rect 1487 15066 1555 15122
rect 1611 15066 1679 15122
rect 1735 15066 1803 15122
rect 1859 15066 1927 15122
rect 1983 15066 2051 15122
rect 2107 15066 2117 15122
rect 305 14998 2117 15066
rect 305 14942 315 14998
rect 371 14942 439 14998
rect 495 14942 563 14998
rect 619 14942 687 14998
rect 743 14942 811 14998
rect 867 14942 935 14998
rect 991 14942 1059 14998
rect 1115 14942 1183 14998
rect 1239 14942 1307 14998
rect 1363 14942 1431 14998
rect 1487 14942 1555 14998
rect 1611 14942 1679 14998
rect 1735 14942 1803 14998
rect 1859 14942 1927 14998
rect 1983 14942 2051 14998
rect 2107 14942 2117 14998
rect 305 14874 2117 14942
rect 305 14818 315 14874
rect 371 14818 439 14874
rect 495 14818 563 14874
rect 619 14818 687 14874
rect 743 14818 811 14874
rect 867 14818 935 14874
rect 991 14818 1059 14874
rect 1115 14818 1183 14874
rect 1239 14818 1307 14874
rect 1363 14818 1431 14874
rect 1487 14818 1555 14874
rect 1611 14818 1679 14874
rect 1735 14818 1803 14874
rect 1859 14818 1927 14874
rect 1983 14818 2051 14874
rect 2107 14818 2117 14874
rect 305 14750 2117 14818
rect 305 14694 315 14750
rect 371 14694 439 14750
rect 495 14694 563 14750
rect 619 14694 687 14750
rect 743 14694 811 14750
rect 867 14694 935 14750
rect 991 14694 1059 14750
rect 1115 14694 1183 14750
rect 1239 14694 1307 14750
rect 1363 14694 1431 14750
rect 1487 14694 1555 14750
rect 1611 14694 1679 14750
rect 1735 14694 1803 14750
rect 1859 14694 1927 14750
rect 1983 14694 2051 14750
rect 2107 14694 2117 14750
rect 305 14626 2117 14694
rect 305 14570 315 14626
rect 371 14570 439 14626
rect 495 14570 563 14626
rect 619 14570 687 14626
rect 743 14570 811 14626
rect 867 14570 935 14626
rect 991 14570 1059 14626
rect 1115 14570 1183 14626
rect 1239 14570 1307 14626
rect 1363 14570 1431 14626
rect 1487 14570 1555 14626
rect 1611 14570 1679 14626
rect 1735 14570 1803 14626
rect 1859 14570 1927 14626
rect 1983 14570 2051 14626
rect 2107 14570 2117 14626
rect 305 14502 2117 14570
rect 305 14446 315 14502
rect 371 14446 439 14502
rect 495 14446 563 14502
rect 619 14446 687 14502
rect 743 14446 811 14502
rect 867 14446 935 14502
rect 991 14446 1059 14502
rect 1115 14446 1183 14502
rect 1239 14446 1307 14502
rect 1363 14446 1431 14502
rect 1487 14446 1555 14502
rect 1611 14446 1679 14502
rect 1735 14446 1803 14502
rect 1859 14446 1927 14502
rect 1983 14446 2051 14502
rect 2107 14446 2117 14502
rect 305 14436 2117 14446
rect 2798 17354 4734 17364
rect 2798 17298 2808 17354
rect 2864 17298 2932 17354
rect 2988 17298 3056 17354
rect 3112 17298 3180 17354
rect 3236 17298 3304 17354
rect 3360 17298 3428 17354
rect 3484 17298 3552 17354
rect 3608 17298 3676 17354
rect 3732 17298 3800 17354
rect 3856 17298 3924 17354
rect 3980 17298 4048 17354
rect 4104 17298 4172 17354
rect 4228 17298 4296 17354
rect 4352 17298 4420 17354
rect 4476 17298 4544 17354
rect 4600 17298 4668 17354
rect 4724 17298 4734 17354
rect 2798 17230 4734 17298
rect 2798 17174 2808 17230
rect 2864 17174 2932 17230
rect 2988 17174 3056 17230
rect 3112 17174 3180 17230
rect 3236 17174 3304 17230
rect 3360 17174 3428 17230
rect 3484 17174 3552 17230
rect 3608 17174 3676 17230
rect 3732 17174 3800 17230
rect 3856 17174 3924 17230
rect 3980 17174 4048 17230
rect 4104 17174 4172 17230
rect 4228 17174 4296 17230
rect 4352 17174 4420 17230
rect 4476 17174 4544 17230
rect 4600 17174 4668 17230
rect 4724 17174 4734 17230
rect 2798 17106 4734 17174
rect 2798 17050 2808 17106
rect 2864 17050 2932 17106
rect 2988 17050 3056 17106
rect 3112 17050 3180 17106
rect 3236 17050 3304 17106
rect 3360 17050 3428 17106
rect 3484 17050 3552 17106
rect 3608 17050 3676 17106
rect 3732 17050 3800 17106
rect 3856 17050 3924 17106
rect 3980 17050 4048 17106
rect 4104 17050 4172 17106
rect 4228 17050 4296 17106
rect 4352 17050 4420 17106
rect 4476 17050 4544 17106
rect 4600 17050 4668 17106
rect 4724 17050 4734 17106
rect 2798 16982 4734 17050
rect 2798 16926 2808 16982
rect 2864 16926 2932 16982
rect 2988 16926 3056 16982
rect 3112 16926 3180 16982
rect 3236 16926 3304 16982
rect 3360 16926 3428 16982
rect 3484 16926 3552 16982
rect 3608 16926 3676 16982
rect 3732 16926 3800 16982
rect 3856 16926 3924 16982
rect 3980 16926 4048 16982
rect 4104 16926 4172 16982
rect 4228 16926 4296 16982
rect 4352 16926 4420 16982
rect 4476 16926 4544 16982
rect 4600 16926 4668 16982
rect 4724 16926 4734 16982
rect 2798 16858 4734 16926
rect 2798 16802 2808 16858
rect 2864 16802 2932 16858
rect 2988 16802 3056 16858
rect 3112 16802 3180 16858
rect 3236 16802 3304 16858
rect 3360 16802 3428 16858
rect 3484 16802 3552 16858
rect 3608 16802 3676 16858
rect 3732 16802 3800 16858
rect 3856 16802 3924 16858
rect 3980 16802 4048 16858
rect 4104 16802 4172 16858
rect 4228 16802 4296 16858
rect 4352 16802 4420 16858
rect 4476 16802 4544 16858
rect 4600 16802 4668 16858
rect 4724 16802 4734 16858
rect 2798 16734 4734 16802
rect 2798 16678 2808 16734
rect 2864 16678 2932 16734
rect 2988 16678 3056 16734
rect 3112 16678 3180 16734
rect 3236 16678 3304 16734
rect 3360 16678 3428 16734
rect 3484 16678 3552 16734
rect 3608 16678 3676 16734
rect 3732 16678 3800 16734
rect 3856 16678 3924 16734
rect 3980 16678 4048 16734
rect 4104 16678 4172 16734
rect 4228 16678 4296 16734
rect 4352 16678 4420 16734
rect 4476 16678 4544 16734
rect 4600 16678 4668 16734
rect 4724 16678 4734 16734
rect 2798 16610 4734 16678
rect 2798 16554 2808 16610
rect 2864 16554 2932 16610
rect 2988 16554 3056 16610
rect 3112 16554 3180 16610
rect 3236 16554 3304 16610
rect 3360 16554 3428 16610
rect 3484 16554 3552 16610
rect 3608 16554 3676 16610
rect 3732 16554 3800 16610
rect 3856 16554 3924 16610
rect 3980 16554 4048 16610
rect 4104 16554 4172 16610
rect 4228 16554 4296 16610
rect 4352 16554 4420 16610
rect 4476 16554 4544 16610
rect 4600 16554 4668 16610
rect 4724 16554 4734 16610
rect 2798 16486 4734 16554
rect 2798 16430 2808 16486
rect 2864 16430 2932 16486
rect 2988 16430 3056 16486
rect 3112 16430 3180 16486
rect 3236 16430 3304 16486
rect 3360 16430 3428 16486
rect 3484 16430 3552 16486
rect 3608 16430 3676 16486
rect 3732 16430 3800 16486
rect 3856 16430 3924 16486
rect 3980 16430 4048 16486
rect 4104 16430 4172 16486
rect 4228 16430 4296 16486
rect 4352 16430 4420 16486
rect 4476 16430 4544 16486
rect 4600 16430 4668 16486
rect 4724 16430 4734 16486
rect 2798 16362 4734 16430
rect 2798 16306 2808 16362
rect 2864 16306 2932 16362
rect 2988 16306 3056 16362
rect 3112 16306 3180 16362
rect 3236 16306 3304 16362
rect 3360 16306 3428 16362
rect 3484 16306 3552 16362
rect 3608 16306 3676 16362
rect 3732 16306 3800 16362
rect 3856 16306 3924 16362
rect 3980 16306 4048 16362
rect 4104 16306 4172 16362
rect 4228 16306 4296 16362
rect 4352 16306 4420 16362
rect 4476 16306 4544 16362
rect 4600 16306 4668 16362
rect 4724 16306 4734 16362
rect 2798 16238 4734 16306
rect 2798 16182 2808 16238
rect 2864 16182 2932 16238
rect 2988 16182 3056 16238
rect 3112 16182 3180 16238
rect 3236 16182 3304 16238
rect 3360 16182 3428 16238
rect 3484 16182 3552 16238
rect 3608 16182 3676 16238
rect 3732 16182 3800 16238
rect 3856 16182 3924 16238
rect 3980 16182 4048 16238
rect 4104 16182 4172 16238
rect 4228 16182 4296 16238
rect 4352 16182 4420 16238
rect 4476 16182 4544 16238
rect 4600 16182 4668 16238
rect 4724 16182 4734 16238
rect 2798 16114 4734 16182
rect 2798 16058 2808 16114
rect 2864 16058 2932 16114
rect 2988 16058 3056 16114
rect 3112 16058 3180 16114
rect 3236 16058 3304 16114
rect 3360 16058 3428 16114
rect 3484 16058 3552 16114
rect 3608 16058 3676 16114
rect 3732 16058 3800 16114
rect 3856 16058 3924 16114
rect 3980 16058 4048 16114
rect 4104 16058 4172 16114
rect 4228 16058 4296 16114
rect 4352 16058 4420 16114
rect 4476 16058 4544 16114
rect 4600 16058 4668 16114
rect 4724 16058 4734 16114
rect 2798 15990 4734 16058
rect 2798 15934 2808 15990
rect 2864 15934 2932 15990
rect 2988 15934 3056 15990
rect 3112 15934 3180 15990
rect 3236 15934 3304 15990
rect 3360 15934 3428 15990
rect 3484 15934 3552 15990
rect 3608 15934 3676 15990
rect 3732 15934 3800 15990
rect 3856 15934 3924 15990
rect 3980 15934 4048 15990
rect 4104 15934 4172 15990
rect 4228 15934 4296 15990
rect 4352 15934 4420 15990
rect 4476 15934 4544 15990
rect 4600 15934 4668 15990
rect 4724 15934 4734 15990
rect 2798 15866 4734 15934
rect 2798 15810 2808 15866
rect 2864 15810 2932 15866
rect 2988 15810 3056 15866
rect 3112 15810 3180 15866
rect 3236 15810 3304 15866
rect 3360 15810 3428 15866
rect 3484 15810 3552 15866
rect 3608 15810 3676 15866
rect 3732 15810 3800 15866
rect 3856 15810 3924 15866
rect 3980 15810 4048 15866
rect 4104 15810 4172 15866
rect 4228 15810 4296 15866
rect 4352 15810 4420 15866
rect 4476 15810 4544 15866
rect 4600 15810 4668 15866
rect 4724 15810 4734 15866
rect 2798 15742 4734 15810
rect 2798 15686 2808 15742
rect 2864 15686 2932 15742
rect 2988 15686 3056 15742
rect 3112 15686 3180 15742
rect 3236 15686 3304 15742
rect 3360 15686 3428 15742
rect 3484 15686 3552 15742
rect 3608 15686 3676 15742
rect 3732 15686 3800 15742
rect 3856 15686 3924 15742
rect 3980 15686 4048 15742
rect 4104 15686 4172 15742
rect 4228 15686 4296 15742
rect 4352 15686 4420 15742
rect 4476 15686 4544 15742
rect 4600 15686 4668 15742
rect 4724 15686 4734 15742
rect 2798 15618 4734 15686
rect 2798 15562 2808 15618
rect 2864 15562 2932 15618
rect 2988 15562 3056 15618
rect 3112 15562 3180 15618
rect 3236 15562 3304 15618
rect 3360 15562 3428 15618
rect 3484 15562 3552 15618
rect 3608 15562 3676 15618
rect 3732 15562 3800 15618
rect 3856 15562 3924 15618
rect 3980 15562 4048 15618
rect 4104 15562 4172 15618
rect 4228 15562 4296 15618
rect 4352 15562 4420 15618
rect 4476 15562 4544 15618
rect 4600 15562 4668 15618
rect 4724 15562 4734 15618
rect 2798 15494 4734 15562
rect 2798 15438 2808 15494
rect 2864 15438 2932 15494
rect 2988 15438 3056 15494
rect 3112 15438 3180 15494
rect 3236 15438 3304 15494
rect 3360 15438 3428 15494
rect 3484 15438 3552 15494
rect 3608 15438 3676 15494
rect 3732 15438 3800 15494
rect 3856 15438 3924 15494
rect 3980 15438 4048 15494
rect 4104 15438 4172 15494
rect 4228 15438 4296 15494
rect 4352 15438 4420 15494
rect 4476 15438 4544 15494
rect 4600 15438 4668 15494
rect 4724 15438 4734 15494
rect 2798 15370 4734 15438
rect 2798 15314 2808 15370
rect 2864 15314 2932 15370
rect 2988 15314 3056 15370
rect 3112 15314 3180 15370
rect 3236 15314 3304 15370
rect 3360 15314 3428 15370
rect 3484 15314 3552 15370
rect 3608 15314 3676 15370
rect 3732 15314 3800 15370
rect 3856 15314 3924 15370
rect 3980 15314 4048 15370
rect 4104 15314 4172 15370
rect 4228 15314 4296 15370
rect 4352 15314 4420 15370
rect 4476 15314 4544 15370
rect 4600 15314 4668 15370
rect 4724 15314 4734 15370
rect 2798 15246 4734 15314
rect 2798 15190 2808 15246
rect 2864 15190 2932 15246
rect 2988 15190 3056 15246
rect 3112 15190 3180 15246
rect 3236 15190 3304 15246
rect 3360 15190 3428 15246
rect 3484 15190 3552 15246
rect 3608 15190 3676 15246
rect 3732 15190 3800 15246
rect 3856 15190 3924 15246
rect 3980 15190 4048 15246
rect 4104 15190 4172 15246
rect 4228 15190 4296 15246
rect 4352 15190 4420 15246
rect 4476 15190 4544 15246
rect 4600 15190 4668 15246
rect 4724 15190 4734 15246
rect 2798 15122 4734 15190
rect 2798 15066 2808 15122
rect 2864 15066 2932 15122
rect 2988 15066 3056 15122
rect 3112 15066 3180 15122
rect 3236 15066 3304 15122
rect 3360 15066 3428 15122
rect 3484 15066 3552 15122
rect 3608 15066 3676 15122
rect 3732 15066 3800 15122
rect 3856 15066 3924 15122
rect 3980 15066 4048 15122
rect 4104 15066 4172 15122
rect 4228 15066 4296 15122
rect 4352 15066 4420 15122
rect 4476 15066 4544 15122
rect 4600 15066 4668 15122
rect 4724 15066 4734 15122
rect 2798 14998 4734 15066
rect 2798 14942 2808 14998
rect 2864 14942 2932 14998
rect 2988 14942 3056 14998
rect 3112 14942 3180 14998
rect 3236 14942 3304 14998
rect 3360 14942 3428 14998
rect 3484 14942 3552 14998
rect 3608 14942 3676 14998
rect 3732 14942 3800 14998
rect 3856 14942 3924 14998
rect 3980 14942 4048 14998
rect 4104 14942 4172 14998
rect 4228 14942 4296 14998
rect 4352 14942 4420 14998
rect 4476 14942 4544 14998
rect 4600 14942 4668 14998
rect 4724 14942 4734 14998
rect 2798 14874 4734 14942
rect 2798 14818 2808 14874
rect 2864 14818 2932 14874
rect 2988 14818 3056 14874
rect 3112 14818 3180 14874
rect 3236 14818 3304 14874
rect 3360 14818 3428 14874
rect 3484 14818 3552 14874
rect 3608 14818 3676 14874
rect 3732 14818 3800 14874
rect 3856 14818 3924 14874
rect 3980 14818 4048 14874
rect 4104 14818 4172 14874
rect 4228 14818 4296 14874
rect 4352 14818 4420 14874
rect 4476 14818 4544 14874
rect 4600 14818 4668 14874
rect 4724 14818 4734 14874
rect 2798 14750 4734 14818
rect 2798 14694 2808 14750
rect 2864 14694 2932 14750
rect 2988 14694 3056 14750
rect 3112 14694 3180 14750
rect 3236 14694 3304 14750
rect 3360 14694 3428 14750
rect 3484 14694 3552 14750
rect 3608 14694 3676 14750
rect 3732 14694 3800 14750
rect 3856 14694 3924 14750
rect 3980 14694 4048 14750
rect 4104 14694 4172 14750
rect 4228 14694 4296 14750
rect 4352 14694 4420 14750
rect 4476 14694 4544 14750
rect 4600 14694 4668 14750
rect 4724 14694 4734 14750
rect 2798 14626 4734 14694
rect 2798 14570 2808 14626
rect 2864 14570 2932 14626
rect 2988 14570 3056 14626
rect 3112 14570 3180 14626
rect 3236 14570 3304 14626
rect 3360 14570 3428 14626
rect 3484 14570 3552 14626
rect 3608 14570 3676 14626
rect 3732 14570 3800 14626
rect 3856 14570 3924 14626
rect 3980 14570 4048 14626
rect 4104 14570 4172 14626
rect 4228 14570 4296 14626
rect 4352 14570 4420 14626
rect 4476 14570 4544 14626
rect 4600 14570 4668 14626
rect 4724 14570 4734 14626
rect 2798 14502 4734 14570
rect 2798 14446 2808 14502
rect 2864 14446 2932 14502
rect 2988 14446 3056 14502
rect 3112 14446 3180 14502
rect 3236 14446 3304 14502
rect 3360 14446 3428 14502
rect 3484 14446 3552 14502
rect 3608 14446 3676 14502
rect 3732 14446 3800 14502
rect 3856 14446 3924 14502
rect 3980 14446 4048 14502
rect 4104 14446 4172 14502
rect 4228 14446 4296 14502
rect 4352 14446 4420 14502
rect 4476 14446 4544 14502
rect 4600 14446 4668 14502
rect 4724 14446 4734 14502
rect 2798 14436 4734 14446
rect 5168 17354 7104 17364
rect 5168 17298 5178 17354
rect 5234 17298 5302 17354
rect 5358 17298 5426 17354
rect 5482 17298 5550 17354
rect 5606 17298 5674 17354
rect 5730 17298 5798 17354
rect 5854 17298 5922 17354
rect 5978 17298 6046 17354
rect 6102 17298 6170 17354
rect 6226 17298 6294 17354
rect 6350 17298 6418 17354
rect 6474 17298 6542 17354
rect 6598 17298 6666 17354
rect 6722 17298 6790 17354
rect 6846 17298 6914 17354
rect 6970 17298 7038 17354
rect 7094 17298 7104 17354
rect 5168 17230 7104 17298
rect 5168 17174 5178 17230
rect 5234 17174 5302 17230
rect 5358 17174 5426 17230
rect 5482 17174 5550 17230
rect 5606 17174 5674 17230
rect 5730 17174 5798 17230
rect 5854 17174 5922 17230
rect 5978 17174 6046 17230
rect 6102 17174 6170 17230
rect 6226 17174 6294 17230
rect 6350 17174 6418 17230
rect 6474 17174 6542 17230
rect 6598 17174 6666 17230
rect 6722 17174 6790 17230
rect 6846 17174 6914 17230
rect 6970 17174 7038 17230
rect 7094 17174 7104 17230
rect 5168 17106 7104 17174
rect 5168 17050 5178 17106
rect 5234 17050 5302 17106
rect 5358 17050 5426 17106
rect 5482 17050 5550 17106
rect 5606 17050 5674 17106
rect 5730 17050 5798 17106
rect 5854 17050 5922 17106
rect 5978 17050 6046 17106
rect 6102 17050 6170 17106
rect 6226 17050 6294 17106
rect 6350 17050 6418 17106
rect 6474 17050 6542 17106
rect 6598 17050 6666 17106
rect 6722 17050 6790 17106
rect 6846 17050 6914 17106
rect 6970 17050 7038 17106
rect 7094 17050 7104 17106
rect 5168 16982 7104 17050
rect 5168 16926 5178 16982
rect 5234 16926 5302 16982
rect 5358 16926 5426 16982
rect 5482 16926 5550 16982
rect 5606 16926 5674 16982
rect 5730 16926 5798 16982
rect 5854 16926 5922 16982
rect 5978 16926 6046 16982
rect 6102 16926 6170 16982
rect 6226 16926 6294 16982
rect 6350 16926 6418 16982
rect 6474 16926 6542 16982
rect 6598 16926 6666 16982
rect 6722 16926 6790 16982
rect 6846 16926 6914 16982
rect 6970 16926 7038 16982
rect 7094 16926 7104 16982
rect 5168 16858 7104 16926
rect 5168 16802 5178 16858
rect 5234 16802 5302 16858
rect 5358 16802 5426 16858
rect 5482 16802 5550 16858
rect 5606 16802 5674 16858
rect 5730 16802 5798 16858
rect 5854 16802 5922 16858
rect 5978 16802 6046 16858
rect 6102 16802 6170 16858
rect 6226 16802 6294 16858
rect 6350 16802 6418 16858
rect 6474 16802 6542 16858
rect 6598 16802 6666 16858
rect 6722 16802 6790 16858
rect 6846 16802 6914 16858
rect 6970 16802 7038 16858
rect 7094 16802 7104 16858
rect 5168 16734 7104 16802
rect 5168 16678 5178 16734
rect 5234 16678 5302 16734
rect 5358 16678 5426 16734
rect 5482 16678 5550 16734
rect 5606 16678 5674 16734
rect 5730 16678 5798 16734
rect 5854 16678 5922 16734
rect 5978 16678 6046 16734
rect 6102 16678 6170 16734
rect 6226 16678 6294 16734
rect 6350 16678 6418 16734
rect 6474 16678 6542 16734
rect 6598 16678 6666 16734
rect 6722 16678 6790 16734
rect 6846 16678 6914 16734
rect 6970 16678 7038 16734
rect 7094 16678 7104 16734
rect 5168 16610 7104 16678
rect 5168 16554 5178 16610
rect 5234 16554 5302 16610
rect 5358 16554 5426 16610
rect 5482 16554 5550 16610
rect 5606 16554 5674 16610
rect 5730 16554 5798 16610
rect 5854 16554 5922 16610
rect 5978 16554 6046 16610
rect 6102 16554 6170 16610
rect 6226 16554 6294 16610
rect 6350 16554 6418 16610
rect 6474 16554 6542 16610
rect 6598 16554 6666 16610
rect 6722 16554 6790 16610
rect 6846 16554 6914 16610
rect 6970 16554 7038 16610
rect 7094 16554 7104 16610
rect 5168 16486 7104 16554
rect 5168 16430 5178 16486
rect 5234 16430 5302 16486
rect 5358 16430 5426 16486
rect 5482 16430 5550 16486
rect 5606 16430 5674 16486
rect 5730 16430 5798 16486
rect 5854 16430 5922 16486
rect 5978 16430 6046 16486
rect 6102 16430 6170 16486
rect 6226 16430 6294 16486
rect 6350 16430 6418 16486
rect 6474 16430 6542 16486
rect 6598 16430 6666 16486
rect 6722 16430 6790 16486
rect 6846 16430 6914 16486
rect 6970 16430 7038 16486
rect 7094 16430 7104 16486
rect 5168 16362 7104 16430
rect 5168 16306 5178 16362
rect 5234 16306 5302 16362
rect 5358 16306 5426 16362
rect 5482 16306 5550 16362
rect 5606 16306 5674 16362
rect 5730 16306 5798 16362
rect 5854 16306 5922 16362
rect 5978 16306 6046 16362
rect 6102 16306 6170 16362
rect 6226 16306 6294 16362
rect 6350 16306 6418 16362
rect 6474 16306 6542 16362
rect 6598 16306 6666 16362
rect 6722 16306 6790 16362
rect 6846 16306 6914 16362
rect 6970 16306 7038 16362
rect 7094 16306 7104 16362
rect 5168 16238 7104 16306
rect 5168 16182 5178 16238
rect 5234 16182 5302 16238
rect 5358 16182 5426 16238
rect 5482 16182 5550 16238
rect 5606 16182 5674 16238
rect 5730 16182 5798 16238
rect 5854 16182 5922 16238
rect 5978 16182 6046 16238
rect 6102 16182 6170 16238
rect 6226 16182 6294 16238
rect 6350 16182 6418 16238
rect 6474 16182 6542 16238
rect 6598 16182 6666 16238
rect 6722 16182 6790 16238
rect 6846 16182 6914 16238
rect 6970 16182 7038 16238
rect 7094 16182 7104 16238
rect 5168 16114 7104 16182
rect 5168 16058 5178 16114
rect 5234 16058 5302 16114
rect 5358 16058 5426 16114
rect 5482 16058 5550 16114
rect 5606 16058 5674 16114
rect 5730 16058 5798 16114
rect 5854 16058 5922 16114
rect 5978 16058 6046 16114
rect 6102 16058 6170 16114
rect 6226 16058 6294 16114
rect 6350 16058 6418 16114
rect 6474 16058 6542 16114
rect 6598 16058 6666 16114
rect 6722 16058 6790 16114
rect 6846 16058 6914 16114
rect 6970 16058 7038 16114
rect 7094 16058 7104 16114
rect 5168 15990 7104 16058
rect 5168 15934 5178 15990
rect 5234 15934 5302 15990
rect 5358 15934 5426 15990
rect 5482 15934 5550 15990
rect 5606 15934 5674 15990
rect 5730 15934 5798 15990
rect 5854 15934 5922 15990
rect 5978 15934 6046 15990
rect 6102 15934 6170 15990
rect 6226 15934 6294 15990
rect 6350 15934 6418 15990
rect 6474 15934 6542 15990
rect 6598 15934 6666 15990
rect 6722 15934 6790 15990
rect 6846 15934 6914 15990
rect 6970 15934 7038 15990
rect 7094 15934 7104 15990
rect 5168 15866 7104 15934
rect 5168 15810 5178 15866
rect 5234 15810 5302 15866
rect 5358 15810 5426 15866
rect 5482 15810 5550 15866
rect 5606 15810 5674 15866
rect 5730 15810 5798 15866
rect 5854 15810 5922 15866
rect 5978 15810 6046 15866
rect 6102 15810 6170 15866
rect 6226 15810 6294 15866
rect 6350 15810 6418 15866
rect 6474 15810 6542 15866
rect 6598 15810 6666 15866
rect 6722 15810 6790 15866
rect 6846 15810 6914 15866
rect 6970 15810 7038 15866
rect 7094 15810 7104 15866
rect 5168 15742 7104 15810
rect 5168 15686 5178 15742
rect 5234 15686 5302 15742
rect 5358 15686 5426 15742
rect 5482 15686 5550 15742
rect 5606 15686 5674 15742
rect 5730 15686 5798 15742
rect 5854 15686 5922 15742
rect 5978 15686 6046 15742
rect 6102 15686 6170 15742
rect 6226 15686 6294 15742
rect 6350 15686 6418 15742
rect 6474 15686 6542 15742
rect 6598 15686 6666 15742
rect 6722 15686 6790 15742
rect 6846 15686 6914 15742
rect 6970 15686 7038 15742
rect 7094 15686 7104 15742
rect 5168 15618 7104 15686
rect 5168 15562 5178 15618
rect 5234 15562 5302 15618
rect 5358 15562 5426 15618
rect 5482 15562 5550 15618
rect 5606 15562 5674 15618
rect 5730 15562 5798 15618
rect 5854 15562 5922 15618
rect 5978 15562 6046 15618
rect 6102 15562 6170 15618
rect 6226 15562 6294 15618
rect 6350 15562 6418 15618
rect 6474 15562 6542 15618
rect 6598 15562 6666 15618
rect 6722 15562 6790 15618
rect 6846 15562 6914 15618
rect 6970 15562 7038 15618
rect 7094 15562 7104 15618
rect 5168 15494 7104 15562
rect 5168 15438 5178 15494
rect 5234 15438 5302 15494
rect 5358 15438 5426 15494
rect 5482 15438 5550 15494
rect 5606 15438 5674 15494
rect 5730 15438 5798 15494
rect 5854 15438 5922 15494
rect 5978 15438 6046 15494
rect 6102 15438 6170 15494
rect 6226 15438 6294 15494
rect 6350 15438 6418 15494
rect 6474 15438 6542 15494
rect 6598 15438 6666 15494
rect 6722 15438 6790 15494
rect 6846 15438 6914 15494
rect 6970 15438 7038 15494
rect 7094 15438 7104 15494
rect 5168 15370 7104 15438
rect 5168 15314 5178 15370
rect 5234 15314 5302 15370
rect 5358 15314 5426 15370
rect 5482 15314 5550 15370
rect 5606 15314 5674 15370
rect 5730 15314 5798 15370
rect 5854 15314 5922 15370
rect 5978 15314 6046 15370
rect 6102 15314 6170 15370
rect 6226 15314 6294 15370
rect 6350 15314 6418 15370
rect 6474 15314 6542 15370
rect 6598 15314 6666 15370
rect 6722 15314 6790 15370
rect 6846 15314 6914 15370
rect 6970 15314 7038 15370
rect 7094 15314 7104 15370
rect 5168 15246 7104 15314
rect 5168 15190 5178 15246
rect 5234 15190 5302 15246
rect 5358 15190 5426 15246
rect 5482 15190 5550 15246
rect 5606 15190 5674 15246
rect 5730 15190 5798 15246
rect 5854 15190 5922 15246
rect 5978 15190 6046 15246
rect 6102 15190 6170 15246
rect 6226 15190 6294 15246
rect 6350 15190 6418 15246
rect 6474 15190 6542 15246
rect 6598 15190 6666 15246
rect 6722 15190 6790 15246
rect 6846 15190 6914 15246
rect 6970 15190 7038 15246
rect 7094 15190 7104 15246
rect 5168 15122 7104 15190
rect 5168 15066 5178 15122
rect 5234 15066 5302 15122
rect 5358 15066 5426 15122
rect 5482 15066 5550 15122
rect 5606 15066 5674 15122
rect 5730 15066 5798 15122
rect 5854 15066 5922 15122
rect 5978 15066 6046 15122
rect 6102 15066 6170 15122
rect 6226 15066 6294 15122
rect 6350 15066 6418 15122
rect 6474 15066 6542 15122
rect 6598 15066 6666 15122
rect 6722 15066 6790 15122
rect 6846 15066 6914 15122
rect 6970 15066 7038 15122
rect 7094 15066 7104 15122
rect 5168 14998 7104 15066
rect 5168 14942 5178 14998
rect 5234 14942 5302 14998
rect 5358 14942 5426 14998
rect 5482 14942 5550 14998
rect 5606 14942 5674 14998
rect 5730 14942 5798 14998
rect 5854 14942 5922 14998
rect 5978 14942 6046 14998
rect 6102 14942 6170 14998
rect 6226 14942 6294 14998
rect 6350 14942 6418 14998
rect 6474 14942 6542 14998
rect 6598 14942 6666 14998
rect 6722 14942 6790 14998
rect 6846 14942 6914 14998
rect 6970 14942 7038 14998
rect 7094 14942 7104 14998
rect 5168 14874 7104 14942
rect 5168 14818 5178 14874
rect 5234 14818 5302 14874
rect 5358 14818 5426 14874
rect 5482 14818 5550 14874
rect 5606 14818 5674 14874
rect 5730 14818 5798 14874
rect 5854 14818 5922 14874
rect 5978 14818 6046 14874
rect 6102 14818 6170 14874
rect 6226 14818 6294 14874
rect 6350 14818 6418 14874
rect 6474 14818 6542 14874
rect 6598 14818 6666 14874
rect 6722 14818 6790 14874
rect 6846 14818 6914 14874
rect 6970 14818 7038 14874
rect 7094 14818 7104 14874
rect 5168 14750 7104 14818
rect 5168 14694 5178 14750
rect 5234 14694 5302 14750
rect 5358 14694 5426 14750
rect 5482 14694 5550 14750
rect 5606 14694 5674 14750
rect 5730 14694 5798 14750
rect 5854 14694 5922 14750
rect 5978 14694 6046 14750
rect 6102 14694 6170 14750
rect 6226 14694 6294 14750
rect 6350 14694 6418 14750
rect 6474 14694 6542 14750
rect 6598 14694 6666 14750
rect 6722 14694 6790 14750
rect 6846 14694 6914 14750
rect 6970 14694 7038 14750
rect 7094 14694 7104 14750
rect 5168 14626 7104 14694
rect 5168 14570 5178 14626
rect 5234 14570 5302 14626
rect 5358 14570 5426 14626
rect 5482 14570 5550 14626
rect 5606 14570 5674 14626
rect 5730 14570 5798 14626
rect 5854 14570 5922 14626
rect 5978 14570 6046 14626
rect 6102 14570 6170 14626
rect 6226 14570 6294 14626
rect 6350 14570 6418 14626
rect 6474 14570 6542 14626
rect 6598 14570 6666 14626
rect 6722 14570 6790 14626
rect 6846 14570 6914 14626
rect 6970 14570 7038 14626
rect 7094 14570 7104 14626
rect 5168 14502 7104 14570
rect 5168 14446 5178 14502
rect 5234 14446 5302 14502
rect 5358 14446 5426 14502
rect 5482 14446 5550 14502
rect 5606 14446 5674 14502
rect 5730 14446 5798 14502
rect 5854 14446 5922 14502
rect 5978 14446 6046 14502
rect 6102 14446 6170 14502
rect 6226 14446 6294 14502
rect 6350 14446 6418 14502
rect 6474 14446 6542 14502
rect 6598 14446 6666 14502
rect 6722 14446 6790 14502
rect 6846 14446 6914 14502
rect 6970 14446 7038 14502
rect 7094 14446 7104 14502
rect 5168 14436 7104 14446
rect 7874 17354 9810 17364
rect 7874 17298 7884 17354
rect 7940 17298 8008 17354
rect 8064 17298 8132 17354
rect 8188 17298 8256 17354
rect 8312 17298 8380 17354
rect 8436 17298 8504 17354
rect 8560 17298 8628 17354
rect 8684 17298 8752 17354
rect 8808 17298 8876 17354
rect 8932 17298 9000 17354
rect 9056 17298 9124 17354
rect 9180 17298 9248 17354
rect 9304 17298 9372 17354
rect 9428 17298 9496 17354
rect 9552 17298 9620 17354
rect 9676 17298 9744 17354
rect 9800 17298 9810 17354
rect 7874 17230 9810 17298
rect 7874 17174 7884 17230
rect 7940 17174 8008 17230
rect 8064 17174 8132 17230
rect 8188 17174 8256 17230
rect 8312 17174 8380 17230
rect 8436 17174 8504 17230
rect 8560 17174 8628 17230
rect 8684 17174 8752 17230
rect 8808 17174 8876 17230
rect 8932 17174 9000 17230
rect 9056 17174 9124 17230
rect 9180 17174 9248 17230
rect 9304 17174 9372 17230
rect 9428 17174 9496 17230
rect 9552 17174 9620 17230
rect 9676 17174 9744 17230
rect 9800 17174 9810 17230
rect 7874 17106 9810 17174
rect 7874 17050 7884 17106
rect 7940 17050 8008 17106
rect 8064 17050 8132 17106
rect 8188 17050 8256 17106
rect 8312 17050 8380 17106
rect 8436 17050 8504 17106
rect 8560 17050 8628 17106
rect 8684 17050 8752 17106
rect 8808 17050 8876 17106
rect 8932 17050 9000 17106
rect 9056 17050 9124 17106
rect 9180 17050 9248 17106
rect 9304 17050 9372 17106
rect 9428 17050 9496 17106
rect 9552 17050 9620 17106
rect 9676 17050 9744 17106
rect 9800 17050 9810 17106
rect 7874 16982 9810 17050
rect 7874 16926 7884 16982
rect 7940 16926 8008 16982
rect 8064 16926 8132 16982
rect 8188 16926 8256 16982
rect 8312 16926 8380 16982
rect 8436 16926 8504 16982
rect 8560 16926 8628 16982
rect 8684 16926 8752 16982
rect 8808 16926 8876 16982
rect 8932 16926 9000 16982
rect 9056 16926 9124 16982
rect 9180 16926 9248 16982
rect 9304 16926 9372 16982
rect 9428 16926 9496 16982
rect 9552 16926 9620 16982
rect 9676 16926 9744 16982
rect 9800 16926 9810 16982
rect 7874 16858 9810 16926
rect 7874 16802 7884 16858
rect 7940 16802 8008 16858
rect 8064 16802 8132 16858
rect 8188 16802 8256 16858
rect 8312 16802 8380 16858
rect 8436 16802 8504 16858
rect 8560 16802 8628 16858
rect 8684 16802 8752 16858
rect 8808 16802 8876 16858
rect 8932 16802 9000 16858
rect 9056 16802 9124 16858
rect 9180 16802 9248 16858
rect 9304 16802 9372 16858
rect 9428 16802 9496 16858
rect 9552 16802 9620 16858
rect 9676 16802 9744 16858
rect 9800 16802 9810 16858
rect 7874 16734 9810 16802
rect 7874 16678 7884 16734
rect 7940 16678 8008 16734
rect 8064 16678 8132 16734
rect 8188 16678 8256 16734
rect 8312 16678 8380 16734
rect 8436 16678 8504 16734
rect 8560 16678 8628 16734
rect 8684 16678 8752 16734
rect 8808 16678 8876 16734
rect 8932 16678 9000 16734
rect 9056 16678 9124 16734
rect 9180 16678 9248 16734
rect 9304 16678 9372 16734
rect 9428 16678 9496 16734
rect 9552 16678 9620 16734
rect 9676 16678 9744 16734
rect 9800 16678 9810 16734
rect 7874 16610 9810 16678
rect 7874 16554 7884 16610
rect 7940 16554 8008 16610
rect 8064 16554 8132 16610
rect 8188 16554 8256 16610
rect 8312 16554 8380 16610
rect 8436 16554 8504 16610
rect 8560 16554 8628 16610
rect 8684 16554 8752 16610
rect 8808 16554 8876 16610
rect 8932 16554 9000 16610
rect 9056 16554 9124 16610
rect 9180 16554 9248 16610
rect 9304 16554 9372 16610
rect 9428 16554 9496 16610
rect 9552 16554 9620 16610
rect 9676 16554 9744 16610
rect 9800 16554 9810 16610
rect 7874 16486 9810 16554
rect 7874 16430 7884 16486
rect 7940 16430 8008 16486
rect 8064 16430 8132 16486
rect 8188 16430 8256 16486
rect 8312 16430 8380 16486
rect 8436 16430 8504 16486
rect 8560 16430 8628 16486
rect 8684 16430 8752 16486
rect 8808 16430 8876 16486
rect 8932 16430 9000 16486
rect 9056 16430 9124 16486
rect 9180 16430 9248 16486
rect 9304 16430 9372 16486
rect 9428 16430 9496 16486
rect 9552 16430 9620 16486
rect 9676 16430 9744 16486
rect 9800 16430 9810 16486
rect 7874 16362 9810 16430
rect 7874 16306 7884 16362
rect 7940 16306 8008 16362
rect 8064 16306 8132 16362
rect 8188 16306 8256 16362
rect 8312 16306 8380 16362
rect 8436 16306 8504 16362
rect 8560 16306 8628 16362
rect 8684 16306 8752 16362
rect 8808 16306 8876 16362
rect 8932 16306 9000 16362
rect 9056 16306 9124 16362
rect 9180 16306 9248 16362
rect 9304 16306 9372 16362
rect 9428 16306 9496 16362
rect 9552 16306 9620 16362
rect 9676 16306 9744 16362
rect 9800 16306 9810 16362
rect 7874 16238 9810 16306
rect 7874 16182 7884 16238
rect 7940 16182 8008 16238
rect 8064 16182 8132 16238
rect 8188 16182 8256 16238
rect 8312 16182 8380 16238
rect 8436 16182 8504 16238
rect 8560 16182 8628 16238
rect 8684 16182 8752 16238
rect 8808 16182 8876 16238
rect 8932 16182 9000 16238
rect 9056 16182 9124 16238
rect 9180 16182 9248 16238
rect 9304 16182 9372 16238
rect 9428 16182 9496 16238
rect 9552 16182 9620 16238
rect 9676 16182 9744 16238
rect 9800 16182 9810 16238
rect 7874 16114 9810 16182
rect 7874 16058 7884 16114
rect 7940 16058 8008 16114
rect 8064 16058 8132 16114
rect 8188 16058 8256 16114
rect 8312 16058 8380 16114
rect 8436 16058 8504 16114
rect 8560 16058 8628 16114
rect 8684 16058 8752 16114
rect 8808 16058 8876 16114
rect 8932 16058 9000 16114
rect 9056 16058 9124 16114
rect 9180 16058 9248 16114
rect 9304 16058 9372 16114
rect 9428 16058 9496 16114
rect 9552 16058 9620 16114
rect 9676 16058 9744 16114
rect 9800 16058 9810 16114
rect 7874 15990 9810 16058
rect 7874 15934 7884 15990
rect 7940 15934 8008 15990
rect 8064 15934 8132 15990
rect 8188 15934 8256 15990
rect 8312 15934 8380 15990
rect 8436 15934 8504 15990
rect 8560 15934 8628 15990
rect 8684 15934 8752 15990
rect 8808 15934 8876 15990
rect 8932 15934 9000 15990
rect 9056 15934 9124 15990
rect 9180 15934 9248 15990
rect 9304 15934 9372 15990
rect 9428 15934 9496 15990
rect 9552 15934 9620 15990
rect 9676 15934 9744 15990
rect 9800 15934 9810 15990
rect 7874 15866 9810 15934
rect 7874 15810 7884 15866
rect 7940 15810 8008 15866
rect 8064 15810 8132 15866
rect 8188 15810 8256 15866
rect 8312 15810 8380 15866
rect 8436 15810 8504 15866
rect 8560 15810 8628 15866
rect 8684 15810 8752 15866
rect 8808 15810 8876 15866
rect 8932 15810 9000 15866
rect 9056 15810 9124 15866
rect 9180 15810 9248 15866
rect 9304 15810 9372 15866
rect 9428 15810 9496 15866
rect 9552 15810 9620 15866
rect 9676 15810 9744 15866
rect 9800 15810 9810 15866
rect 7874 15742 9810 15810
rect 7874 15686 7884 15742
rect 7940 15686 8008 15742
rect 8064 15686 8132 15742
rect 8188 15686 8256 15742
rect 8312 15686 8380 15742
rect 8436 15686 8504 15742
rect 8560 15686 8628 15742
rect 8684 15686 8752 15742
rect 8808 15686 8876 15742
rect 8932 15686 9000 15742
rect 9056 15686 9124 15742
rect 9180 15686 9248 15742
rect 9304 15686 9372 15742
rect 9428 15686 9496 15742
rect 9552 15686 9620 15742
rect 9676 15686 9744 15742
rect 9800 15686 9810 15742
rect 7874 15618 9810 15686
rect 7874 15562 7884 15618
rect 7940 15562 8008 15618
rect 8064 15562 8132 15618
rect 8188 15562 8256 15618
rect 8312 15562 8380 15618
rect 8436 15562 8504 15618
rect 8560 15562 8628 15618
rect 8684 15562 8752 15618
rect 8808 15562 8876 15618
rect 8932 15562 9000 15618
rect 9056 15562 9124 15618
rect 9180 15562 9248 15618
rect 9304 15562 9372 15618
rect 9428 15562 9496 15618
rect 9552 15562 9620 15618
rect 9676 15562 9744 15618
rect 9800 15562 9810 15618
rect 7874 15494 9810 15562
rect 7874 15438 7884 15494
rect 7940 15438 8008 15494
rect 8064 15438 8132 15494
rect 8188 15438 8256 15494
rect 8312 15438 8380 15494
rect 8436 15438 8504 15494
rect 8560 15438 8628 15494
rect 8684 15438 8752 15494
rect 8808 15438 8876 15494
rect 8932 15438 9000 15494
rect 9056 15438 9124 15494
rect 9180 15438 9248 15494
rect 9304 15438 9372 15494
rect 9428 15438 9496 15494
rect 9552 15438 9620 15494
rect 9676 15438 9744 15494
rect 9800 15438 9810 15494
rect 7874 15370 9810 15438
rect 7874 15314 7884 15370
rect 7940 15314 8008 15370
rect 8064 15314 8132 15370
rect 8188 15314 8256 15370
rect 8312 15314 8380 15370
rect 8436 15314 8504 15370
rect 8560 15314 8628 15370
rect 8684 15314 8752 15370
rect 8808 15314 8876 15370
rect 8932 15314 9000 15370
rect 9056 15314 9124 15370
rect 9180 15314 9248 15370
rect 9304 15314 9372 15370
rect 9428 15314 9496 15370
rect 9552 15314 9620 15370
rect 9676 15314 9744 15370
rect 9800 15314 9810 15370
rect 7874 15246 9810 15314
rect 7874 15190 7884 15246
rect 7940 15190 8008 15246
rect 8064 15190 8132 15246
rect 8188 15190 8256 15246
rect 8312 15190 8380 15246
rect 8436 15190 8504 15246
rect 8560 15190 8628 15246
rect 8684 15190 8752 15246
rect 8808 15190 8876 15246
rect 8932 15190 9000 15246
rect 9056 15190 9124 15246
rect 9180 15190 9248 15246
rect 9304 15190 9372 15246
rect 9428 15190 9496 15246
rect 9552 15190 9620 15246
rect 9676 15190 9744 15246
rect 9800 15190 9810 15246
rect 7874 15122 9810 15190
rect 7874 15066 7884 15122
rect 7940 15066 8008 15122
rect 8064 15066 8132 15122
rect 8188 15066 8256 15122
rect 8312 15066 8380 15122
rect 8436 15066 8504 15122
rect 8560 15066 8628 15122
rect 8684 15066 8752 15122
rect 8808 15066 8876 15122
rect 8932 15066 9000 15122
rect 9056 15066 9124 15122
rect 9180 15066 9248 15122
rect 9304 15066 9372 15122
rect 9428 15066 9496 15122
rect 9552 15066 9620 15122
rect 9676 15066 9744 15122
rect 9800 15066 9810 15122
rect 7874 14998 9810 15066
rect 7874 14942 7884 14998
rect 7940 14942 8008 14998
rect 8064 14942 8132 14998
rect 8188 14942 8256 14998
rect 8312 14942 8380 14998
rect 8436 14942 8504 14998
rect 8560 14942 8628 14998
rect 8684 14942 8752 14998
rect 8808 14942 8876 14998
rect 8932 14942 9000 14998
rect 9056 14942 9124 14998
rect 9180 14942 9248 14998
rect 9304 14942 9372 14998
rect 9428 14942 9496 14998
rect 9552 14942 9620 14998
rect 9676 14942 9744 14998
rect 9800 14942 9810 14998
rect 7874 14874 9810 14942
rect 7874 14818 7884 14874
rect 7940 14818 8008 14874
rect 8064 14818 8132 14874
rect 8188 14818 8256 14874
rect 8312 14818 8380 14874
rect 8436 14818 8504 14874
rect 8560 14818 8628 14874
rect 8684 14818 8752 14874
rect 8808 14818 8876 14874
rect 8932 14818 9000 14874
rect 9056 14818 9124 14874
rect 9180 14818 9248 14874
rect 9304 14818 9372 14874
rect 9428 14818 9496 14874
rect 9552 14818 9620 14874
rect 9676 14818 9744 14874
rect 9800 14818 9810 14874
rect 7874 14750 9810 14818
rect 7874 14694 7884 14750
rect 7940 14694 8008 14750
rect 8064 14694 8132 14750
rect 8188 14694 8256 14750
rect 8312 14694 8380 14750
rect 8436 14694 8504 14750
rect 8560 14694 8628 14750
rect 8684 14694 8752 14750
rect 8808 14694 8876 14750
rect 8932 14694 9000 14750
rect 9056 14694 9124 14750
rect 9180 14694 9248 14750
rect 9304 14694 9372 14750
rect 9428 14694 9496 14750
rect 9552 14694 9620 14750
rect 9676 14694 9744 14750
rect 9800 14694 9810 14750
rect 7874 14626 9810 14694
rect 7874 14570 7884 14626
rect 7940 14570 8008 14626
rect 8064 14570 8132 14626
rect 8188 14570 8256 14626
rect 8312 14570 8380 14626
rect 8436 14570 8504 14626
rect 8560 14570 8628 14626
rect 8684 14570 8752 14626
rect 8808 14570 8876 14626
rect 8932 14570 9000 14626
rect 9056 14570 9124 14626
rect 9180 14570 9248 14626
rect 9304 14570 9372 14626
rect 9428 14570 9496 14626
rect 9552 14570 9620 14626
rect 9676 14570 9744 14626
rect 9800 14570 9810 14626
rect 7874 14502 9810 14570
rect 7874 14446 7884 14502
rect 7940 14446 8008 14502
rect 8064 14446 8132 14502
rect 8188 14446 8256 14502
rect 8312 14446 8380 14502
rect 8436 14446 8504 14502
rect 8560 14446 8628 14502
rect 8684 14446 8752 14502
rect 8808 14446 8876 14502
rect 8932 14446 9000 14502
rect 9056 14446 9124 14502
rect 9180 14446 9248 14502
rect 9304 14446 9372 14502
rect 9428 14446 9496 14502
rect 9552 14446 9620 14502
rect 9676 14446 9744 14502
rect 9800 14446 9810 14502
rect 7874 14436 9810 14446
rect 10244 17354 12180 17364
rect 10244 17298 10254 17354
rect 10310 17298 10378 17354
rect 10434 17298 10502 17354
rect 10558 17298 10626 17354
rect 10682 17298 10750 17354
rect 10806 17298 10874 17354
rect 10930 17298 10998 17354
rect 11054 17298 11122 17354
rect 11178 17298 11246 17354
rect 11302 17298 11370 17354
rect 11426 17298 11494 17354
rect 11550 17298 11618 17354
rect 11674 17298 11742 17354
rect 11798 17298 11866 17354
rect 11922 17298 11990 17354
rect 12046 17298 12114 17354
rect 12170 17298 12180 17354
rect 10244 17230 12180 17298
rect 10244 17174 10254 17230
rect 10310 17174 10378 17230
rect 10434 17174 10502 17230
rect 10558 17174 10626 17230
rect 10682 17174 10750 17230
rect 10806 17174 10874 17230
rect 10930 17174 10998 17230
rect 11054 17174 11122 17230
rect 11178 17174 11246 17230
rect 11302 17174 11370 17230
rect 11426 17174 11494 17230
rect 11550 17174 11618 17230
rect 11674 17174 11742 17230
rect 11798 17174 11866 17230
rect 11922 17174 11990 17230
rect 12046 17174 12114 17230
rect 12170 17174 12180 17230
rect 10244 17106 12180 17174
rect 10244 17050 10254 17106
rect 10310 17050 10378 17106
rect 10434 17050 10502 17106
rect 10558 17050 10626 17106
rect 10682 17050 10750 17106
rect 10806 17050 10874 17106
rect 10930 17050 10998 17106
rect 11054 17050 11122 17106
rect 11178 17050 11246 17106
rect 11302 17050 11370 17106
rect 11426 17050 11494 17106
rect 11550 17050 11618 17106
rect 11674 17050 11742 17106
rect 11798 17050 11866 17106
rect 11922 17050 11990 17106
rect 12046 17050 12114 17106
rect 12170 17050 12180 17106
rect 10244 16982 12180 17050
rect 10244 16926 10254 16982
rect 10310 16926 10378 16982
rect 10434 16926 10502 16982
rect 10558 16926 10626 16982
rect 10682 16926 10750 16982
rect 10806 16926 10874 16982
rect 10930 16926 10998 16982
rect 11054 16926 11122 16982
rect 11178 16926 11246 16982
rect 11302 16926 11370 16982
rect 11426 16926 11494 16982
rect 11550 16926 11618 16982
rect 11674 16926 11742 16982
rect 11798 16926 11866 16982
rect 11922 16926 11990 16982
rect 12046 16926 12114 16982
rect 12170 16926 12180 16982
rect 10244 16858 12180 16926
rect 10244 16802 10254 16858
rect 10310 16802 10378 16858
rect 10434 16802 10502 16858
rect 10558 16802 10626 16858
rect 10682 16802 10750 16858
rect 10806 16802 10874 16858
rect 10930 16802 10998 16858
rect 11054 16802 11122 16858
rect 11178 16802 11246 16858
rect 11302 16802 11370 16858
rect 11426 16802 11494 16858
rect 11550 16802 11618 16858
rect 11674 16802 11742 16858
rect 11798 16802 11866 16858
rect 11922 16802 11990 16858
rect 12046 16802 12114 16858
rect 12170 16802 12180 16858
rect 10244 16734 12180 16802
rect 10244 16678 10254 16734
rect 10310 16678 10378 16734
rect 10434 16678 10502 16734
rect 10558 16678 10626 16734
rect 10682 16678 10750 16734
rect 10806 16678 10874 16734
rect 10930 16678 10998 16734
rect 11054 16678 11122 16734
rect 11178 16678 11246 16734
rect 11302 16678 11370 16734
rect 11426 16678 11494 16734
rect 11550 16678 11618 16734
rect 11674 16678 11742 16734
rect 11798 16678 11866 16734
rect 11922 16678 11990 16734
rect 12046 16678 12114 16734
rect 12170 16678 12180 16734
rect 10244 16610 12180 16678
rect 10244 16554 10254 16610
rect 10310 16554 10378 16610
rect 10434 16554 10502 16610
rect 10558 16554 10626 16610
rect 10682 16554 10750 16610
rect 10806 16554 10874 16610
rect 10930 16554 10998 16610
rect 11054 16554 11122 16610
rect 11178 16554 11246 16610
rect 11302 16554 11370 16610
rect 11426 16554 11494 16610
rect 11550 16554 11618 16610
rect 11674 16554 11742 16610
rect 11798 16554 11866 16610
rect 11922 16554 11990 16610
rect 12046 16554 12114 16610
rect 12170 16554 12180 16610
rect 10244 16486 12180 16554
rect 10244 16430 10254 16486
rect 10310 16430 10378 16486
rect 10434 16430 10502 16486
rect 10558 16430 10626 16486
rect 10682 16430 10750 16486
rect 10806 16430 10874 16486
rect 10930 16430 10998 16486
rect 11054 16430 11122 16486
rect 11178 16430 11246 16486
rect 11302 16430 11370 16486
rect 11426 16430 11494 16486
rect 11550 16430 11618 16486
rect 11674 16430 11742 16486
rect 11798 16430 11866 16486
rect 11922 16430 11990 16486
rect 12046 16430 12114 16486
rect 12170 16430 12180 16486
rect 10244 16362 12180 16430
rect 10244 16306 10254 16362
rect 10310 16306 10378 16362
rect 10434 16306 10502 16362
rect 10558 16306 10626 16362
rect 10682 16306 10750 16362
rect 10806 16306 10874 16362
rect 10930 16306 10998 16362
rect 11054 16306 11122 16362
rect 11178 16306 11246 16362
rect 11302 16306 11370 16362
rect 11426 16306 11494 16362
rect 11550 16306 11618 16362
rect 11674 16306 11742 16362
rect 11798 16306 11866 16362
rect 11922 16306 11990 16362
rect 12046 16306 12114 16362
rect 12170 16306 12180 16362
rect 10244 16238 12180 16306
rect 10244 16182 10254 16238
rect 10310 16182 10378 16238
rect 10434 16182 10502 16238
rect 10558 16182 10626 16238
rect 10682 16182 10750 16238
rect 10806 16182 10874 16238
rect 10930 16182 10998 16238
rect 11054 16182 11122 16238
rect 11178 16182 11246 16238
rect 11302 16182 11370 16238
rect 11426 16182 11494 16238
rect 11550 16182 11618 16238
rect 11674 16182 11742 16238
rect 11798 16182 11866 16238
rect 11922 16182 11990 16238
rect 12046 16182 12114 16238
rect 12170 16182 12180 16238
rect 10244 16114 12180 16182
rect 10244 16058 10254 16114
rect 10310 16058 10378 16114
rect 10434 16058 10502 16114
rect 10558 16058 10626 16114
rect 10682 16058 10750 16114
rect 10806 16058 10874 16114
rect 10930 16058 10998 16114
rect 11054 16058 11122 16114
rect 11178 16058 11246 16114
rect 11302 16058 11370 16114
rect 11426 16058 11494 16114
rect 11550 16058 11618 16114
rect 11674 16058 11742 16114
rect 11798 16058 11866 16114
rect 11922 16058 11990 16114
rect 12046 16058 12114 16114
rect 12170 16058 12180 16114
rect 10244 15990 12180 16058
rect 10244 15934 10254 15990
rect 10310 15934 10378 15990
rect 10434 15934 10502 15990
rect 10558 15934 10626 15990
rect 10682 15934 10750 15990
rect 10806 15934 10874 15990
rect 10930 15934 10998 15990
rect 11054 15934 11122 15990
rect 11178 15934 11246 15990
rect 11302 15934 11370 15990
rect 11426 15934 11494 15990
rect 11550 15934 11618 15990
rect 11674 15934 11742 15990
rect 11798 15934 11866 15990
rect 11922 15934 11990 15990
rect 12046 15934 12114 15990
rect 12170 15934 12180 15990
rect 10244 15866 12180 15934
rect 10244 15810 10254 15866
rect 10310 15810 10378 15866
rect 10434 15810 10502 15866
rect 10558 15810 10626 15866
rect 10682 15810 10750 15866
rect 10806 15810 10874 15866
rect 10930 15810 10998 15866
rect 11054 15810 11122 15866
rect 11178 15810 11246 15866
rect 11302 15810 11370 15866
rect 11426 15810 11494 15866
rect 11550 15810 11618 15866
rect 11674 15810 11742 15866
rect 11798 15810 11866 15866
rect 11922 15810 11990 15866
rect 12046 15810 12114 15866
rect 12170 15810 12180 15866
rect 10244 15742 12180 15810
rect 10244 15686 10254 15742
rect 10310 15686 10378 15742
rect 10434 15686 10502 15742
rect 10558 15686 10626 15742
rect 10682 15686 10750 15742
rect 10806 15686 10874 15742
rect 10930 15686 10998 15742
rect 11054 15686 11122 15742
rect 11178 15686 11246 15742
rect 11302 15686 11370 15742
rect 11426 15686 11494 15742
rect 11550 15686 11618 15742
rect 11674 15686 11742 15742
rect 11798 15686 11866 15742
rect 11922 15686 11990 15742
rect 12046 15686 12114 15742
rect 12170 15686 12180 15742
rect 10244 15618 12180 15686
rect 10244 15562 10254 15618
rect 10310 15562 10378 15618
rect 10434 15562 10502 15618
rect 10558 15562 10626 15618
rect 10682 15562 10750 15618
rect 10806 15562 10874 15618
rect 10930 15562 10998 15618
rect 11054 15562 11122 15618
rect 11178 15562 11246 15618
rect 11302 15562 11370 15618
rect 11426 15562 11494 15618
rect 11550 15562 11618 15618
rect 11674 15562 11742 15618
rect 11798 15562 11866 15618
rect 11922 15562 11990 15618
rect 12046 15562 12114 15618
rect 12170 15562 12180 15618
rect 10244 15494 12180 15562
rect 10244 15438 10254 15494
rect 10310 15438 10378 15494
rect 10434 15438 10502 15494
rect 10558 15438 10626 15494
rect 10682 15438 10750 15494
rect 10806 15438 10874 15494
rect 10930 15438 10998 15494
rect 11054 15438 11122 15494
rect 11178 15438 11246 15494
rect 11302 15438 11370 15494
rect 11426 15438 11494 15494
rect 11550 15438 11618 15494
rect 11674 15438 11742 15494
rect 11798 15438 11866 15494
rect 11922 15438 11990 15494
rect 12046 15438 12114 15494
rect 12170 15438 12180 15494
rect 10244 15370 12180 15438
rect 10244 15314 10254 15370
rect 10310 15314 10378 15370
rect 10434 15314 10502 15370
rect 10558 15314 10626 15370
rect 10682 15314 10750 15370
rect 10806 15314 10874 15370
rect 10930 15314 10998 15370
rect 11054 15314 11122 15370
rect 11178 15314 11246 15370
rect 11302 15314 11370 15370
rect 11426 15314 11494 15370
rect 11550 15314 11618 15370
rect 11674 15314 11742 15370
rect 11798 15314 11866 15370
rect 11922 15314 11990 15370
rect 12046 15314 12114 15370
rect 12170 15314 12180 15370
rect 10244 15246 12180 15314
rect 10244 15190 10254 15246
rect 10310 15190 10378 15246
rect 10434 15190 10502 15246
rect 10558 15190 10626 15246
rect 10682 15190 10750 15246
rect 10806 15190 10874 15246
rect 10930 15190 10998 15246
rect 11054 15190 11122 15246
rect 11178 15190 11246 15246
rect 11302 15190 11370 15246
rect 11426 15190 11494 15246
rect 11550 15190 11618 15246
rect 11674 15190 11742 15246
rect 11798 15190 11866 15246
rect 11922 15190 11990 15246
rect 12046 15190 12114 15246
rect 12170 15190 12180 15246
rect 10244 15122 12180 15190
rect 10244 15066 10254 15122
rect 10310 15066 10378 15122
rect 10434 15066 10502 15122
rect 10558 15066 10626 15122
rect 10682 15066 10750 15122
rect 10806 15066 10874 15122
rect 10930 15066 10998 15122
rect 11054 15066 11122 15122
rect 11178 15066 11246 15122
rect 11302 15066 11370 15122
rect 11426 15066 11494 15122
rect 11550 15066 11618 15122
rect 11674 15066 11742 15122
rect 11798 15066 11866 15122
rect 11922 15066 11990 15122
rect 12046 15066 12114 15122
rect 12170 15066 12180 15122
rect 10244 14998 12180 15066
rect 10244 14942 10254 14998
rect 10310 14942 10378 14998
rect 10434 14942 10502 14998
rect 10558 14942 10626 14998
rect 10682 14942 10750 14998
rect 10806 14942 10874 14998
rect 10930 14942 10998 14998
rect 11054 14942 11122 14998
rect 11178 14942 11246 14998
rect 11302 14942 11370 14998
rect 11426 14942 11494 14998
rect 11550 14942 11618 14998
rect 11674 14942 11742 14998
rect 11798 14942 11866 14998
rect 11922 14942 11990 14998
rect 12046 14942 12114 14998
rect 12170 14942 12180 14998
rect 10244 14874 12180 14942
rect 10244 14818 10254 14874
rect 10310 14818 10378 14874
rect 10434 14818 10502 14874
rect 10558 14818 10626 14874
rect 10682 14818 10750 14874
rect 10806 14818 10874 14874
rect 10930 14818 10998 14874
rect 11054 14818 11122 14874
rect 11178 14818 11246 14874
rect 11302 14818 11370 14874
rect 11426 14818 11494 14874
rect 11550 14818 11618 14874
rect 11674 14818 11742 14874
rect 11798 14818 11866 14874
rect 11922 14818 11990 14874
rect 12046 14818 12114 14874
rect 12170 14818 12180 14874
rect 10244 14750 12180 14818
rect 10244 14694 10254 14750
rect 10310 14694 10378 14750
rect 10434 14694 10502 14750
rect 10558 14694 10626 14750
rect 10682 14694 10750 14750
rect 10806 14694 10874 14750
rect 10930 14694 10998 14750
rect 11054 14694 11122 14750
rect 11178 14694 11246 14750
rect 11302 14694 11370 14750
rect 11426 14694 11494 14750
rect 11550 14694 11618 14750
rect 11674 14694 11742 14750
rect 11798 14694 11866 14750
rect 11922 14694 11990 14750
rect 12046 14694 12114 14750
rect 12170 14694 12180 14750
rect 10244 14626 12180 14694
rect 10244 14570 10254 14626
rect 10310 14570 10378 14626
rect 10434 14570 10502 14626
rect 10558 14570 10626 14626
rect 10682 14570 10750 14626
rect 10806 14570 10874 14626
rect 10930 14570 10998 14626
rect 11054 14570 11122 14626
rect 11178 14570 11246 14626
rect 11302 14570 11370 14626
rect 11426 14570 11494 14626
rect 11550 14570 11618 14626
rect 11674 14570 11742 14626
rect 11798 14570 11866 14626
rect 11922 14570 11990 14626
rect 12046 14570 12114 14626
rect 12170 14570 12180 14626
rect 10244 14502 12180 14570
rect 10244 14446 10254 14502
rect 10310 14446 10378 14502
rect 10434 14446 10502 14502
rect 10558 14446 10626 14502
rect 10682 14446 10750 14502
rect 10806 14446 10874 14502
rect 10930 14446 10998 14502
rect 11054 14446 11122 14502
rect 11178 14446 11246 14502
rect 11302 14446 11370 14502
rect 11426 14446 11494 14502
rect 11550 14446 11618 14502
rect 11674 14446 11742 14502
rect 11798 14446 11866 14502
rect 11922 14446 11990 14502
rect 12046 14446 12114 14502
rect 12170 14446 12180 14502
rect 10244 14436 12180 14446
rect 12861 17354 14673 17364
rect 12861 17298 12871 17354
rect 12927 17298 12995 17354
rect 13051 17298 13119 17354
rect 13175 17298 13243 17354
rect 13299 17298 13367 17354
rect 13423 17298 13491 17354
rect 13547 17298 13615 17354
rect 13671 17298 13739 17354
rect 13795 17298 13863 17354
rect 13919 17298 13987 17354
rect 14043 17298 14111 17354
rect 14167 17298 14235 17354
rect 14291 17298 14359 17354
rect 14415 17298 14483 17354
rect 14539 17298 14607 17354
rect 14663 17298 14673 17354
rect 12861 17230 14673 17298
rect 12861 17174 12871 17230
rect 12927 17174 12995 17230
rect 13051 17174 13119 17230
rect 13175 17174 13243 17230
rect 13299 17174 13367 17230
rect 13423 17174 13491 17230
rect 13547 17174 13615 17230
rect 13671 17174 13739 17230
rect 13795 17174 13863 17230
rect 13919 17174 13987 17230
rect 14043 17174 14111 17230
rect 14167 17174 14235 17230
rect 14291 17174 14359 17230
rect 14415 17174 14483 17230
rect 14539 17174 14607 17230
rect 14663 17174 14673 17230
rect 12861 17106 14673 17174
rect 12861 17050 12871 17106
rect 12927 17050 12995 17106
rect 13051 17050 13119 17106
rect 13175 17050 13243 17106
rect 13299 17050 13367 17106
rect 13423 17050 13491 17106
rect 13547 17050 13615 17106
rect 13671 17050 13739 17106
rect 13795 17050 13863 17106
rect 13919 17050 13987 17106
rect 14043 17050 14111 17106
rect 14167 17050 14235 17106
rect 14291 17050 14359 17106
rect 14415 17050 14483 17106
rect 14539 17050 14607 17106
rect 14663 17050 14673 17106
rect 12861 16982 14673 17050
rect 12861 16926 12871 16982
rect 12927 16926 12995 16982
rect 13051 16926 13119 16982
rect 13175 16926 13243 16982
rect 13299 16926 13367 16982
rect 13423 16926 13491 16982
rect 13547 16926 13615 16982
rect 13671 16926 13739 16982
rect 13795 16926 13863 16982
rect 13919 16926 13987 16982
rect 14043 16926 14111 16982
rect 14167 16926 14235 16982
rect 14291 16926 14359 16982
rect 14415 16926 14483 16982
rect 14539 16926 14607 16982
rect 14663 16926 14673 16982
rect 12861 16858 14673 16926
rect 12861 16802 12871 16858
rect 12927 16802 12995 16858
rect 13051 16802 13119 16858
rect 13175 16802 13243 16858
rect 13299 16802 13367 16858
rect 13423 16802 13491 16858
rect 13547 16802 13615 16858
rect 13671 16802 13739 16858
rect 13795 16802 13863 16858
rect 13919 16802 13987 16858
rect 14043 16802 14111 16858
rect 14167 16802 14235 16858
rect 14291 16802 14359 16858
rect 14415 16802 14483 16858
rect 14539 16802 14607 16858
rect 14663 16802 14673 16858
rect 12861 16734 14673 16802
rect 12861 16678 12871 16734
rect 12927 16678 12995 16734
rect 13051 16678 13119 16734
rect 13175 16678 13243 16734
rect 13299 16678 13367 16734
rect 13423 16678 13491 16734
rect 13547 16678 13615 16734
rect 13671 16678 13739 16734
rect 13795 16678 13863 16734
rect 13919 16678 13987 16734
rect 14043 16678 14111 16734
rect 14167 16678 14235 16734
rect 14291 16678 14359 16734
rect 14415 16678 14483 16734
rect 14539 16678 14607 16734
rect 14663 16678 14673 16734
rect 12861 16610 14673 16678
rect 12861 16554 12871 16610
rect 12927 16554 12995 16610
rect 13051 16554 13119 16610
rect 13175 16554 13243 16610
rect 13299 16554 13367 16610
rect 13423 16554 13491 16610
rect 13547 16554 13615 16610
rect 13671 16554 13739 16610
rect 13795 16554 13863 16610
rect 13919 16554 13987 16610
rect 14043 16554 14111 16610
rect 14167 16554 14235 16610
rect 14291 16554 14359 16610
rect 14415 16554 14483 16610
rect 14539 16554 14607 16610
rect 14663 16554 14673 16610
rect 12861 16486 14673 16554
rect 12861 16430 12871 16486
rect 12927 16430 12995 16486
rect 13051 16430 13119 16486
rect 13175 16430 13243 16486
rect 13299 16430 13367 16486
rect 13423 16430 13491 16486
rect 13547 16430 13615 16486
rect 13671 16430 13739 16486
rect 13795 16430 13863 16486
rect 13919 16430 13987 16486
rect 14043 16430 14111 16486
rect 14167 16430 14235 16486
rect 14291 16430 14359 16486
rect 14415 16430 14483 16486
rect 14539 16430 14607 16486
rect 14663 16430 14673 16486
rect 12861 16362 14673 16430
rect 12861 16306 12871 16362
rect 12927 16306 12995 16362
rect 13051 16306 13119 16362
rect 13175 16306 13243 16362
rect 13299 16306 13367 16362
rect 13423 16306 13491 16362
rect 13547 16306 13615 16362
rect 13671 16306 13739 16362
rect 13795 16306 13863 16362
rect 13919 16306 13987 16362
rect 14043 16306 14111 16362
rect 14167 16306 14235 16362
rect 14291 16306 14359 16362
rect 14415 16306 14483 16362
rect 14539 16306 14607 16362
rect 14663 16306 14673 16362
rect 12861 16238 14673 16306
rect 12861 16182 12871 16238
rect 12927 16182 12995 16238
rect 13051 16182 13119 16238
rect 13175 16182 13243 16238
rect 13299 16182 13367 16238
rect 13423 16182 13491 16238
rect 13547 16182 13615 16238
rect 13671 16182 13739 16238
rect 13795 16182 13863 16238
rect 13919 16182 13987 16238
rect 14043 16182 14111 16238
rect 14167 16182 14235 16238
rect 14291 16182 14359 16238
rect 14415 16182 14483 16238
rect 14539 16182 14607 16238
rect 14663 16182 14673 16238
rect 12861 16114 14673 16182
rect 12861 16058 12871 16114
rect 12927 16058 12995 16114
rect 13051 16058 13119 16114
rect 13175 16058 13243 16114
rect 13299 16058 13367 16114
rect 13423 16058 13491 16114
rect 13547 16058 13615 16114
rect 13671 16058 13739 16114
rect 13795 16058 13863 16114
rect 13919 16058 13987 16114
rect 14043 16058 14111 16114
rect 14167 16058 14235 16114
rect 14291 16058 14359 16114
rect 14415 16058 14483 16114
rect 14539 16058 14607 16114
rect 14663 16058 14673 16114
rect 12861 15990 14673 16058
rect 12861 15934 12871 15990
rect 12927 15934 12995 15990
rect 13051 15934 13119 15990
rect 13175 15934 13243 15990
rect 13299 15934 13367 15990
rect 13423 15934 13491 15990
rect 13547 15934 13615 15990
rect 13671 15934 13739 15990
rect 13795 15934 13863 15990
rect 13919 15934 13987 15990
rect 14043 15934 14111 15990
rect 14167 15934 14235 15990
rect 14291 15934 14359 15990
rect 14415 15934 14483 15990
rect 14539 15934 14607 15990
rect 14663 15934 14673 15990
rect 12861 15866 14673 15934
rect 12861 15810 12871 15866
rect 12927 15810 12995 15866
rect 13051 15810 13119 15866
rect 13175 15810 13243 15866
rect 13299 15810 13367 15866
rect 13423 15810 13491 15866
rect 13547 15810 13615 15866
rect 13671 15810 13739 15866
rect 13795 15810 13863 15866
rect 13919 15810 13987 15866
rect 14043 15810 14111 15866
rect 14167 15810 14235 15866
rect 14291 15810 14359 15866
rect 14415 15810 14483 15866
rect 14539 15810 14607 15866
rect 14663 15810 14673 15866
rect 12861 15742 14673 15810
rect 12861 15686 12871 15742
rect 12927 15686 12995 15742
rect 13051 15686 13119 15742
rect 13175 15686 13243 15742
rect 13299 15686 13367 15742
rect 13423 15686 13491 15742
rect 13547 15686 13615 15742
rect 13671 15686 13739 15742
rect 13795 15686 13863 15742
rect 13919 15686 13987 15742
rect 14043 15686 14111 15742
rect 14167 15686 14235 15742
rect 14291 15686 14359 15742
rect 14415 15686 14483 15742
rect 14539 15686 14607 15742
rect 14663 15686 14673 15742
rect 12861 15618 14673 15686
rect 12861 15562 12871 15618
rect 12927 15562 12995 15618
rect 13051 15562 13119 15618
rect 13175 15562 13243 15618
rect 13299 15562 13367 15618
rect 13423 15562 13491 15618
rect 13547 15562 13615 15618
rect 13671 15562 13739 15618
rect 13795 15562 13863 15618
rect 13919 15562 13987 15618
rect 14043 15562 14111 15618
rect 14167 15562 14235 15618
rect 14291 15562 14359 15618
rect 14415 15562 14483 15618
rect 14539 15562 14607 15618
rect 14663 15562 14673 15618
rect 12861 15494 14673 15562
rect 12861 15438 12871 15494
rect 12927 15438 12995 15494
rect 13051 15438 13119 15494
rect 13175 15438 13243 15494
rect 13299 15438 13367 15494
rect 13423 15438 13491 15494
rect 13547 15438 13615 15494
rect 13671 15438 13739 15494
rect 13795 15438 13863 15494
rect 13919 15438 13987 15494
rect 14043 15438 14111 15494
rect 14167 15438 14235 15494
rect 14291 15438 14359 15494
rect 14415 15438 14483 15494
rect 14539 15438 14607 15494
rect 14663 15438 14673 15494
rect 12861 15370 14673 15438
rect 12861 15314 12871 15370
rect 12927 15314 12995 15370
rect 13051 15314 13119 15370
rect 13175 15314 13243 15370
rect 13299 15314 13367 15370
rect 13423 15314 13491 15370
rect 13547 15314 13615 15370
rect 13671 15314 13739 15370
rect 13795 15314 13863 15370
rect 13919 15314 13987 15370
rect 14043 15314 14111 15370
rect 14167 15314 14235 15370
rect 14291 15314 14359 15370
rect 14415 15314 14483 15370
rect 14539 15314 14607 15370
rect 14663 15314 14673 15370
rect 12861 15246 14673 15314
rect 12861 15190 12871 15246
rect 12927 15190 12995 15246
rect 13051 15190 13119 15246
rect 13175 15190 13243 15246
rect 13299 15190 13367 15246
rect 13423 15190 13491 15246
rect 13547 15190 13615 15246
rect 13671 15190 13739 15246
rect 13795 15190 13863 15246
rect 13919 15190 13987 15246
rect 14043 15190 14111 15246
rect 14167 15190 14235 15246
rect 14291 15190 14359 15246
rect 14415 15190 14483 15246
rect 14539 15190 14607 15246
rect 14663 15190 14673 15246
rect 12861 15122 14673 15190
rect 12861 15066 12871 15122
rect 12927 15066 12995 15122
rect 13051 15066 13119 15122
rect 13175 15066 13243 15122
rect 13299 15066 13367 15122
rect 13423 15066 13491 15122
rect 13547 15066 13615 15122
rect 13671 15066 13739 15122
rect 13795 15066 13863 15122
rect 13919 15066 13987 15122
rect 14043 15066 14111 15122
rect 14167 15066 14235 15122
rect 14291 15066 14359 15122
rect 14415 15066 14483 15122
rect 14539 15066 14607 15122
rect 14663 15066 14673 15122
rect 12861 14998 14673 15066
rect 12861 14942 12871 14998
rect 12927 14942 12995 14998
rect 13051 14942 13119 14998
rect 13175 14942 13243 14998
rect 13299 14942 13367 14998
rect 13423 14942 13491 14998
rect 13547 14942 13615 14998
rect 13671 14942 13739 14998
rect 13795 14942 13863 14998
rect 13919 14942 13987 14998
rect 14043 14942 14111 14998
rect 14167 14942 14235 14998
rect 14291 14942 14359 14998
rect 14415 14942 14483 14998
rect 14539 14942 14607 14998
rect 14663 14942 14673 14998
rect 12861 14874 14673 14942
rect 12861 14818 12871 14874
rect 12927 14818 12995 14874
rect 13051 14818 13119 14874
rect 13175 14818 13243 14874
rect 13299 14818 13367 14874
rect 13423 14818 13491 14874
rect 13547 14818 13615 14874
rect 13671 14818 13739 14874
rect 13795 14818 13863 14874
rect 13919 14818 13987 14874
rect 14043 14818 14111 14874
rect 14167 14818 14235 14874
rect 14291 14818 14359 14874
rect 14415 14818 14483 14874
rect 14539 14818 14607 14874
rect 14663 14818 14673 14874
rect 12861 14750 14673 14818
rect 12861 14694 12871 14750
rect 12927 14694 12995 14750
rect 13051 14694 13119 14750
rect 13175 14694 13243 14750
rect 13299 14694 13367 14750
rect 13423 14694 13491 14750
rect 13547 14694 13615 14750
rect 13671 14694 13739 14750
rect 13795 14694 13863 14750
rect 13919 14694 13987 14750
rect 14043 14694 14111 14750
rect 14167 14694 14235 14750
rect 14291 14694 14359 14750
rect 14415 14694 14483 14750
rect 14539 14694 14607 14750
rect 14663 14694 14673 14750
rect 12861 14626 14673 14694
rect 12861 14570 12871 14626
rect 12927 14570 12995 14626
rect 13051 14570 13119 14626
rect 13175 14570 13243 14626
rect 13299 14570 13367 14626
rect 13423 14570 13491 14626
rect 13547 14570 13615 14626
rect 13671 14570 13739 14626
rect 13795 14570 13863 14626
rect 13919 14570 13987 14626
rect 14043 14570 14111 14626
rect 14167 14570 14235 14626
rect 14291 14570 14359 14626
rect 14415 14570 14483 14626
rect 14539 14570 14607 14626
rect 14663 14570 14673 14626
rect 12861 14502 14673 14570
rect 12861 14446 12871 14502
rect 12927 14446 12995 14502
rect 13051 14446 13119 14502
rect 13175 14446 13243 14502
rect 13299 14446 13367 14502
rect 13423 14446 13491 14502
rect 13547 14446 13615 14502
rect 13671 14446 13739 14502
rect 13795 14446 13863 14502
rect 13919 14446 13987 14502
rect 14043 14446 14111 14502
rect 14167 14446 14235 14502
rect 14291 14446 14359 14502
rect 14415 14446 14483 14502
rect 14539 14446 14607 14502
rect 14663 14446 14673 14502
rect 12861 14436 14673 14446
rect 2481 14148 2681 14158
rect 2481 14092 2491 14148
rect 2547 14092 2615 14148
rect 2671 14092 2681 14148
rect 2481 14024 2681 14092
rect 2481 13968 2491 14024
rect 2547 13968 2615 14024
rect 2671 13968 2681 14024
rect 2481 13900 2681 13968
rect 2481 13844 2491 13900
rect 2547 13844 2615 13900
rect 2671 13844 2681 13900
rect 2481 13776 2681 13844
rect 2481 13720 2491 13776
rect 2547 13720 2615 13776
rect 2671 13720 2681 13776
rect 2481 13652 2681 13720
rect 2481 13596 2491 13652
rect 2547 13596 2615 13652
rect 2671 13596 2681 13652
rect 2481 13528 2681 13596
rect 2481 13472 2491 13528
rect 2547 13472 2615 13528
rect 2671 13472 2681 13528
rect 2481 13404 2681 13472
rect 2481 13348 2491 13404
rect 2547 13348 2615 13404
rect 2671 13348 2681 13404
rect 2481 13280 2681 13348
rect 2481 13224 2491 13280
rect 2547 13224 2615 13280
rect 2671 13224 2681 13280
rect 2481 13156 2681 13224
rect 2481 13100 2491 13156
rect 2547 13100 2615 13156
rect 2671 13100 2681 13156
rect 2481 13032 2681 13100
rect 2481 12976 2491 13032
rect 2547 12976 2615 13032
rect 2671 12976 2681 13032
rect 2481 12908 2681 12976
rect 2481 12852 2491 12908
rect 2547 12852 2615 12908
rect 2671 12852 2681 12908
rect 2481 12842 2681 12852
rect 4851 14148 5051 14158
rect 4851 14092 4861 14148
rect 4917 14092 4985 14148
rect 5041 14092 5051 14148
rect 4851 14024 5051 14092
rect 4851 13968 4861 14024
rect 4917 13968 4985 14024
rect 5041 13968 5051 14024
rect 4851 13900 5051 13968
rect 4851 13844 4861 13900
rect 4917 13844 4985 13900
rect 5041 13844 5051 13900
rect 4851 13776 5051 13844
rect 4851 13720 4861 13776
rect 4917 13720 4985 13776
rect 5041 13720 5051 13776
rect 4851 13652 5051 13720
rect 4851 13596 4861 13652
rect 4917 13596 4985 13652
rect 5041 13596 5051 13652
rect 4851 13528 5051 13596
rect 4851 13472 4861 13528
rect 4917 13472 4985 13528
rect 5041 13472 5051 13528
rect 4851 13404 5051 13472
rect 4851 13348 4861 13404
rect 4917 13348 4985 13404
rect 5041 13348 5051 13404
rect 4851 13280 5051 13348
rect 4851 13224 4861 13280
rect 4917 13224 4985 13280
rect 5041 13224 5051 13280
rect 4851 13156 5051 13224
rect 4851 13100 4861 13156
rect 4917 13100 4985 13156
rect 5041 13100 5051 13156
rect 4851 13032 5051 13100
rect 4851 12976 4861 13032
rect 4917 12976 4985 13032
rect 5041 12976 5051 13032
rect 4851 12908 5051 12976
rect 4851 12852 4861 12908
rect 4917 12852 4985 12908
rect 5041 12852 5051 12908
rect 4851 12842 5051 12852
rect 7265 14148 7713 14158
rect 7265 14092 7275 14148
rect 7331 14092 7399 14148
rect 7455 14092 7523 14148
rect 7579 14092 7647 14148
rect 7703 14092 7713 14148
rect 7265 14024 7713 14092
rect 7265 13968 7275 14024
rect 7331 13968 7399 14024
rect 7455 13968 7523 14024
rect 7579 13968 7647 14024
rect 7703 13968 7713 14024
rect 7265 13900 7713 13968
rect 7265 13844 7275 13900
rect 7331 13844 7399 13900
rect 7455 13844 7523 13900
rect 7579 13844 7647 13900
rect 7703 13844 7713 13900
rect 7265 13776 7713 13844
rect 7265 13720 7275 13776
rect 7331 13720 7399 13776
rect 7455 13720 7523 13776
rect 7579 13720 7647 13776
rect 7703 13720 7713 13776
rect 7265 13652 7713 13720
rect 7265 13596 7275 13652
rect 7331 13596 7399 13652
rect 7455 13596 7523 13652
rect 7579 13596 7647 13652
rect 7703 13596 7713 13652
rect 7265 13528 7713 13596
rect 7265 13472 7275 13528
rect 7331 13472 7399 13528
rect 7455 13472 7523 13528
rect 7579 13472 7647 13528
rect 7703 13472 7713 13528
rect 7265 13404 7713 13472
rect 7265 13348 7275 13404
rect 7331 13348 7399 13404
rect 7455 13348 7523 13404
rect 7579 13348 7647 13404
rect 7703 13348 7713 13404
rect 7265 13280 7713 13348
rect 7265 13224 7275 13280
rect 7331 13224 7399 13280
rect 7455 13224 7523 13280
rect 7579 13224 7647 13280
rect 7703 13224 7713 13280
rect 7265 13156 7713 13224
rect 7265 13100 7275 13156
rect 7331 13100 7399 13156
rect 7455 13100 7523 13156
rect 7579 13100 7647 13156
rect 7703 13100 7713 13156
rect 7265 13032 7713 13100
rect 7265 12976 7275 13032
rect 7331 12976 7399 13032
rect 7455 12976 7523 13032
rect 7579 12976 7647 13032
rect 7703 12976 7713 13032
rect 7265 12908 7713 12976
rect 7265 12852 7275 12908
rect 7331 12852 7399 12908
rect 7455 12852 7523 12908
rect 7579 12852 7647 12908
rect 7703 12852 7713 12908
rect 7265 12842 7713 12852
rect 9927 14148 10127 14158
rect 9927 14092 9937 14148
rect 9993 14092 10061 14148
rect 10117 14092 10127 14148
rect 9927 14024 10127 14092
rect 9927 13968 9937 14024
rect 9993 13968 10061 14024
rect 10117 13968 10127 14024
rect 9927 13900 10127 13968
rect 9927 13844 9937 13900
rect 9993 13844 10061 13900
rect 10117 13844 10127 13900
rect 9927 13776 10127 13844
rect 9927 13720 9937 13776
rect 9993 13720 10061 13776
rect 10117 13720 10127 13776
rect 9927 13652 10127 13720
rect 9927 13596 9937 13652
rect 9993 13596 10061 13652
rect 10117 13596 10127 13652
rect 9927 13528 10127 13596
rect 9927 13472 9937 13528
rect 9993 13472 10061 13528
rect 10117 13472 10127 13528
rect 9927 13404 10127 13472
rect 9927 13348 9937 13404
rect 9993 13348 10061 13404
rect 10117 13348 10127 13404
rect 9927 13280 10127 13348
rect 9927 13224 9937 13280
rect 9993 13224 10061 13280
rect 10117 13224 10127 13280
rect 9927 13156 10127 13224
rect 9927 13100 9937 13156
rect 9993 13100 10061 13156
rect 10117 13100 10127 13156
rect 9927 13032 10127 13100
rect 9927 12976 9937 13032
rect 9993 12976 10061 13032
rect 10117 12976 10127 13032
rect 9927 12908 10127 12976
rect 9927 12852 9937 12908
rect 9993 12852 10061 12908
rect 10117 12852 10127 12908
rect 9927 12842 10127 12852
rect 12297 14148 12497 14158
rect 12297 14092 12307 14148
rect 12363 14092 12431 14148
rect 12487 14092 12497 14148
rect 12297 14024 12497 14092
rect 12297 13968 12307 14024
rect 12363 13968 12431 14024
rect 12487 13968 12497 14024
rect 12297 13900 12497 13968
rect 12297 13844 12307 13900
rect 12363 13844 12431 13900
rect 12487 13844 12497 13900
rect 12297 13776 12497 13844
rect 12297 13720 12307 13776
rect 12363 13720 12431 13776
rect 12487 13720 12497 13776
rect 12297 13652 12497 13720
rect 12297 13596 12307 13652
rect 12363 13596 12431 13652
rect 12487 13596 12497 13652
rect 12297 13528 12497 13596
rect 12297 13472 12307 13528
rect 12363 13472 12431 13528
rect 12487 13472 12497 13528
rect 12297 13404 12497 13472
rect 12297 13348 12307 13404
rect 12363 13348 12431 13404
rect 12487 13348 12497 13404
rect 12297 13280 12497 13348
rect 12297 13224 12307 13280
rect 12363 13224 12431 13280
rect 12487 13224 12497 13280
rect 12297 13156 12497 13224
rect 12297 13100 12307 13156
rect 12363 13100 12431 13156
rect 12487 13100 12497 13156
rect 12297 13032 12497 13100
rect 12297 12976 12307 13032
rect 12363 12976 12431 13032
rect 12487 12976 12497 13032
rect 12297 12908 12497 12976
rect 12297 12852 12307 12908
rect 12363 12852 12431 12908
rect 12487 12852 12497 12908
rect 12297 12842 12497 12852
rect 305 12548 2117 12558
rect 305 12492 315 12548
rect 371 12492 439 12548
rect 495 12492 563 12548
rect 619 12492 687 12548
rect 743 12492 811 12548
rect 867 12492 935 12548
rect 991 12492 1059 12548
rect 1115 12492 1183 12548
rect 1239 12492 1307 12548
rect 1363 12492 1431 12548
rect 1487 12492 1555 12548
rect 1611 12492 1679 12548
rect 1735 12492 1803 12548
rect 1859 12492 1927 12548
rect 1983 12492 2051 12548
rect 2107 12492 2117 12548
rect 305 12424 2117 12492
rect 305 12368 315 12424
rect 371 12368 439 12424
rect 495 12368 563 12424
rect 619 12368 687 12424
rect 743 12368 811 12424
rect 867 12368 935 12424
rect 991 12368 1059 12424
rect 1115 12368 1183 12424
rect 1239 12368 1307 12424
rect 1363 12368 1431 12424
rect 1487 12368 1555 12424
rect 1611 12368 1679 12424
rect 1735 12368 1803 12424
rect 1859 12368 1927 12424
rect 1983 12368 2051 12424
rect 2107 12368 2117 12424
rect 305 12300 2117 12368
rect 305 12244 315 12300
rect 371 12244 439 12300
rect 495 12244 563 12300
rect 619 12244 687 12300
rect 743 12244 811 12300
rect 867 12244 935 12300
rect 991 12244 1059 12300
rect 1115 12244 1183 12300
rect 1239 12244 1307 12300
rect 1363 12244 1431 12300
rect 1487 12244 1555 12300
rect 1611 12244 1679 12300
rect 1735 12244 1803 12300
rect 1859 12244 1927 12300
rect 1983 12244 2051 12300
rect 2107 12244 2117 12300
rect 305 12176 2117 12244
rect 305 12120 315 12176
rect 371 12120 439 12176
rect 495 12120 563 12176
rect 619 12120 687 12176
rect 743 12120 811 12176
rect 867 12120 935 12176
rect 991 12120 1059 12176
rect 1115 12120 1183 12176
rect 1239 12120 1307 12176
rect 1363 12120 1431 12176
rect 1487 12120 1555 12176
rect 1611 12120 1679 12176
rect 1735 12120 1803 12176
rect 1859 12120 1927 12176
rect 1983 12120 2051 12176
rect 2107 12120 2117 12176
rect 305 12052 2117 12120
rect 305 11996 315 12052
rect 371 11996 439 12052
rect 495 11996 563 12052
rect 619 11996 687 12052
rect 743 11996 811 12052
rect 867 11996 935 12052
rect 991 11996 1059 12052
rect 1115 11996 1183 12052
rect 1239 11996 1307 12052
rect 1363 11996 1431 12052
rect 1487 11996 1555 12052
rect 1611 11996 1679 12052
rect 1735 11996 1803 12052
rect 1859 11996 1927 12052
rect 1983 11996 2051 12052
rect 2107 11996 2117 12052
rect 305 11928 2117 11996
rect 305 11872 315 11928
rect 371 11872 439 11928
rect 495 11872 563 11928
rect 619 11872 687 11928
rect 743 11872 811 11928
rect 867 11872 935 11928
rect 991 11872 1059 11928
rect 1115 11872 1183 11928
rect 1239 11872 1307 11928
rect 1363 11872 1431 11928
rect 1487 11872 1555 11928
rect 1611 11872 1679 11928
rect 1735 11872 1803 11928
rect 1859 11872 1927 11928
rect 1983 11872 2051 11928
rect 2107 11872 2117 11928
rect 305 11804 2117 11872
rect 305 11748 315 11804
rect 371 11748 439 11804
rect 495 11748 563 11804
rect 619 11748 687 11804
rect 743 11748 811 11804
rect 867 11748 935 11804
rect 991 11748 1059 11804
rect 1115 11748 1183 11804
rect 1239 11748 1307 11804
rect 1363 11748 1431 11804
rect 1487 11748 1555 11804
rect 1611 11748 1679 11804
rect 1735 11748 1803 11804
rect 1859 11748 1927 11804
rect 1983 11748 2051 11804
rect 2107 11748 2117 11804
rect 305 11680 2117 11748
rect 305 11624 315 11680
rect 371 11624 439 11680
rect 495 11624 563 11680
rect 619 11624 687 11680
rect 743 11624 811 11680
rect 867 11624 935 11680
rect 991 11624 1059 11680
rect 1115 11624 1183 11680
rect 1239 11624 1307 11680
rect 1363 11624 1431 11680
rect 1487 11624 1555 11680
rect 1611 11624 1679 11680
rect 1735 11624 1803 11680
rect 1859 11624 1927 11680
rect 1983 11624 2051 11680
rect 2107 11624 2117 11680
rect 305 11556 2117 11624
rect 305 11500 315 11556
rect 371 11500 439 11556
rect 495 11500 563 11556
rect 619 11500 687 11556
rect 743 11500 811 11556
rect 867 11500 935 11556
rect 991 11500 1059 11556
rect 1115 11500 1183 11556
rect 1239 11500 1307 11556
rect 1363 11500 1431 11556
rect 1487 11500 1555 11556
rect 1611 11500 1679 11556
rect 1735 11500 1803 11556
rect 1859 11500 1927 11556
rect 1983 11500 2051 11556
rect 2107 11500 2117 11556
rect 305 11432 2117 11500
rect 305 11376 315 11432
rect 371 11376 439 11432
rect 495 11376 563 11432
rect 619 11376 687 11432
rect 743 11376 811 11432
rect 867 11376 935 11432
rect 991 11376 1059 11432
rect 1115 11376 1183 11432
rect 1239 11376 1307 11432
rect 1363 11376 1431 11432
rect 1487 11376 1555 11432
rect 1611 11376 1679 11432
rect 1735 11376 1803 11432
rect 1859 11376 1927 11432
rect 1983 11376 2051 11432
rect 2107 11376 2117 11432
rect 305 11308 2117 11376
rect 305 11252 315 11308
rect 371 11252 439 11308
rect 495 11252 563 11308
rect 619 11252 687 11308
rect 743 11252 811 11308
rect 867 11252 935 11308
rect 991 11252 1059 11308
rect 1115 11252 1183 11308
rect 1239 11252 1307 11308
rect 1363 11252 1431 11308
rect 1487 11252 1555 11308
rect 1611 11252 1679 11308
rect 1735 11252 1803 11308
rect 1859 11252 1927 11308
rect 1983 11252 2051 11308
rect 2107 11252 2117 11308
rect 305 11242 2117 11252
rect 2798 12548 4734 12558
rect 2798 12492 2808 12548
rect 2864 12492 2932 12548
rect 2988 12492 3056 12548
rect 3112 12492 3180 12548
rect 3236 12492 3304 12548
rect 3360 12492 3428 12548
rect 3484 12492 3552 12548
rect 3608 12492 3676 12548
rect 3732 12492 3800 12548
rect 3856 12492 3924 12548
rect 3980 12492 4048 12548
rect 4104 12492 4172 12548
rect 4228 12492 4296 12548
rect 4352 12492 4420 12548
rect 4476 12492 4544 12548
rect 4600 12492 4668 12548
rect 4724 12492 4734 12548
rect 2798 12424 4734 12492
rect 2798 12368 2808 12424
rect 2864 12368 2932 12424
rect 2988 12368 3056 12424
rect 3112 12368 3180 12424
rect 3236 12368 3304 12424
rect 3360 12368 3428 12424
rect 3484 12368 3552 12424
rect 3608 12368 3676 12424
rect 3732 12368 3800 12424
rect 3856 12368 3924 12424
rect 3980 12368 4048 12424
rect 4104 12368 4172 12424
rect 4228 12368 4296 12424
rect 4352 12368 4420 12424
rect 4476 12368 4544 12424
rect 4600 12368 4668 12424
rect 4724 12368 4734 12424
rect 2798 12300 4734 12368
rect 2798 12244 2808 12300
rect 2864 12244 2932 12300
rect 2988 12244 3056 12300
rect 3112 12244 3180 12300
rect 3236 12244 3304 12300
rect 3360 12244 3428 12300
rect 3484 12244 3552 12300
rect 3608 12244 3676 12300
rect 3732 12244 3800 12300
rect 3856 12244 3924 12300
rect 3980 12244 4048 12300
rect 4104 12244 4172 12300
rect 4228 12244 4296 12300
rect 4352 12244 4420 12300
rect 4476 12244 4544 12300
rect 4600 12244 4668 12300
rect 4724 12244 4734 12300
rect 2798 12176 4734 12244
rect 2798 12120 2808 12176
rect 2864 12120 2932 12176
rect 2988 12120 3056 12176
rect 3112 12120 3180 12176
rect 3236 12120 3304 12176
rect 3360 12120 3428 12176
rect 3484 12120 3552 12176
rect 3608 12120 3676 12176
rect 3732 12120 3800 12176
rect 3856 12120 3924 12176
rect 3980 12120 4048 12176
rect 4104 12120 4172 12176
rect 4228 12120 4296 12176
rect 4352 12120 4420 12176
rect 4476 12120 4544 12176
rect 4600 12120 4668 12176
rect 4724 12120 4734 12176
rect 2798 12052 4734 12120
rect 2798 11996 2808 12052
rect 2864 11996 2932 12052
rect 2988 11996 3056 12052
rect 3112 11996 3180 12052
rect 3236 11996 3304 12052
rect 3360 11996 3428 12052
rect 3484 11996 3552 12052
rect 3608 11996 3676 12052
rect 3732 11996 3800 12052
rect 3856 11996 3924 12052
rect 3980 11996 4048 12052
rect 4104 11996 4172 12052
rect 4228 11996 4296 12052
rect 4352 11996 4420 12052
rect 4476 11996 4544 12052
rect 4600 11996 4668 12052
rect 4724 11996 4734 12052
rect 2798 11928 4734 11996
rect 2798 11872 2808 11928
rect 2864 11872 2932 11928
rect 2988 11872 3056 11928
rect 3112 11872 3180 11928
rect 3236 11872 3304 11928
rect 3360 11872 3428 11928
rect 3484 11872 3552 11928
rect 3608 11872 3676 11928
rect 3732 11872 3800 11928
rect 3856 11872 3924 11928
rect 3980 11872 4048 11928
rect 4104 11872 4172 11928
rect 4228 11872 4296 11928
rect 4352 11872 4420 11928
rect 4476 11872 4544 11928
rect 4600 11872 4668 11928
rect 4724 11872 4734 11928
rect 2798 11804 4734 11872
rect 2798 11748 2808 11804
rect 2864 11748 2932 11804
rect 2988 11748 3056 11804
rect 3112 11748 3180 11804
rect 3236 11748 3304 11804
rect 3360 11748 3428 11804
rect 3484 11748 3552 11804
rect 3608 11748 3676 11804
rect 3732 11748 3800 11804
rect 3856 11748 3924 11804
rect 3980 11748 4048 11804
rect 4104 11748 4172 11804
rect 4228 11748 4296 11804
rect 4352 11748 4420 11804
rect 4476 11748 4544 11804
rect 4600 11748 4668 11804
rect 4724 11748 4734 11804
rect 2798 11680 4734 11748
rect 2798 11624 2808 11680
rect 2864 11624 2932 11680
rect 2988 11624 3056 11680
rect 3112 11624 3180 11680
rect 3236 11624 3304 11680
rect 3360 11624 3428 11680
rect 3484 11624 3552 11680
rect 3608 11624 3676 11680
rect 3732 11624 3800 11680
rect 3856 11624 3924 11680
rect 3980 11624 4048 11680
rect 4104 11624 4172 11680
rect 4228 11624 4296 11680
rect 4352 11624 4420 11680
rect 4476 11624 4544 11680
rect 4600 11624 4668 11680
rect 4724 11624 4734 11680
rect 2798 11556 4734 11624
rect 2798 11500 2808 11556
rect 2864 11500 2932 11556
rect 2988 11500 3056 11556
rect 3112 11500 3180 11556
rect 3236 11500 3304 11556
rect 3360 11500 3428 11556
rect 3484 11500 3552 11556
rect 3608 11500 3676 11556
rect 3732 11500 3800 11556
rect 3856 11500 3924 11556
rect 3980 11500 4048 11556
rect 4104 11500 4172 11556
rect 4228 11500 4296 11556
rect 4352 11500 4420 11556
rect 4476 11500 4544 11556
rect 4600 11500 4668 11556
rect 4724 11500 4734 11556
rect 2798 11432 4734 11500
rect 2798 11376 2808 11432
rect 2864 11376 2932 11432
rect 2988 11376 3056 11432
rect 3112 11376 3180 11432
rect 3236 11376 3304 11432
rect 3360 11376 3428 11432
rect 3484 11376 3552 11432
rect 3608 11376 3676 11432
rect 3732 11376 3800 11432
rect 3856 11376 3924 11432
rect 3980 11376 4048 11432
rect 4104 11376 4172 11432
rect 4228 11376 4296 11432
rect 4352 11376 4420 11432
rect 4476 11376 4544 11432
rect 4600 11376 4668 11432
rect 4724 11376 4734 11432
rect 2798 11308 4734 11376
rect 2798 11252 2808 11308
rect 2864 11252 2932 11308
rect 2988 11252 3056 11308
rect 3112 11252 3180 11308
rect 3236 11252 3304 11308
rect 3360 11252 3428 11308
rect 3484 11252 3552 11308
rect 3608 11252 3676 11308
rect 3732 11252 3800 11308
rect 3856 11252 3924 11308
rect 3980 11252 4048 11308
rect 4104 11252 4172 11308
rect 4228 11252 4296 11308
rect 4352 11252 4420 11308
rect 4476 11252 4544 11308
rect 4600 11252 4668 11308
rect 4724 11252 4734 11308
rect 2798 11242 4734 11252
rect 5168 12548 7104 12558
rect 5168 12492 5178 12548
rect 5234 12492 5302 12548
rect 5358 12492 5426 12548
rect 5482 12492 5550 12548
rect 5606 12492 5674 12548
rect 5730 12492 5798 12548
rect 5854 12492 5922 12548
rect 5978 12492 6046 12548
rect 6102 12492 6170 12548
rect 6226 12492 6294 12548
rect 6350 12492 6418 12548
rect 6474 12492 6542 12548
rect 6598 12492 6666 12548
rect 6722 12492 6790 12548
rect 6846 12492 6914 12548
rect 6970 12492 7038 12548
rect 7094 12492 7104 12548
rect 5168 12424 7104 12492
rect 5168 12368 5178 12424
rect 5234 12368 5302 12424
rect 5358 12368 5426 12424
rect 5482 12368 5550 12424
rect 5606 12368 5674 12424
rect 5730 12368 5798 12424
rect 5854 12368 5922 12424
rect 5978 12368 6046 12424
rect 6102 12368 6170 12424
rect 6226 12368 6294 12424
rect 6350 12368 6418 12424
rect 6474 12368 6542 12424
rect 6598 12368 6666 12424
rect 6722 12368 6790 12424
rect 6846 12368 6914 12424
rect 6970 12368 7038 12424
rect 7094 12368 7104 12424
rect 5168 12300 7104 12368
rect 5168 12244 5178 12300
rect 5234 12244 5302 12300
rect 5358 12244 5426 12300
rect 5482 12244 5550 12300
rect 5606 12244 5674 12300
rect 5730 12244 5798 12300
rect 5854 12244 5922 12300
rect 5978 12244 6046 12300
rect 6102 12244 6170 12300
rect 6226 12244 6294 12300
rect 6350 12244 6418 12300
rect 6474 12244 6542 12300
rect 6598 12244 6666 12300
rect 6722 12244 6790 12300
rect 6846 12244 6914 12300
rect 6970 12244 7038 12300
rect 7094 12244 7104 12300
rect 5168 12176 7104 12244
rect 5168 12120 5178 12176
rect 5234 12120 5302 12176
rect 5358 12120 5426 12176
rect 5482 12120 5550 12176
rect 5606 12120 5674 12176
rect 5730 12120 5798 12176
rect 5854 12120 5922 12176
rect 5978 12120 6046 12176
rect 6102 12120 6170 12176
rect 6226 12120 6294 12176
rect 6350 12120 6418 12176
rect 6474 12120 6542 12176
rect 6598 12120 6666 12176
rect 6722 12120 6790 12176
rect 6846 12120 6914 12176
rect 6970 12120 7038 12176
rect 7094 12120 7104 12176
rect 5168 12052 7104 12120
rect 5168 11996 5178 12052
rect 5234 11996 5302 12052
rect 5358 11996 5426 12052
rect 5482 11996 5550 12052
rect 5606 11996 5674 12052
rect 5730 11996 5798 12052
rect 5854 11996 5922 12052
rect 5978 11996 6046 12052
rect 6102 11996 6170 12052
rect 6226 11996 6294 12052
rect 6350 11996 6418 12052
rect 6474 11996 6542 12052
rect 6598 11996 6666 12052
rect 6722 11996 6790 12052
rect 6846 11996 6914 12052
rect 6970 11996 7038 12052
rect 7094 11996 7104 12052
rect 5168 11928 7104 11996
rect 5168 11872 5178 11928
rect 5234 11872 5302 11928
rect 5358 11872 5426 11928
rect 5482 11872 5550 11928
rect 5606 11872 5674 11928
rect 5730 11872 5798 11928
rect 5854 11872 5922 11928
rect 5978 11872 6046 11928
rect 6102 11872 6170 11928
rect 6226 11872 6294 11928
rect 6350 11872 6418 11928
rect 6474 11872 6542 11928
rect 6598 11872 6666 11928
rect 6722 11872 6790 11928
rect 6846 11872 6914 11928
rect 6970 11872 7038 11928
rect 7094 11872 7104 11928
rect 5168 11804 7104 11872
rect 5168 11748 5178 11804
rect 5234 11748 5302 11804
rect 5358 11748 5426 11804
rect 5482 11748 5550 11804
rect 5606 11748 5674 11804
rect 5730 11748 5798 11804
rect 5854 11748 5922 11804
rect 5978 11748 6046 11804
rect 6102 11748 6170 11804
rect 6226 11748 6294 11804
rect 6350 11748 6418 11804
rect 6474 11748 6542 11804
rect 6598 11748 6666 11804
rect 6722 11748 6790 11804
rect 6846 11748 6914 11804
rect 6970 11748 7038 11804
rect 7094 11748 7104 11804
rect 5168 11680 7104 11748
rect 5168 11624 5178 11680
rect 5234 11624 5302 11680
rect 5358 11624 5426 11680
rect 5482 11624 5550 11680
rect 5606 11624 5674 11680
rect 5730 11624 5798 11680
rect 5854 11624 5922 11680
rect 5978 11624 6046 11680
rect 6102 11624 6170 11680
rect 6226 11624 6294 11680
rect 6350 11624 6418 11680
rect 6474 11624 6542 11680
rect 6598 11624 6666 11680
rect 6722 11624 6790 11680
rect 6846 11624 6914 11680
rect 6970 11624 7038 11680
rect 7094 11624 7104 11680
rect 5168 11556 7104 11624
rect 5168 11500 5178 11556
rect 5234 11500 5302 11556
rect 5358 11500 5426 11556
rect 5482 11500 5550 11556
rect 5606 11500 5674 11556
rect 5730 11500 5798 11556
rect 5854 11500 5922 11556
rect 5978 11500 6046 11556
rect 6102 11500 6170 11556
rect 6226 11500 6294 11556
rect 6350 11500 6418 11556
rect 6474 11500 6542 11556
rect 6598 11500 6666 11556
rect 6722 11500 6790 11556
rect 6846 11500 6914 11556
rect 6970 11500 7038 11556
rect 7094 11500 7104 11556
rect 5168 11432 7104 11500
rect 5168 11376 5178 11432
rect 5234 11376 5302 11432
rect 5358 11376 5426 11432
rect 5482 11376 5550 11432
rect 5606 11376 5674 11432
rect 5730 11376 5798 11432
rect 5854 11376 5922 11432
rect 5978 11376 6046 11432
rect 6102 11376 6170 11432
rect 6226 11376 6294 11432
rect 6350 11376 6418 11432
rect 6474 11376 6542 11432
rect 6598 11376 6666 11432
rect 6722 11376 6790 11432
rect 6846 11376 6914 11432
rect 6970 11376 7038 11432
rect 7094 11376 7104 11432
rect 5168 11308 7104 11376
rect 5168 11252 5178 11308
rect 5234 11252 5302 11308
rect 5358 11252 5426 11308
rect 5482 11252 5550 11308
rect 5606 11252 5674 11308
rect 5730 11252 5798 11308
rect 5854 11252 5922 11308
rect 5978 11252 6046 11308
rect 6102 11252 6170 11308
rect 6226 11252 6294 11308
rect 6350 11252 6418 11308
rect 6474 11252 6542 11308
rect 6598 11252 6666 11308
rect 6722 11252 6790 11308
rect 6846 11252 6914 11308
rect 6970 11252 7038 11308
rect 7094 11252 7104 11308
rect 5168 11242 7104 11252
rect 7874 12548 9810 12558
rect 7874 12492 7884 12548
rect 7940 12492 8008 12548
rect 8064 12492 8132 12548
rect 8188 12492 8256 12548
rect 8312 12492 8380 12548
rect 8436 12492 8504 12548
rect 8560 12492 8628 12548
rect 8684 12492 8752 12548
rect 8808 12492 8876 12548
rect 8932 12492 9000 12548
rect 9056 12492 9124 12548
rect 9180 12492 9248 12548
rect 9304 12492 9372 12548
rect 9428 12492 9496 12548
rect 9552 12492 9620 12548
rect 9676 12492 9744 12548
rect 9800 12492 9810 12548
rect 7874 12424 9810 12492
rect 7874 12368 7884 12424
rect 7940 12368 8008 12424
rect 8064 12368 8132 12424
rect 8188 12368 8256 12424
rect 8312 12368 8380 12424
rect 8436 12368 8504 12424
rect 8560 12368 8628 12424
rect 8684 12368 8752 12424
rect 8808 12368 8876 12424
rect 8932 12368 9000 12424
rect 9056 12368 9124 12424
rect 9180 12368 9248 12424
rect 9304 12368 9372 12424
rect 9428 12368 9496 12424
rect 9552 12368 9620 12424
rect 9676 12368 9744 12424
rect 9800 12368 9810 12424
rect 7874 12300 9810 12368
rect 7874 12244 7884 12300
rect 7940 12244 8008 12300
rect 8064 12244 8132 12300
rect 8188 12244 8256 12300
rect 8312 12244 8380 12300
rect 8436 12244 8504 12300
rect 8560 12244 8628 12300
rect 8684 12244 8752 12300
rect 8808 12244 8876 12300
rect 8932 12244 9000 12300
rect 9056 12244 9124 12300
rect 9180 12244 9248 12300
rect 9304 12244 9372 12300
rect 9428 12244 9496 12300
rect 9552 12244 9620 12300
rect 9676 12244 9744 12300
rect 9800 12244 9810 12300
rect 7874 12176 9810 12244
rect 7874 12120 7884 12176
rect 7940 12120 8008 12176
rect 8064 12120 8132 12176
rect 8188 12120 8256 12176
rect 8312 12120 8380 12176
rect 8436 12120 8504 12176
rect 8560 12120 8628 12176
rect 8684 12120 8752 12176
rect 8808 12120 8876 12176
rect 8932 12120 9000 12176
rect 9056 12120 9124 12176
rect 9180 12120 9248 12176
rect 9304 12120 9372 12176
rect 9428 12120 9496 12176
rect 9552 12120 9620 12176
rect 9676 12120 9744 12176
rect 9800 12120 9810 12176
rect 7874 12052 9810 12120
rect 7874 11996 7884 12052
rect 7940 11996 8008 12052
rect 8064 11996 8132 12052
rect 8188 11996 8256 12052
rect 8312 11996 8380 12052
rect 8436 11996 8504 12052
rect 8560 11996 8628 12052
rect 8684 11996 8752 12052
rect 8808 11996 8876 12052
rect 8932 11996 9000 12052
rect 9056 11996 9124 12052
rect 9180 11996 9248 12052
rect 9304 11996 9372 12052
rect 9428 11996 9496 12052
rect 9552 11996 9620 12052
rect 9676 11996 9744 12052
rect 9800 11996 9810 12052
rect 7874 11928 9810 11996
rect 7874 11872 7884 11928
rect 7940 11872 8008 11928
rect 8064 11872 8132 11928
rect 8188 11872 8256 11928
rect 8312 11872 8380 11928
rect 8436 11872 8504 11928
rect 8560 11872 8628 11928
rect 8684 11872 8752 11928
rect 8808 11872 8876 11928
rect 8932 11872 9000 11928
rect 9056 11872 9124 11928
rect 9180 11872 9248 11928
rect 9304 11872 9372 11928
rect 9428 11872 9496 11928
rect 9552 11872 9620 11928
rect 9676 11872 9744 11928
rect 9800 11872 9810 11928
rect 7874 11804 9810 11872
rect 7874 11748 7884 11804
rect 7940 11748 8008 11804
rect 8064 11748 8132 11804
rect 8188 11748 8256 11804
rect 8312 11748 8380 11804
rect 8436 11748 8504 11804
rect 8560 11748 8628 11804
rect 8684 11748 8752 11804
rect 8808 11748 8876 11804
rect 8932 11748 9000 11804
rect 9056 11748 9124 11804
rect 9180 11748 9248 11804
rect 9304 11748 9372 11804
rect 9428 11748 9496 11804
rect 9552 11748 9620 11804
rect 9676 11748 9744 11804
rect 9800 11748 9810 11804
rect 7874 11680 9810 11748
rect 7874 11624 7884 11680
rect 7940 11624 8008 11680
rect 8064 11624 8132 11680
rect 8188 11624 8256 11680
rect 8312 11624 8380 11680
rect 8436 11624 8504 11680
rect 8560 11624 8628 11680
rect 8684 11624 8752 11680
rect 8808 11624 8876 11680
rect 8932 11624 9000 11680
rect 9056 11624 9124 11680
rect 9180 11624 9248 11680
rect 9304 11624 9372 11680
rect 9428 11624 9496 11680
rect 9552 11624 9620 11680
rect 9676 11624 9744 11680
rect 9800 11624 9810 11680
rect 7874 11556 9810 11624
rect 7874 11500 7884 11556
rect 7940 11500 8008 11556
rect 8064 11500 8132 11556
rect 8188 11500 8256 11556
rect 8312 11500 8380 11556
rect 8436 11500 8504 11556
rect 8560 11500 8628 11556
rect 8684 11500 8752 11556
rect 8808 11500 8876 11556
rect 8932 11500 9000 11556
rect 9056 11500 9124 11556
rect 9180 11500 9248 11556
rect 9304 11500 9372 11556
rect 9428 11500 9496 11556
rect 9552 11500 9620 11556
rect 9676 11500 9744 11556
rect 9800 11500 9810 11556
rect 7874 11432 9810 11500
rect 7874 11376 7884 11432
rect 7940 11376 8008 11432
rect 8064 11376 8132 11432
rect 8188 11376 8256 11432
rect 8312 11376 8380 11432
rect 8436 11376 8504 11432
rect 8560 11376 8628 11432
rect 8684 11376 8752 11432
rect 8808 11376 8876 11432
rect 8932 11376 9000 11432
rect 9056 11376 9124 11432
rect 9180 11376 9248 11432
rect 9304 11376 9372 11432
rect 9428 11376 9496 11432
rect 9552 11376 9620 11432
rect 9676 11376 9744 11432
rect 9800 11376 9810 11432
rect 7874 11308 9810 11376
rect 7874 11252 7884 11308
rect 7940 11252 8008 11308
rect 8064 11252 8132 11308
rect 8188 11252 8256 11308
rect 8312 11252 8380 11308
rect 8436 11252 8504 11308
rect 8560 11252 8628 11308
rect 8684 11252 8752 11308
rect 8808 11252 8876 11308
rect 8932 11252 9000 11308
rect 9056 11252 9124 11308
rect 9180 11252 9248 11308
rect 9304 11252 9372 11308
rect 9428 11252 9496 11308
rect 9552 11252 9620 11308
rect 9676 11252 9744 11308
rect 9800 11252 9810 11308
rect 7874 11242 9810 11252
rect 10244 12548 12180 12558
rect 10244 12492 10254 12548
rect 10310 12492 10378 12548
rect 10434 12492 10502 12548
rect 10558 12492 10626 12548
rect 10682 12492 10750 12548
rect 10806 12492 10874 12548
rect 10930 12492 10998 12548
rect 11054 12492 11122 12548
rect 11178 12492 11246 12548
rect 11302 12492 11370 12548
rect 11426 12492 11494 12548
rect 11550 12492 11618 12548
rect 11674 12492 11742 12548
rect 11798 12492 11866 12548
rect 11922 12492 11990 12548
rect 12046 12492 12114 12548
rect 12170 12492 12180 12548
rect 10244 12424 12180 12492
rect 10244 12368 10254 12424
rect 10310 12368 10378 12424
rect 10434 12368 10502 12424
rect 10558 12368 10626 12424
rect 10682 12368 10750 12424
rect 10806 12368 10874 12424
rect 10930 12368 10998 12424
rect 11054 12368 11122 12424
rect 11178 12368 11246 12424
rect 11302 12368 11370 12424
rect 11426 12368 11494 12424
rect 11550 12368 11618 12424
rect 11674 12368 11742 12424
rect 11798 12368 11866 12424
rect 11922 12368 11990 12424
rect 12046 12368 12114 12424
rect 12170 12368 12180 12424
rect 10244 12300 12180 12368
rect 10244 12244 10254 12300
rect 10310 12244 10378 12300
rect 10434 12244 10502 12300
rect 10558 12244 10626 12300
rect 10682 12244 10750 12300
rect 10806 12244 10874 12300
rect 10930 12244 10998 12300
rect 11054 12244 11122 12300
rect 11178 12244 11246 12300
rect 11302 12244 11370 12300
rect 11426 12244 11494 12300
rect 11550 12244 11618 12300
rect 11674 12244 11742 12300
rect 11798 12244 11866 12300
rect 11922 12244 11990 12300
rect 12046 12244 12114 12300
rect 12170 12244 12180 12300
rect 10244 12176 12180 12244
rect 10244 12120 10254 12176
rect 10310 12120 10378 12176
rect 10434 12120 10502 12176
rect 10558 12120 10626 12176
rect 10682 12120 10750 12176
rect 10806 12120 10874 12176
rect 10930 12120 10998 12176
rect 11054 12120 11122 12176
rect 11178 12120 11246 12176
rect 11302 12120 11370 12176
rect 11426 12120 11494 12176
rect 11550 12120 11618 12176
rect 11674 12120 11742 12176
rect 11798 12120 11866 12176
rect 11922 12120 11990 12176
rect 12046 12120 12114 12176
rect 12170 12120 12180 12176
rect 10244 12052 12180 12120
rect 10244 11996 10254 12052
rect 10310 11996 10378 12052
rect 10434 11996 10502 12052
rect 10558 11996 10626 12052
rect 10682 11996 10750 12052
rect 10806 11996 10874 12052
rect 10930 11996 10998 12052
rect 11054 11996 11122 12052
rect 11178 11996 11246 12052
rect 11302 11996 11370 12052
rect 11426 11996 11494 12052
rect 11550 11996 11618 12052
rect 11674 11996 11742 12052
rect 11798 11996 11866 12052
rect 11922 11996 11990 12052
rect 12046 11996 12114 12052
rect 12170 11996 12180 12052
rect 10244 11928 12180 11996
rect 10244 11872 10254 11928
rect 10310 11872 10378 11928
rect 10434 11872 10502 11928
rect 10558 11872 10626 11928
rect 10682 11872 10750 11928
rect 10806 11872 10874 11928
rect 10930 11872 10998 11928
rect 11054 11872 11122 11928
rect 11178 11872 11246 11928
rect 11302 11872 11370 11928
rect 11426 11872 11494 11928
rect 11550 11872 11618 11928
rect 11674 11872 11742 11928
rect 11798 11872 11866 11928
rect 11922 11872 11990 11928
rect 12046 11872 12114 11928
rect 12170 11872 12180 11928
rect 10244 11804 12180 11872
rect 10244 11748 10254 11804
rect 10310 11748 10378 11804
rect 10434 11748 10502 11804
rect 10558 11748 10626 11804
rect 10682 11748 10750 11804
rect 10806 11748 10874 11804
rect 10930 11748 10998 11804
rect 11054 11748 11122 11804
rect 11178 11748 11246 11804
rect 11302 11748 11370 11804
rect 11426 11748 11494 11804
rect 11550 11748 11618 11804
rect 11674 11748 11742 11804
rect 11798 11748 11866 11804
rect 11922 11748 11990 11804
rect 12046 11748 12114 11804
rect 12170 11748 12180 11804
rect 10244 11680 12180 11748
rect 10244 11624 10254 11680
rect 10310 11624 10378 11680
rect 10434 11624 10502 11680
rect 10558 11624 10626 11680
rect 10682 11624 10750 11680
rect 10806 11624 10874 11680
rect 10930 11624 10998 11680
rect 11054 11624 11122 11680
rect 11178 11624 11246 11680
rect 11302 11624 11370 11680
rect 11426 11624 11494 11680
rect 11550 11624 11618 11680
rect 11674 11624 11742 11680
rect 11798 11624 11866 11680
rect 11922 11624 11990 11680
rect 12046 11624 12114 11680
rect 12170 11624 12180 11680
rect 10244 11556 12180 11624
rect 10244 11500 10254 11556
rect 10310 11500 10378 11556
rect 10434 11500 10502 11556
rect 10558 11500 10626 11556
rect 10682 11500 10750 11556
rect 10806 11500 10874 11556
rect 10930 11500 10998 11556
rect 11054 11500 11122 11556
rect 11178 11500 11246 11556
rect 11302 11500 11370 11556
rect 11426 11500 11494 11556
rect 11550 11500 11618 11556
rect 11674 11500 11742 11556
rect 11798 11500 11866 11556
rect 11922 11500 11990 11556
rect 12046 11500 12114 11556
rect 12170 11500 12180 11556
rect 10244 11432 12180 11500
rect 10244 11376 10254 11432
rect 10310 11376 10378 11432
rect 10434 11376 10502 11432
rect 10558 11376 10626 11432
rect 10682 11376 10750 11432
rect 10806 11376 10874 11432
rect 10930 11376 10998 11432
rect 11054 11376 11122 11432
rect 11178 11376 11246 11432
rect 11302 11376 11370 11432
rect 11426 11376 11494 11432
rect 11550 11376 11618 11432
rect 11674 11376 11742 11432
rect 11798 11376 11866 11432
rect 11922 11376 11990 11432
rect 12046 11376 12114 11432
rect 12170 11376 12180 11432
rect 10244 11308 12180 11376
rect 10244 11252 10254 11308
rect 10310 11252 10378 11308
rect 10434 11252 10502 11308
rect 10558 11252 10626 11308
rect 10682 11252 10750 11308
rect 10806 11252 10874 11308
rect 10930 11252 10998 11308
rect 11054 11252 11122 11308
rect 11178 11252 11246 11308
rect 11302 11252 11370 11308
rect 11426 11252 11494 11308
rect 11550 11252 11618 11308
rect 11674 11252 11742 11308
rect 11798 11252 11866 11308
rect 11922 11252 11990 11308
rect 12046 11252 12114 11308
rect 12170 11252 12180 11308
rect 10244 11242 12180 11252
rect 12861 12548 14673 12558
rect 12861 12492 12871 12548
rect 12927 12492 12995 12548
rect 13051 12492 13119 12548
rect 13175 12492 13243 12548
rect 13299 12492 13367 12548
rect 13423 12492 13491 12548
rect 13547 12492 13615 12548
rect 13671 12492 13739 12548
rect 13795 12492 13863 12548
rect 13919 12492 13987 12548
rect 14043 12492 14111 12548
rect 14167 12492 14235 12548
rect 14291 12492 14359 12548
rect 14415 12492 14483 12548
rect 14539 12492 14607 12548
rect 14663 12492 14673 12548
rect 12861 12424 14673 12492
rect 12861 12368 12871 12424
rect 12927 12368 12995 12424
rect 13051 12368 13119 12424
rect 13175 12368 13243 12424
rect 13299 12368 13367 12424
rect 13423 12368 13491 12424
rect 13547 12368 13615 12424
rect 13671 12368 13739 12424
rect 13795 12368 13863 12424
rect 13919 12368 13987 12424
rect 14043 12368 14111 12424
rect 14167 12368 14235 12424
rect 14291 12368 14359 12424
rect 14415 12368 14483 12424
rect 14539 12368 14607 12424
rect 14663 12368 14673 12424
rect 12861 12300 14673 12368
rect 12861 12244 12871 12300
rect 12927 12244 12995 12300
rect 13051 12244 13119 12300
rect 13175 12244 13243 12300
rect 13299 12244 13367 12300
rect 13423 12244 13491 12300
rect 13547 12244 13615 12300
rect 13671 12244 13739 12300
rect 13795 12244 13863 12300
rect 13919 12244 13987 12300
rect 14043 12244 14111 12300
rect 14167 12244 14235 12300
rect 14291 12244 14359 12300
rect 14415 12244 14483 12300
rect 14539 12244 14607 12300
rect 14663 12244 14673 12300
rect 12861 12176 14673 12244
rect 12861 12120 12871 12176
rect 12927 12120 12995 12176
rect 13051 12120 13119 12176
rect 13175 12120 13243 12176
rect 13299 12120 13367 12176
rect 13423 12120 13491 12176
rect 13547 12120 13615 12176
rect 13671 12120 13739 12176
rect 13795 12120 13863 12176
rect 13919 12120 13987 12176
rect 14043 12120 14111 12176
rect 14167 12120 14235 12176
rect 14291 12120 14359 12176
rect 14415 12120 14483 12176
rect 14539 12120 14607 12176
rect 14663 12120 14673 12176
rect 12861 12052 14673 12120
rect 12861 11996 12871 12052
rect 12927 11996 12995 12052
rect 13051 11996 13119 12052
rect 13175 11996 13243 12052
rect 13299 11996 13367 12052
rect 13423 11996 13491 12052
rect 13547 11996 13615 12052
rect 13671 11996 13739 12052
rect 13795 11996 13863 12052
rect 13919 11996 13987 12052
rect 14043 11996 14111 12052
rect 14167 11996 14235 12052
rect 14291 11996 14359 12052
rect 14415 11996 14483 12052
rect 14539 11996 14607 12052
rect 14663 11996 14673 12052
rect 12861 11928 14673 11996
rect 12861 11872 12871 11928
rect 12927 11872 12995 11928
rect 13051 11872 13119 11928
rect 13175 11872 13243 11928
rect 13299 11872 13367 11928
rect 13423 11872 13491 11928
rect 13547 11872 13615 11928
rect 13671 11872 13739 11928
rect 13795 11872 13863 11928
rect 13919 11872 13987 11928
rect 14043 11872 14111 11928
rect 14167 11872 14235 11928
rect 14291 11872 14359 11928
rect 14415 11872 14483 11928
rect 14539 11872 14607 11928
rect 14663 11872 14673 11928
rect 12861 11804 14673 11872
rect 12861 11748 12871 11804
rect 12927 11748 12995 11804
rect 13051 11748 13119 11804
rect 13175 11748 13243 11804
rect 13299 11748 13367 11804
rect 13423 11748 13491 11804
rect 13547 11748 13615 11804
rect 13671 11748 13739 11804
rect 13795 11748 13863 11804
rect 13919 11748 13987 11804
rect 14043 11748 14111 11804
rect 14167 11748 14235 11804
rect 14291 11748 14359 11804
rect 14415 11748 14483 11804
rect 14539 11748 14607 11804
rect 14663 11748 14673 11804
rect 12861 11680 14673 11748
rect 12861 11624 12871 11680
rect 12927 11624 12995 11680
rect 13051 11624 13119 11680
rect 13175 11624 13243 11680
rect 13299 11624 13367 11680
rect 13423 11624 13491 11680
rect 13547 11624 13615 11680
rect 13671 11624 13739 11680
rect 13795 11624 13863 11680
rect 13919 11624 13987 11680
rect 14043 11624 14111 11680
rect 14167 11624 14235 11680
rect 14291 11624 14359 11680
rect 14415 11624 14483 11680
rect 14539 11624 14607 11680
rect 14663 11624 14673 11680
rect 12861 11556 14673 11624
rect 12861 11500 12871 11556
rect 12927 11500 12995 11556
rect 13051 11500 13119 11556
rect 13175 11500 13243 11556
rect 13299 11500 13367 11556
rect 13423 11500 13491 11556
rect 13547 11500 13615 11556
rect 13671 11500 13739 11556
rect 13795 11500 13863 11556
rect 13919 11500 13987 11556
rect 14043 11500 14111 11556
rect 14167 11500 14235 11556
rect 14291 11500 14359 11556
rect 14415 11500 14483 11556
rect 14539 11500 14607 11556
rect 14663 11500 14673 11556
rect 12861 11432 14673 11500
rect 12861 11376 12871 11432
rect 12927 11376 12995 11432
rect 13051 11376 13119 11432
rect 13175 11376 13243 11432
rect 13299 11376 13367 11432
rect 13423 11376 13491 11432
rect 13547 11376 13615 11432
rect 13671 11376 13739 11432
rect 13795 11376 13863 11432
rect 13919 11376 13987 11432
rect 14043 11376 14111 11432
rect 14167 11376 14235 11432
rect 14291 11376 14359 11432
rect 14415 11376 14483 11432
rect 14539 11376 14607 11432
rect 14663 11376 14673 11432
rect 12861 11308 14673 11376
rect 12861 11252 12871 11308
rect 12927 11252 12995 11308
rect 13051 11252 13119 11308
rect 13175 11252 13243 11308
rect 13299 11252 13367 11308
rect 13423 11252 13491 11308
rect 13547 11252 13615 11308
rect 13671 11252 13739 11308
rect 13795 11252 13863 11308
rect 13919 11252 13987 11308
rect 14043 11252 14111 11308
rect 14167 11252 14235 11308
rect 14291 11252 14359 11308
rect 14415 11252 14483 11308
rect 14539 11252 14607 11308
rect 14663 11252 14673 11308
rect 12861 11242 14673 11252
rect 2481 10954 2681 10964
rect 2481 10898 2491 10954
rect 2547 10898 2615 10954
rect 2671 10898 2681 10954
rect 2481 10830 2681 10898
rect 2481 10774 2491 10830
rect 2547 10774 2615 10830
rect 2671 10774 2681 10830
rect 2481 10706 2681 10774
rect 2481 10650 2491 10706
rect 2547 10650 2615 10706
rect 2671 10650 2681 10706
rect 2481 10582 2681 10650
rect 2481 10526 2491 10582
rect 2547 10526 2615 10582
rect 2671 10526 2681 10582
rect 2481 10458 2681 10526
rect 2481 10402 2491 10458
rect 2547 10402 2615 10458
rect 2671 10402 2681 10458
rect 2481 10334 2681 10402
rect 2481 10278 2491 10334
rect 2547 10278 2615 10334
rect 2671 10278 2681 10334
rect 2481 10210 2681 10278
rect 2481 10154 2491 10210
rect 2547 10154 2615 10210
rect 2671 10154 2681 10210
rect 2481 10086 2681 10154
rect 2481 10030 2491 10086
rect 2547 10030 2615 10086
rect 2671 10030 2681 10086
rect 2481 9962 2681 10030
rect 2481 9906 2491 9962
rect 2547 9906 2615 9962
rect 2671 9906 2681 9962
rect 2481 9838 2681 9906
rect 2481 9782 2491 9838
rect 2547 9782 2615 9838
rect 2671 9782 2681 9838
rect 2481 9714 2681 9782
rect 2481 9658 2491 9714
rect 2547 9658 2615 9714
rect 2671 9658 2681 9714
rect 2481 9590 2681 9658
rect 2481 9534 2491 9590
rect 2547 9534 2615 9590
rect 2671 9534 2681 9590
rect 2481 9466 2681 9534
rect 2481 9410 2491 9466
rect 2547 9410 2615 9466
rect 2671 9410 2681 9466
rect 2481 9342 2681 9410
rect 2481 9286 2491 9342
rect 2547 9286 2615 9342
rect 2671 9286 2681 9342
rect 2481 9218 2681 9286
rect 2481 9162 2491 9218
rect 2547 9162 2615 9218
rect 2671 9162 2681 9218
rect 2481 9094 2681 9162
rect 2481 9038 2491 9094
rect 2547 9038 2615 9094
rect 2671 9038 2681 9094
rect 2481 8970 2681 9038
rect 2481 8914 2491 8970
rect 2547 8914 2615 8970
rect 2671 8914 2681 8970
rect 2481 8846 2681 8914
rect 2481 8790 2491 8846
rect 2547 8790 2615 8846
rect 2671 8790 2681 8846
rect 2481 8722 2681 8790
rect 2481 8666 2491 8722
rect 2547 8666 2615 8722
rect 2671 8666 2681 8722
rect 2481 8598 2681 8666
rect 2481 8542 2491 8598
rect 2547 8542 2615 8598
rect 2671 8542 2681 8598
rect 2481 8474 2681 8542
rect 2481 8418 2491 8474
rect 2547 8418 2615 8474
rect 2671 8418 2681 8474
rect 2481 8350 2681 8418
rect 2481 8294 2491 8350
rect 2547 8294 2615 8350
rect 2671 8294 2681 8350
rect 2481 8226 2681 8294
rect 2481 8170 2491 8226
rect 2547 8170 2615 8226
rect 2671 8170 2681 8226
rect 2481 8102 2681 8170
rect 2481 8046 2491 8102
rect 2547 8046 2615 8102
rect 2671 8046 2681 8102
rect 2481 8036 2681 8046
rect 4851 10954 5051 10964
rect 4851 10898 4861 10954
rect 4917 10898 4985 10954
rect 5041 10898 5051 10954
rect 4851 10830 5051 10898
rect 4851 10774 4861 10830
rect 4917 10774 4985 10830
rect 5041 10774 5051 10830
rect 4851 10706 5051 10774
rect 4851 10650 4861 10706
rect 4917 10650 4985 10706
rect 5041 10650 5051 10706
rect 4851 10582 5051 10650
rect 4851 10526 4861 10582
rect 4917 10526 4985 10582
rect 5041 10526 5051 10582
rect 4851 10458 5051 10526
rect 4851 10402 4861 10458
rect 4917 10402 4985 10458
rect 5041 10402 5051 10458
rect 4851 10334 5051 10402
rect 4851 10278 4861 10334
rect 4917 10278 4985 10334
rect 5041 10278 5051 10334
rect 4851 10210 5051 10278
rect 4851 10154 4861 10210
rect 4917 10154 4985 10210
rect 5041 10154 5051 10210
rect 4851 10086 5051 10154
rect 4851 10030 4861 10086
rect 4917 10030 4985 10086
rect 5041 10030 5051 10086
rect 4851 9962 5051 10030
rect 4851 9906 4861 9962
rect 4917 9906 4985 9962
rect 5041 9906 5051 9962
rect 4851 9838 5051 9906
rect 4851 9782 4861 9838
rect 4917 9782 4985 9838
rect 5041 9782 5051 9838
rect 4851 9714 5051 9782
rect 4851 9658 4861 9714
rect 4917 9658 4985 9714
rect 5041 9658 5051 9714
rect 4851 9590 5051 9658
rect 4851 9534 4861 9590
rect 4917 9534 4985 9590
rect 5041 9534 5051 9590
rect 4851 9466 5051 9534
rect 4851 9410 4861 9466
rect 4917 9410 4985 9466
rect 5041 9410 5051 9466
rect 4851 9342 5051 9410
rect 4851 9286 4861 9342
rect 4917 9286 4985 9342
rect 5041 9286 5051 9342
rect 4851 9218 5051 9286
rect 4851 9162 4861 9218
rect 4917 9162 4985 9218
rect 5041 9162 5051 9218
rect 4851 9094 5051 9162
rect 4851 9038 4861 9094
rect 4917 9038 4985 9094
rect 5041 9038 5051 9094
rect 4851 8970 5051 9038
rect 4851 8914 4861 8970
rect 4917 8914 4985 8970
rect 5041 8914 5051 8970
rect 4851 8846 5051 8914
rect 4851 8790 4861 8846
rect 4917 8790 4985 8846
rect 5041 8790 5051 8846
rect 4851 8722 5051 8790
rect 4851 8666 4861 8722
rect 4917 8666 4985 8722
rect 5041 8666 5051 8722
rect 4851 8598 5051 8666
rect 4851 8542 4861 8598
rect 4917 8542 4985 8598
rect 5041 8542 5051 8598
rect 4851 8474 5051 8542
rect 4851 8418 4861 8474
rect 4917 8418 4985 8474
rect 5041 8418 5051 8474
rect 4851 8350 5051 8418
rect 4851 8294 4861 8350
rect 4917 8294 4985 8350
rect 5041 8294 5051 8350
rect 4851 8226 5051 8294
rect 4851 8170 4861 8226
rect 4917 8170 4985 8226
rect 5041 8170 5051 8226
rect 4851 8102 5051 8170
rect 4851 8046 4861 8102
rect 4917 8046 4985 8102
rect 5041 8046 5051 8102
rect 4851 8036 5051 8046
rect 7265 10954 7713 10964
rect 7265 10898 7275 10954
rect 7331 10898 7399 10954
rect 7455 10898 7523 10954
rect 7579 10898 7647 10954
rect 7703 10898 7713 10954
rect 7265 10830 7713 10898
rect 7265 10774 7275 10830
rect 7331 10774 7399 10830
rect 7455 10774 7523 10830
rect 7579 10774 7647 10830
rect 7703 10774 7713 10830
rect 7265 10706 7713 10774
rect 7265 10650 7275 10706
rect 7331 10650 7399 10706
rect 7455 10650 7523 10706
rect 7579 10650 7647 10706
rect 7703 10650 7713 10706
rect 7265 10582 7713 10650
rect 7265 10526 7275 10582
rect 7331 10526 7399 10582
rect 7455 10526 7523 10582
rect 7579 10526 7647 10582
rect 7703 10526 7713 10582
rect 7265 10458 7713 10526
rect 7265 10402 7275 10458
rect 7331 10402 7399 10458
rect 7455 10402 7523 10458
rect 7579 10402 7647 10458
rect 7703 10402 7713 10458
rect 7265 10334 7713 10402
rect 7265 10278 7275 10334
rect 7331 10278 7399 10334
rect 7455 10278 7523 10334
rect 7579 10278 7647 10334
rect 7703 10278 7713 10334
rect 7265 10210 7713 10278
rect 7265 10154 7275 10210
rect 7331 10154 7399 10210
rect 7455 10154 7523 10210
rect 7579 10154 7647 10210
rect 7703 10154 7713 10210
rect 7265 10086 7713 10154
rect 7265 10030 7275 10086
rect 7331 10030 7399 10086
rect 7455 10030 7523 10086
rect 7579 10030 7647 10086
rect 7703 10030 7713 10086
rect 7265 9962 7713 10030
rect 7265 9906 7275 9962
rect 7331 9906 7399 9962
rect 7455 9906 7523 9962
rect 7579 9906 7647 9962
rect 7703 9906 7713 9962
rect 7265 9838 7713 9906
rect 7265 9782 7275 9838
rect 7331 9782 7399 9838
rect 7455 9782 7523 9838
rect 7579 9782 7647 9838
rect 7703 9782 7713 9838
rect 7265 9714 7713 9782
rect 7265 9658 7275 9714
rect 7331 9658 7399 9714
rect 7455 9658 7523 9714
rect 7579 9658 7647 9714
rect 7703 9658 7713 9714
rect 7265 9590 7713 9658
rect 7265 9534 7275 9590
rect 7331 9534 7399 9590
rect 7455 9534 7523 9590
rect 7579 9534 7647 9590
rect 7703 9534 7713 9590
rect 7265 9466 7713 9534
rect 7265 9410 7275 9466
rect 7331 9410 7399 9466
rect 7455 9410 7523 9466
rect 7579 9410 7647 9466
rect 7703 9410 7713 9466
rect 7265 9342 7713 9410
rect 7265 9286 7275 9342
rect 7331 9286 7399 9342
rect 7455 9286 7523 9342
rect 7579 9286 7647 9342
rect 7703 9286 7713 9342
rect 7265 9218 7713 9286
rect 7265 9162 7275 9218
rect 7331 9162 7399 9218
rect 7455 9162 7523 9218
rect 7579 9162 7647 9218
rect 7703 9162 7713 9218
rect 7265 9094 7713 9162
rect 7265 9038 7275 9094
rect 7331 9038 7399 9094
rect 7455 9038 7523 9094
rect 7579 9038 7647 9094
rect 7703 9038 7713 9094
rect 7265 8970 7713 9038
rect 7265 8914 7275 8970
rect 7331 8914 7399 8970
rect 7455 8914 7523 8970
rect 7579 8914 7647 8970
rect 7703 8914 7713 8970
rect 7265 8846 7713 8914
rect 7265 8790 7275 8846
rect 7331 8790 7399 8846
rect 7455 8790 7523 8846
rect 7579 8790 7647 8846
rect 7703 8790 7713 8846
rect 7265 8722 7713 8790
rect 7265 8666 7275 8722
rect 7331 8666 7399 8722
rect 7455 8666 7523 8722
rect 7579 8666 7647 8722
rect 7703 8666 7713 8722
rect 7265 8598 7713 8666
rect 7265 8542 7275 8598
rect 7331 8542 7399 8598
rect 7455 8542 7523 8598
rect 7579 8542 7647 8598
rect 7703 8542 7713 8598
rect 7265 8474 7713 8542
rect 7265 8418 7275 8474
rect 7331 8418 7399 8474
rect 7455 8418 7523 8474
rect 7579 8418 7647 8474
rect 7703 8418 7713 8474
rect 7265 8350 7713 8418
rect 7265 8294 7275 8350
rect 7331 8294 7399 8350
rect 7455 8294 7523 8350
rect 7579 8294 7647 8350
rect 7703 8294 7713 8350
rect 7265 8226 7713 8294
rect 7265 8170 7275 8226
rect 7331 8170 7399 8226
rect 7455 8170 7523 8226
rect 7579 8170 7647 8226
rect 7703 8170 7713 8226
rect 7265 8102 7713 8170
rect 7265 8046 7275 8102
rect 7331 8046 7399 8102
rect 7455 8046 7523 8102
rect 7579 8046 7647 8102
rect 7703 8046 7713 8102
rect 7265 8036 7713 8046
rect 9927 10954 10127 10964
rect 9927 10898 9937 10954
rect 9993 10898 10061 10954
rect 10117 10898 10127 10954
rect 9927 10830 10127 10898
rect 9927 10774 9937 10830
rect 9993 10774 10061 10830
rect 10117 10774 10127 10830
rect 9927 10706 10127 10774
rect 9927 10650 9937 10706
rect 9993 10650 10061 10706
rect 10117 10650 10127 10706
rect 9927 10582 10127 10650
rect 9927 10526 9937 10582
rect 9993 10526 10061 10582
rect 10117 10526 10127 10582
rect 9927 10458 10127 10526
rect 9927 10402 9937 10458
rect 9993 10402 10061 10458
rect 10117 10402 10127 10458
rect 9927 10334 10127 10402
rect 9927 10278 9937 10334
rect 9993 10278 10061 10334
rect 10117 10278 10127 10334
rect 9927 10210 10127 10278
rect 9927 10154 9937 10210
rect 9993 10154 10061 10210
rect 10117 10154 10127 10210
rect 9927 10086 10127 10154
rect 9927 10030 9937 10086
rect 9993 10030 10061 10086
rect 10117 10030 10127 10086
rect 9927 9962 10127 10030
rect 9927 9906 9937 9962
rect 9993 9906 10061 9962
rect 10117 9906 10127 9962
rect 9927 9838 10127 9906
rect 9927 9782 9937 9838
rect 9993 9782 10061 9838
rect 10117 9782 10127 9838
rect 9927 9714 10127 9782
rect 9927 9658 9937 9714
rect 9993 9658 10061 9714
rect 10117 9658 10127 9714
rect 9927 9590 10127 9658
rect 9927 9534 9937 9590
rect 9993 9534 10061 9590
rect 10117 9534 10127 9590
rect 9927 9466 10127 9534
rect 9927 9410 9937 9466
rect 9993 9410 10061 9466
rect 10117 9410 10127 9466
rect 9927 9342 10127 9410
rect 9927 9286 9937 9342
rect 9993 9286 10061 9342
rect 10117 9286 10127 9342
rect 9927 9218 10127 9286
rect 9927 9162 9937 9218
rect 9993 9162 10061 9218
rect 10117 9162 10127 9218
rect 9927 9094 10127 9162
rect 9927 9038 9937 9094
rect 9993 9038 10061 9094
rect 10117 9038 10127 9094
rect 9927 8970 10127 9038
rect 9927 8914 9937 8970
rect 9993 8914 10061 8970
rect 10117 8914 10127 8970
rect 9927 8846 10127 8914
rect 9927 8790 9937 8846
rect 9993 8790 10061 8846
rect 10117 8790 10127 8846
rect 9927 8722 10127 8790
rect 9927 8666 9937 8722
rect 9993 8666 10061 8722
rect 10117 8666 10127 8722
rect 9927 8598 10127 8666
rect 9927 8542 9937 8598
rect 9993 8542 10061 8598
rect 10117 8542 10127 8598
rect 9927 8474 10127 8542
rect 9927 8418 9937 8474
rect 9993 8418 10061 8474
rect 10117 8418 10127 8474
rect 9927 8350 10127 8418
rect 9927 8294 9937 8350
rect 9993 8294 10061 8350
rect 10117 8294 10127 8350
rect 9927 8226 10127 8294
rect 9927 8170 9937 8226
rect 9993 8170 10061 8226
rect 10117 8170 10127 8226
rect 9927 8102 10127 8170
rect 9927 8046 9937 8102
rect 9993 8046 10061 8102
rect 10117 8046 10127 8102
rect 9927 8036 10127 8046
rect 12297 10954 12497 10964
rect 12297 10898 12307 10954
rect 12363 10898 12431 10954
rect 12487 10898 12497 10954
rect 12297 10830 12497 10898
rect 12297 10774 12307 10830
rect 12363 10774 12431 10830
rect 12487 10774 12497 10830
rect 12297 10706 12497 10774
rect 12297 10650 12307 10706
rect 12363 10650 12431 10706
rect 12487 10650 12497 10706
rect 12297 10582 12497 10650
rect 12297 10526 12307 10582
rect 12363 10526 12431 10582
rect 12487 10526 12497 10582
rect 12297 10458 12497 10526
rect 12297 10402 12307 10458
rect 12363 10402 12431 10458
rect 12487 10402 12497 10458
rect 12297 10334 12497 10402
rect 12297 10278 12307 10334
rect 12363 10278 12431 10334
rect 12487 10278 12497 10334
rect 12297 10210 12497 10278
rect 12297 10154 12307 10210
rect 12363 10154 12431 10210
rect 12487 10154 12497 10210
rect 12297 10086 12497 10154
rect 12297 10030 12307 10086
rect 12363 10030 12431 10086
rect 12487 10030 12497 10086
rect 12297 9962 12497 10030
rect 12297 9906 12307 9962
rect 12363 9906 12431 9962
rect 12487 9906 12497 9962
rect 12297 9838 12497 9906
rect 12297 9782 12307 9838
rect 12363 9782 12431 9838
rect 12487 9782 12497 9838
rect 12297 9714 12497 9782
rect 12297 9658 12307 9714
rect 12363 9658 12431 9714
rect 12487 9658 12497 9714
rect 12297 9590 12497 9658
rect 12297 9534 12307 9590
rect 12363 9534 12431 9590
rect 12487 9534 12497 9590
rect 12297 9466 12497 9534
rect 12297 9410 12307 9466
rect 12363 9410 12431 9466
rect 12487 9410 12497 9466
rect 12297 9342 12497 9410
rect 12297 9286 12307 9342
rect 12363 9286 12431 9342
rect 12487 9286 12497 9342
rect 12297 9218 12497 9286
rect 12297 9162 12307 9218
rect 12363 9162 12431 9218
rect 12487 9162 12497 9218
rect 12297 9094 12497 9162
rect 12297 9038 12307 9094
rect 12363 9038 12431 9094
rect 12487 9038 12497 9094
rect 12297 8970 12497 9038
rect 12297 8914 12307 8970
rect 12363 8914 12431 8970
rect 12487 8914 12497 8970
rect 12297 8846 12497 8914
rect 12297 8790 12307 8846
rect 12363 8790 12431 8846
rect 12487 8790 12497 8846
rect 12297 8722 12497 8790
rect 12297 8666 12307 8722
rect 12363 8666 12431 8722
rect 12487 8666 12497 8722
rect 12297 8598 12497 8666
rect 12297 8542 12307 8598
rect 12363 8542 12431 8598
rect 12487 8542 12497 8598
rect 12297 8474 12497 8542
rect 12297 8418 12307 8474
rect 12363 8418 12431 8474
rect 12487 8418 12497 8474
rect 12297 8350 12497 8418
rect 12297 8294 12307 8350
rect 12363 8294 12431 8350
rect 12487 8294 12497 8350
rect 12297 8226 12497 8294
rect 12297 8170 12307 8226
rect 12363 8170 12431 8226
rect 12487 8170 12497 8226
rect 12297 8102 12497 8170
rect 12297 8046 12307 8102
rect 12363 8046 12431 8102
rect 12487 8046 12497 8102
rect 12297 8036 12497 8046
rect 2481 7754 2681 7764
rect 2481 7698 2491 7754
rect 2547 7698 2615 7754
rect 2671 7698 2681 7754
rect 2481 7630 2681 7698
rect 2481 7574 2491 7630
rect 2547 7574 2615 7630
rect 2671 7574 2681 7630
rect 2481 7506 2681 7574
rect 2481 7450 2491 7506
rect 2547 7450 2615 7506
rect 2671 7450 2681 7506
rect 2481 7382 2681 7450
rect 2481 7326 2491 7382
rect 2547 7326 2615 7382
rect 2671 7326 2681 7382
rect 2481 7258 2681 7326
rect 2481 7202 2491 7258
rect 2547 7202 2615 7258
rect 2671 7202 2681 7258
rect 2481 7134 2681 7202
rect 2481 7078 2491 7134
rect 2547 7078 2615 7134
rect 2671 7078 2681 7134
rect 2481 7010 2681 7078
rect 2481 6954 2491 7010
rect 2547 6954 2615 7010
rect 2671 6954 2681 7010
rect 2481 6886 2681 6954
rect 2481 6830 2491 6886
rect 2547 6830 2615 6886
rect 2671 6830 2681 6886
rect 2481 6762 2681 6830
rect 2481 6706 2491 6762
rect 2547 6706 2615 6762
rect 2671 6706 2681 6762
rect 2481 6638 2681 6706
rect 2481 6582 2491 6638
rect 2547 6582 2615 6638
rect 2671 6582 2681 6638
rect 2481 6514 2681 6582
rect 2481 6458 2491 6514
rect 2547 6458 2615 6514
rect 2671 6458 2681 6514
rect 2481 6390 2681 6458
rect 2481 6334 2491 6390
rect 2547 6334 2615 6390
rect 2671 6334 2681 6390
rect 2481 6266 2681 6334
rect 2481 6210 2491 6266
rect 2547 6210 2615 6266
rect 2671 6210 2681 6266
rect 2481 6142 2681 6210
rect 2481 6086 2491 6142
rect 2547 6086 2615 6142
rect 2671 6086 2681 6142
rect 2481 6018 2681 6086
rect 2481 5962 2491 6018
rect 2547 5962 2615 6018
rect 2671 5962 2681 6018
rect 2481 5894 2681 5962
rect 2481 5838 2491 5894
rect 2547 5838 2615 5894
rect 2671 5838 2681 5894
rect 2481 5770 2681 5838
rect 2481 5714 2491 5770
rect 2547 5714 2615 5770
rect 2671 5714 2681 5770
rect 2481 5646 2681 5714
rect 2481 5590 2491 5646
rect 2547 5590 2615 5646
rect 2671 5590 2681 5646
rect 2481 5522 2681 5590
rect 2481 5466 2491 5522
rect 2547 5466 2615 5522
rect 2671 5466 2681 5522
rect 2481 5398 2681 5466
rect 2481 5342 2491 5398
rect 2547 5342 2615 5398
rect 2671 5342 2681 5398
rect 2481 5274 2681 5342
rect 2481 5218 2491 5274
rect 2547 5218 2615 5274
rect 2671 5218 2681 5274
rect 2481 5150 2681 5218
rect 2481 5094 2491 5150
rect 2547 5094 2615 5150
rect 2671 5094 2681 5150
rect 2481 5026 2681 5094
rect 2481 4970 2491 5026
rect 2547 4970 2615 5026
rect 2671 4970 2681 5026
rect 2481 4902 2681 4970
rect 2481 4846 2491 4902
rect 2547 4846 2615 4902
rect 2671 4846 2681 4902
rect 2481 4836 2681 4846
rect 4851 7754 5051 7764
rect 4851 7698 4861 7754
rect 4917 7698 4985 7754
rect 5041 7698 5051 7754
rect 4851 7630 5051 7698
rect 4851 7574 4861 7630
rect 4917 7574 4985 7630
rect 5041 7574 5051 7630
rect 4851 7506 5051 7574
rect 4851 7450 4861 7506
rect 4917 7450 4985 7506
rect 5041 7450 5051 7506
rect 4851 7382 5051 7450
rect 4851 7326 4861 7382
rect 4917 7326 4985 7382
rect 5041 7326 5051 7382
rect 4851 7258 5051 7326
rect 4851 7202 4861 7258
rect 4917 7202 4985 7258
rect 5041 7202 5051 7258
rect 4851 7134 5051 7202
rect 4851 7078 4861 7134
rect 4917 7078 4985 7134
rect 5041 7078 5051 7134
rect 4851 7010 5051 7078
rect 4851 6954 4861 7010
rect 4917 6954 4985 7010
rect 5041 6954 5051 7010
rect 4851 6886 5051 6954
rect 4851 6830 4861 6886
rect 4917 6830 4985 6886
rect 5041 6830 5051 6886
rect 4851 6762 5051 6830
rect 4851 6706 4861 6762
rect 4917 6706 4985 6762
rect 5041 6706 5051 6762
rect 4851 6638 5051 6706
rect 4851 6582 4861 6638
rect 4917 6582 4985 6638
rect 5041 6582 5051 6638
rect 4851 6514 5051 6582
rect 4851 6458 4861 6514
rect 4917 6458 4985 6514
rect 5041 6458 5051 6514
rect 4851 6390 5051 6458
rect 4851 6334 4861 6390
rect 4917 6334 4985 6390
rect 5041 6334 5051 6390
rect 4851 6266 5051 6334
rect 4851 6210 4861 6266
rect 4917 6210 4985 6266
rect 5041 6210 5051 6266
rect 4851 6142 5051 6210
rect 4851 6086 4861 6142
rect 4917 6086 4985 6142
rect 5041 6086 5051 6142
rect 4851 6018 5051 6086
rect 4851 5962 4861 6018
rect 4917 5962 4985 6018
rect 5041 5962 5051 6018
rect 4851 5894 5051 5962
rect 4851 5838 4861 5894
rect 4917 5838 4985 5894
rect 5041 5838 5051 5894
rect 4851 5770 5051 5838
rect 4851 5714 4861 5770
rect 4917 5714 4985 5770
rect 5041 5714 5051 5770
rect 4851 5646 5051 5714
rect 4851 5590 4861 5646
rect 4917 5590 4985 5646
rect 5041 5590 5051 5646
rect 4851 5522 5051 5590
rect 4851 5466 4861 5522
rect 4917 5466 4985 5522
rect 5041 5466 5051 5522
rect 4851 5398 5051 5466
rect 4851 5342 4861 5398
rect 4917 5342 4985 5398
rect 5041 5342 5051 5398
rect 4851 5274 5051 5342
rect 4851 5218 4861 5274
rect 4917 5218 4985 5274
rect 5041 5218 5051 5274
rect 4851 5150 5051 5218
rect 4851 5094 4861 5150
rect 4917 5094 4985 5150
rect 5041 5094 5051 5150
rect 4851 5026 5051 5094
rect 4851 4970 4861 5026
rect 4917 4970 4985 5026
rect 5041 4970 5051 5026
rect 4851 4902 5051 4970
rect 4851 4846 4861 4902
rect 4917 4846 4985 4902
rect 5041 4846 5051 4902
rect 4851 4836 5051 4846
rect 7265 7754 7713 7764
rect 7265 7698 7275 7754
rect 7331 7698 7399 7754
rect 7455 7698 7523 7754
rect 7579 7698 7647 7754
rect 7703 7698 7713 7754
rect 7265 7630 7713 7698
rect 7265 7574 7275 7630
rect 7331 7574 7399 7630
rect 7455 7574 7523 7630
rect 7579 7574 7647 7630
rect 7703 7574 7713 7630
rect 7265 7506 7713 7574
rect 7265 7450 7275 7506
rect 7331 7450 7399 7506
rect 7455 7450 7523 7506
rect 7579 7450 7647 7506
rect 7703 7450 7713 7506
rect 7265 7382 7713 7450
rect 7265 7326 7275 7382
rect 7331 7326 7399 7382
rect 7455 7326 7523 7382
rect 7579 7326 7647 7382
rect 7703 7326 7713 7382
rect 7265 7258 7713 7326
rect 7265 7202 7275 7258
rect 7331 7202 7399 7258
rect 7455 7202 7523 7258
rect 7579 7202 7647 7258
rect 7703 7202 7713 7258
rect 7265 7134 7713 7202
rect 7265 7078 7275 7134
rect 7331 7078 7399 7134
rect 7455 7078 7523 7134
rect 7579 7078 7647 7134
rect 7703 7078 7713 7134
rect 7265 7010 7713 7078
rect 7265 6954 7275 7010
rect 7331 6954 7399 7010
rect 7455 6954 7523 7010
rect 7579 6954 7647 7010
rect 7703 6954 7713 7010
rect 7265 6886 7713 6954
rect 7265 6830 7275 6886
rect 7331 6830 7399 6886
rect 7455 6830 7523 6886
rect 7579 6830 7647 6886
rect 7703 6830 7713 6886
rect 7265 6762 7713 6830
rect 7265 6706 7275 6762
rect 7331 6706 7399 6762
rect 7455 6706 7523 6762
rect 7579 6706 7647 6762
rect 7703 6706 7713 6762
rect 7265 6638 7713 6706
rect 7265 6582 7275 6638
rect 7331 6582 7399 6638
rect 7455 6582 7523 6638
rect 7579 6582 7647 6638
rect 7703 6582 7713 6638
rect 7265 6514 7713 6582
rect 7265 6458 7275 6514
rect 7331 6458 7399 6514
rect 7455 6458 7523 6514
rect 7579 6458 7647 6514
rect 7703 6458 7713 6514
rect 7265 6390 7713 6458
rect 7265 6334 7275 6390
rect 7331 6334 7399 6390
rect 7455 6334 7523 6390
rect 7579 6334 7647 6390
rect 7703 6334 7713 6390
rect 7265 6266 7713 6334
rect 7265 6210 7275 6266
rect 7331 6210 7399 6266
rect 7455 6210 7523 6266
rect 7579 6210 7647 6266
rect 7703 6210 7713 6266
rect 7265 6142 7713 6210
rect 7265 6086 7275 6142
rect 7331 6086 7399 6142
rect 7455 6086 7523 6142
rect 7579 6086 7647 6142
rect 7703 6086 7713 6142
rect 7265 6018 7713 6086
rect 7265 5962 7275 6018
rect 7331 5962 7399 6018
rect 7455 5962 7523 6018
rect 7579 5962 7647 6018
rect 7703 5962 7713 6018
rect 7265 5894 7713 5962
rect 7265 5838 7275 5894
rect 7331 5838 7399 5894
rect 7455 5838 7523 5894
rect 7579 5838 7647 5894
rect 7703 5838 7713 5894
rect 7265 5770 7713 5838
rect 7265 5714 7275 5770
rect 7331 5714 7399 5770
rect 7455 5714 7523 5770
rect 7579 5714 7647 5770
rect 7703 5714 7713 5770
rect 7265 5646 7713 5714
rect 7265 5590 7275 5646
rect 7331 5590 7399 5646
rect 7455 5590 7523 5646
rect 7579 5590 7647 5646
rect 7703 5590 7713 5646
rect 7265 5522 7713 5590
rect 7265 5466 7275 5522
rect 7331 5466 7399 5522
rect 7455 5466 7523 5522
rect 7579 5466 7647 5522
rect 7703 5466 7713 5522
rect 7265 5398 7713 5466
rect 7265 5342 7275 5398
rect 7331 5342 7399 5398
rect 7455 5342 7523 5398
rect 7579 5342 7647 5398
rect 7703 5342 7713 5398
rect 7265 5274 7713 5342
rect 7265 5218 7275 5274
rect 7331 5218 7399 5274
rect 7455 5218 7523 5274
rect 7579 5218 7647 5274
rect 7703 5218 7713 5274
rect 7265 5150 7713 5218
rect 7265 5094 7275 5150
rect 7331 5094 7399 5150
rect 7455 5094 7523 5150
rect 7579 5094 7647 5150
rect 7703 5094 7713 5150
rect 7265 5026 7713 5094
rect 7265 4970 7275 5026
rect 7331 4970 7399 5026
rect 7455 4970 7523 5026
rect 7579 4970 7647 5026
rect 7703 4970 7713 5026
rect 7265 4902 7713 4970
rect 7265 4846 7275 4902
rect 7331 4846 7399 4902
rect 7455 4846 7523 4902
rect 7579 4846 7647 4902
rect 7703 4846 7713 4902
rect 7265 4836 7713 4846
rect 9927 7754 10127 7764
rect 9927 7698 9937 7754
rect 9993 7698 10061 7754
rect 10117 7698 10127 7754
rect 9927 7630 10127 7698
rect 9927 7574 9937 7630
rect 9993 7574 10061 7630
rect 10117 7574 10127 7630
rect 9927 7506 10127 7574
rect 9927 7450 9937 7506
rect 9993 7450 10061 7506
rect 10117 7450 10127 7506
rect 9927 7382 10127 7450
rect 9927 7326 9937 7382
rect 9993 7326 10061 7382
rect 10117 7326 10127 7382
rect 9927 7258 10127 7326
rect 9927 7202 9937 7258
rect 9993 7202 10061 7258
rect 10117 7202 10127 7258
rect 9927 7134 10127 7202
rect 9927 7078 9937 7134
rect 9993 7078 10061 7134
rect 10117 7078 10127 7134
rect 9927 7010 10127 7078
rect 9927 6954 9937 7010
rect 9993 6954 10061 7010
rect 10117 6954 10127 7010
rect 9927 6886 10127 6954
rect 9927 6830 9937 6886
rect 9993 6830 10061 6886
rect 10117 6830 10127 6886
rect 9927 6762 10127 6830
rect 9927 6706 9937 6762
rect 9993 6706 10061 6762
rect 10117 6706 10127 6762
rect 9927 6638 10127 6706
rect 9927 6582 9937 6638
rect 9993 6582 10061 6638
rect 10117 6582 10127 6638
rect 9927 6514 10127 6582
rect 9927 6458 9937 6514
rect 9993 6458 10061 6514
rect 10117 6458 10127 6514
rect 9927 6390 10127 6458
rect 9927 6334 9937 6390
rect 9993 6334 10061 6390
rect 10117 6334 10127 6390
rect 9927 6266 10127 6334
rect 9927 6210 9937 6266
rect 9993 6210 10061 6266
rect 10117 6210 10127 6266
rect 9927 6142 10127 6210
rect 9927 6086 9937 6142
rect 9993 6086 10061 6142
rect 10117 6086 10127 6142
rect 9927 6018 10127 6086
rect 9927 5962 9937 6018
rect 9993 5962 10061 6018
rect 10117 5962 10127 6018
rect 9927 5894 10127 5962
rect 9927 5838 9937 5894
rect 9993 5838 10061 5894
rect 10117 5838 10127 5894
rect 9927 5770 10127 5838
rect 9927 5714 9937 5770
rect 9993 5714 10061 5770
rect 10117 5714 10127 5770
rect 9927 5646 10127 5714
rect 9927 5590 9937 5646
rect 9993 5590 10061 5646
rect 10117 5590 10127 5646
rect 9927 5522 10127 5590
rect 9927 5466 9937 5522
rect 9993 5466 10061 5522
rect 10117 5466 10127 5522
rect 9927 5398 10127 5466
rect 9927 5342 9937 5398
rect 9993 5342 10061 5398
rect 10117 5342 10127 5398
rect 9927 5274 10127 5342
rect 9927 5218 9937 5274
rect 9993 5218 10061 5274
rect 10117 5218 10127 5274
rect 9927 5150 10127 5218
rect 9927 5094 9937 5150
rect 9993 5094 10061 5150
rect 10117 5094 10127 5150
rect 9927 5026 10127 5094
rect 9927 4970 9937 5026
rect 9993 4970 10061 5026
rect 10117 4970 10127 5026
rect 9927 4902 10127 4970
rect 9927 4846 9937 4902
rect 9993 4846 10061 4902
rect 10117 4846 10127 4902
rect 9927 4836 10127 4846
rect 12297 7754 12497 7764
rect 12297 7698 12307 7754
rect 12363 7698 12431 7754
rect 12487 7698 12497 7754
rect 12297 7630 12497 7698
rect 12297 7574 12307 7630
rect 12363 7574 12431 7630
rect 12487 7574 12497 7630
rect 12297 7506 12497 7574
rect 12297 7450 12307 7506
rect 12363 7450 12431 7506
rect 12487 7450 12497 7506
rect 12297 7382 12497 7450
rect 12297 7326 12307 7382
rect 12363 7326 12431 7382
rect 12487 7326 12497 7382
rect 12297 7258 12497 7326
rect 12297 7202 12307 7258
rect 12363 7202 12431 7258
rect 12487 7202 12497 7258
rect 12297 7134 12497 7202
rect 12297 7078 12307 7134
rect 12363 7078 12431 7134
rect 12487 7078 12497 7134
rect 12297 7010 12497 7078
rect 12297 6954 12307 7010
rect 12363 6954 12431 7010
rect 12487 6954 12497 7010
rect 12297 6886 12497 6954
rect 12297 6830 12307 6886
rect 12363 6830 12431 6886
rect 12487 6830 12497 6886
rect 12297 6762 12497 6830
rect 12297 6706 12307 6762
rect 12363 6706 12431 6762
rect 12487 6706 12497 6762
rect 12297 6638 12497 6706
rect 12297 6582 12307 6638
rect 12363 6582 12431 6638
rect 12487 6582 12497 6638
rect 12297 6514 12497 6582
rect 12297 6458 12307 6514
rect 12363 6458 12431 6514
rect 12487 6458 12497 6514
rect 12297 6390 12497 6458
rect 12297 6334 12307 6390
rect 12363 6334 12431 6390
rect 12487 6334 12497 6390
rect 12297 6266 12497 6334
rect 12297 6210 12307 6266
rect 12363 6210 12431 6266
rect 12487 6210 12497 6266
rect 12297 6142 12497 6210
rect 12297 6086 12307 6142
rect 12363 6086 12431 6142
rect 12487 6086 12497 6142
rect 12297 6018 12497 6086
rect 12297 5962 12307 6018
rect 12363 5962 12431 6018
rect 12487 5962 12497 6018
rect 12297 5894 12497 5962
rect 12297 5838 12307 5894
rect 12363 5838 12431 5894
rect 12487 5838 12497 5894
rect 12297 5770 12497 5838
rect 12297 5714 12307 5770
rect 12363 5714 12431 5770
rect 12487 5714 12497 5770
rect 12297 5646 12497 5714
rect 12297 5590 12307 5646
rect 12363 5590 12431 5646
rect 12487 5590 12497 5646
rect 12297 5522 12497 5590
rect 12297 5466 12307 5522
rect 12363 5466 12431 5522
rect 12487 5466 12497 5522
rect 12297 5398 12497 5466
rect 12297 5342 12307 5398
rect 12363 5342 12431 5398
rect 12487 5342 12497 5398
rect 12297 5274 12497 5342
rect 12297 5218 12307 5274
rect 12363 5218 12431 5274
rect 12487 5218 12497 5274
rect 12297 5150 12497 5218
rect 12297 5094 12307 5150
rect 12363 5094 12431 5150
rect 12487 5094 12497 5150
rect 12297 5026 12497 5094
rect 12297 4970 12307 5026
rect 12363 4970 12431 5026
rect 12487 4970 12497 5026
rect 12297 4902 12497 4970
rect 12297 4846 12307 4902
rect 12363 4846 12431 4902
rect 12487 4846 12497 4902
rect 12297 4836 12497 4846
rect 2481 4554 2681 4564
rect 2481 4498 2491 4554
rect 2547 4498 2615 4554
rect 2671 4498 2681 4554
rect 2481 4430 2681 4498
rect 2481 4374 2491 4430
rect 2547 4374 2615 4430
rect 2671 4374 2681 4430
rect 2481 4306 2681 4374
rect 2481 4250 2491 4306
rect 2547 4250 2615 4306
rect 2671 4250 2681 4306
rect 2481 4182 2681 4250
rect 2481 4126 2491 4182
rect 2547 4126 2615 4182
rect 2671 4126 2681 4182
rect 2481 4058 2681 4126
rect 2481 4002 2491 4058
rect 2547 4002 2615 4058
rect 2671 4002 2681 4058
rect 2481 3934 2681 4002
rect 2481 3878 2491 3934
rect 2547 3878 2615 3934
rect 2671 3878 2681 3934
rect 2481 3810 2681 3878
rect 2481 3754 2491 3810
rect 2547 3754 2615 3810
rect 2671 3754 2681 3810
rect 2481 3686 2681 3754
rect 2481 3630 2491 3686
rect 2547 3630 2615 3686
rect 2671 3630 2681 3686
rect 2481 3562 2681 3630
rect 2481 3506 2491 3562
rect 2547 3506 2615 3562
rect 2671 3506 2681 3562
rect 2481 3438 2681 3506
rect 2481 3382 2491 3438
rect 2547 3382 2615 3438
rect 2671 3382 2681 3438
rect 2481 3314 2681 3382
rect 2481 3258 2491 3314
rect 2547 3258 2615 3314
rect 2671 3258 2681 3314
rect 2481 3190 2681 3258
rect 2481 3134 2491 3190
rect 2547 3134 2615 3190
rect 2671 3134 2681 3190
rect 2481 3066 2681 3134
rect 2481 3010 2491 3066
rect 2547 3010 2615 3066
rect 2671 3010 2681 3066
rect 2481 2942 2681 3010
rect 2481 2886 2491 2942
rect 2547 2886 2615 2942
rect 2671 2886 2681 2942
rect 2481 2818 2681 2886
rect 2481 2762 2491 2818
rect 2547 2762 2615 2818
rect 2671 2762 2681 2818
rect 2481 2694 2681 2762
rect 2481 2638 2491 2694
rect 2547 2638 2615 2694
rect 2671 2638 2681 2694
rect 2481 2570 2681 2638
rect 2481 2514 2491 2570
rect 2547 2514 2615 2570
rect 2671 2514 2681 2570
rect 2481 2446 2681 2514
rect 2481 2390 2491 2446
rect 2547 2390 2615 2446
rect 2671 2390 2681 2446
rect 2481 2322 2681 2390
rect 2481 2266 2491 2322
rect 2547 2266 2615 2322
rect 2671 2266 2681 2322
rect 2481 2198 2681 2266
rect 2481 2142 2491 2198
rect 2547 2142 2615 2198
rect 2671 2142 2681 2198
rect 2481 2074 2681 2142
rect 2481 2018 2491 2074
rect 2547 2018 2615 2074
rect 2671 2018 2681 2074
rect 2481 1950 2681 2018
rect 2481 1894 2491 1950
rect 2547 1894 2615 1950
rect 2671 1894 2681 1950
rect 2481 1826 2681 1894
rect 2481 1770 2491 1826
rect 2547 1770 2615 1826
rect 2671 1770 2681 1826
rect 2481 1702 2681 1770
rect 2481 1646 2491 1702
rect 2547 1646 2615 1702
rect 2671 1646 2681 1702
rect 2481 1636 2681 1646
rect 4851 4554 5051 4564
rect 4851 4498 4861 4554
rect 4917 4498 4985 4554
rect 5041 4498 5051 4554
rect 4851 4430 5051 4498
rect 4851 4374 4861 4430
rect 4917 4374 4985 4430
rect 5041 4374 5051 4430
rect 4851 4306 5051 4374
rect 4851 4250 4861 4306
rect 4917 4250 4985 4306
rect 5041 4250 5051 4306
rect 4851 4182 5051 4250
rect 4851 4126 4861 4182
rect 4917 4126 4985 4182
rect 5041 4126 5051 4182
rect 4851 4058 5051 4126
rect 4851 4002 4861 4058
rect 4917 4002 4985 4058
rect 5041 4002 5051 4058
rect 4851 3934 5051 4002
rect 4851 3878 4861 3934
rect 4917 3878 4985 3934
rect 5041 3878 5051 3934
rect 4851 3810 5051 3878
rect 4851 3754 4861 3810
rect 4917 3754 4985 3810
rect 5041 3754 5051 3810
rect 4851 3686 5051 3754
rect 4851 3630 4861 3686
rect 4917 3630 4985 3686
rect 5041 3630 5051 3686
rect 4851 3562 5051 3630
rect 4851 3506 4861 3562
rect 4917 3506 4985 3562
rect 5041 3506 5051 3562
rect 4851 3438 5051 3506
rect 4851 3382 4861 3438
rect 4917 3382 4985 3438
rect 5041 3382 5051 3438
rect 4851 3314 5051 3382
rect 4851 3258 4861 3314
rect 4917 3258 4985 3314
rect 5041 3258 5051 3314
rect 4851 3190 5051 3258
rect 4851 3134 4861 3190
rect 4917 3134 4985 3190
rect 5041 3134 5051 3190
rect 4851 3066 5051 3134
rect 4851 3010 4861 3066
rect 4917 3010 4985 3066
rect 5041 3010 5051 3066
rect 4851 2942 5051 3010
rect 4851 2886 4861 2942
rect 4917 2886 4985 2942
rect 5041 2886 5051 2942
rect 4851 2818 5051 2886
rect 4851 2762 4861 2818
rect 4917 2762 4985 2818
rect 5041 2762 5051 2818
rect 4851 2694 5051 2762
rect 4851 2638 4861 2694
rect 4917 2638 4985 2694
rect 5041 2638 5051 2694
rect 4851 2570 5051 2638
rect 4851 2514 4861 2570
rect 4917 2514 4985 2570
rect 5041 2514 5051 2570
rect 4851 2446 5051 2514
rect 4851 2390 4861 2446
rect 4917 2390 4985 2446
rect 5041 2390 5051 2446
rect 4851 2322 5051 2390
rect 4851 2266 4861 2322
rect 4917 2266 4985 2322
rect 5041 2266 5051 2322
rect 4851 2198 5051 2266
rect 4851 2142 4861 2198
rect 4917 2142 4985 2198
rect 5041 2142 5051 2198
rect 4851 2074 5051 2142
rect 4851 2018 4861 2074
rect 4917 2018 4985 2074
rect 5041 2018 5051 2074
rect 4851 1950 5051 2018
rect 4851 1894 4861 1950
rect 4917 1894 4985 1950
rect 5041 1894 5051 1950
rect 4851 1826 5051 1894
rect 4851 1770 4861 1826
rect 4917 1770 4985 1826
rect 5041 1770 5051 1826
rect 4851 1702 5051 1770
rect 4851 1646 4861 1702
rect 4917 1646 4985 1702
rect 5041 1646 5051 1702
rect 4851 1636 5051 1646
rect 7265 4554 7713 4564
rect 7265 4498 7275 4554
rect 7331 4498 7399 4554
rect 7455 4498 7523 4554
rect 7579 4498 7647 4554
rect 7703 4498 7713 4554
rect 7265 4430 7713 4498
rect 7265 4374 7275 4430
rect 7331 4374 7399 4430
rect 7455 4374 7523 4430
rect 7579 4374 7647 4430
rect 7703 4374 7713 4430
rect 7265 4306 7713 4374
rect 7265 4250 7275 4306
rect 7331 4250 7399 4306
rect 7455 4250 7523 4306
rect 7579 4250 7647 4306
rect 7703 4250 7713 4306
rect 7265 4182 7713 4250
rect 7265 4126 7275 4182
rect 7331 4126 7399 4182
rect 7455 4126 7523 4182
rect 7579 4126 7647 4182
rect 7703 4126 7713 4182
rect 7265 4058 7713 4126
rect 7265 4002 7275 4058
rect 7331 4002 7399 4058
rect 7455 4002 7523 4058
rect 7579 4002 7647 4058
rect 7703 4002 7713 4058
rect 7265 3934 7713 4002
rect 7265 3878 7275 3934
rect 7331 3878 7399 3934
rect 7455 3878 7523 3934
rect 7579 3878 7647 3934
rect 7703 3878 7713 3934
rect 7265 3810 7713 3878
rect 7265 3754 7275 3810
rect 7331 3754 7399 3810
rect 7455 3754 7523 3810
rect 7579 3754 7647 3810
rect 7703 3754 7713 3810
rect 7265 3686 7713 3754
rect 7265 3630 7275 3686
rect 7331 3630 7399 3686
rect 7455 3630 7523 3686
rect 7579 3630 7647 3686
rect 7703 3630 7713 3686
rect 7265 3562 7713 3630
rect 7265 3506 7275 3562
rect 7331 3506 7399 3562
rect 7455 3506 7523 3562
rect 7579 3506 7647 3562
rect 7703 3506 7713 3562
rect 7265 3438 7713 3506
rect 7265 3382 7275 3438
rect 7331 3382 7399 3438
rect 7455 3382 7523 3438
rect 7579 3382 7647 3438
rect 7703 3382 7713 3438
rect 7265 3314 7713 3382
rect 7265 3258 7275 3314
rect 7331 3258 7399 3314
rect 7455 3258 7523 3314
rect 7579 3258 7647 3314
rect 7703 3258 7713 3314
rect 7265 3190 7713 3258
rect 7265 3134 7275 3190
rect 7331 3134 7399 3190
rect 7455 3134 7523 3190
rect 7579 3134 7647 3190
rect 7703 3134 7713 3190
rect 7265 3066 7713 3134
rect 7265 3010 7275 3066
rect 7331 3010 7399 3066
rect 7455 3010 7523 3066
rect 7579 3010 7647 3066
rect 7703 3010 7713 3066
rect 7265 2942 7713 3010
rect 7265 2886 7275 2942
rect 7331 2886 7399 2942
rect 7455 2886 7523 2942
rect 7579 2886 7647 2942
rect 7703 2886 7713 2942
rect 7265 2818 7713 2886
rect 7265 2762 7275 2818
rect 7331 2762 7399 2818
rect 7455 2762 7523 2818
rect 7579 2762 7647 2818
rect 7703 2762 7713 2818
rect 7265 2694 7713 2762
rect 7265 2638 7275 2694
rect 7331 2638 7399 2694
rect 7455 2638 7523 2694
rect 7579 2638 7647 2694
rect 7703 2638 7713 2694
rect 7265 2570 7713 2638
rect 7265 2514 7275 2570
rect 7331 2514 7399 2570
rect 7455 2514 7523 2570
rect 7579 2514 7647 2570
rect 7703 2514 7713 2570
rect 7265 2446 7713 2514
rect 7265 2390 7275 2446
rect 7331 2390 7399 2446
rect 7455 2390 7523 2446
rect 7579 2390 7647 2446
rect 7703 2390 7713 2446
rect 7265 2322 7713 2390
rect 7265 2266 7275 2322
rect 7331 2266 7399 2322
rect 7455 2266 7523 2322
rect 7579 2266 7647 2322
rect 7703 2266 7713 2322
rect 7265 2198 7713 2266
rect 7265 2142 7275 2198
rect 7331 2142 7399 2198
rect 7455 2142 7523 2198
rect 7579 2142 7647 2198
rect 7703 2142 7713 2198
rect 7265 2074 7713 2142
rect 7265 2018 7275 2074
rect 7331 2018 7399 2074
rect 7455 2018 7523 2074
rect 7579 2018 7647 2074
rect 7703 2018 7713 2074
rect 7265 1950 7713 2018
rect 7265 1894 7275 1950
rect 7331 1894 7399 1950
rect 7455 1894 7523 1950
rect 7579 1894 7647 1950
rect 7703 1894 7713 1950
rect 7265 1826 7713 1894
rect 7265 1770 7275 1826
rect 7331 1770 7399 1826
rect 7455 1770 7523 1826
rect 7579 1770 7647 1826
rect 7703 1770 7713 1826
rect 7265 1702 7713 1770
rect 7265 1646 7275 1702
rect 7331 1646 7399 1702
rect 7455 1646 7523 1702
rect 7579 1646 7647 1702
rect 7703 1646 7713 1702
rect 7265 1636 7713 1646
rect 9927 4554 10127 4564
rect 9927 4498 9937 4554
rect 9993 4498 10061 4554
rect 10117 4498 10127 4554
rect 9927 4430 10127 4498
rect 9927 4374 9937 4430
rect 9993 4374 10061 4430
rect 10117 4374 10127 4430
rect 9927 4306 10127 4374
rect 9927 4250 9937 4306
rect 9993 4250 10061 4306
rect 10117 4250 10127 4306
rect 9927 4182 10127 4250
rect 9927 4126 9937 4182
rect 9993 4126 10061 4182
rect 10117 4126 10127 4182
rect 9927 4058 10127 4126
rect 9927 4002 9937 4058
rect 9993 4002 10061 4058
rect 10117 4002 10127 4058
rect 9927 3934 10127 4002
rect 9927 3878 9937 3934
rect 9993 3878 10061 3934
rect 10117 3878 10127 3934
rect 9927 3810 10127 3878
rect 9927 3754 9937 3810
rect 9993 3754 10061 3810
rect 10117 3754 10127 3810
rect 9927 3686 10127 3754
rect 9927 3630 9937 3686
rect 9993 3630 10061 3686
rect 10117 3630 10127 3686
rect 9927 3562 10127 3630
rect 9927 3506 9937 3562
rect 9993 3506 10061 3562
rect 10117 3506 10127 3562
rect 9927 3438 10127 3506
rect 9927 3382 9937 3438
rect 9993 3382 10061 3438
rect 10117 3382 10127 3438
rect 9927 3314 10127 3382
rect 9927 3258 9937 3314
rect 9993 3258 10061 3314
rect 10117 3258 10127 3314
rect 9927 3190 10127 3258
rect 9927 3134 9937 3190
rect 9993 3134 10061 3190
rect 10117 3134 10127 3190
rect 9927 3066 10127 3134
rect 9927 3010 9937 3066
rect 9993 3010 10061 3066
rect 10117 3010 10127 3066
rect 9927 2942 10127 3010
rect 9927 2886 9937 2942
rect 9993 2886 10061 2942
rect 10117 2886 10127 2942
rect 9927 2818 10127 2886
rect 9927 2762 9937 2818
rect 9993 2762 10061 2818
rect 10117 2762 10127 2818
rect 9927 2694 10127 2762
rect 9927 2638 9937 2694
rect 9993 2638 10061 2694
rect 10117 2638 10127 2694
rect 9927 2570 10127 2638
rect 9927 2514 9937 2570
rect 9993 2514 10061 2570
rect 10117 2514 10127 2570
rect 9927 2446 10127 2514
rect 9927 2390 9937 2446
rect 9993 2390 10061 2446
rect 10117 2390 10127 2446
rect 9927 2322 10127 2390
rect 9927 2266 9937 2322
rect 9993 2266 10061 2322
rect 10117 2266 10127 2322
rect 9927 2198 10127 2266
rect 9927 2142 9937 2198
rect 9993 2142 10061 2198
rect 10117 2142 10127 2198
rect 9927 2074 10127 2142
rect 9927 2018 9937 2074
rect 9993 2018 10061 2074
rect 10117 2018 10127 2074
rect 9927 1950 10127 2018
rect 9927 1894 9937 1950
rect 9993 1894 10061 1950
rect 10117 1894 10127 1950
rect 9927 1826 10127 1894
rect 9927 1770 9937 1826
rect 9993 1770 10061 1826
rect 10117 1770 10127 1826
rect 9927 1702 10127 1770
rect 9927 1646 9937 1702
rect 9993 1646 10061 1702
rect 10117 1646 10127 1702
rect 9927 1636 10127 1646
rect 12297 4554 12497 4564
rect 12297 4498 12307 4554
rect 12363 4498 12431 4554
rect 12487 4498 12497 4554
rect 12297 4430 12497 4498
rect 12297 4374 12307 4430
rect 12363 4374 12431 4430
rect 12487 4374 12497 4430
rect 12297 4306 12497 4374
rect 12297 4250 12307 4306
rect 12363 4250 12431 4306
rect 12487 4250 12497 4306
rect 12297 4182 12497 4250
rect 12297 4126 12307 4182
rect 12363 4126 12431 4182
rect 12487 4126 12497 4182
rect 12297 4058 12497 4126
rect 12297 4002 12307 4058
rect 12363 4002 12431 4058
rect 12487 4002 12497 4058
rect 12297 3934 12497 4002
rect 12297 3878 12307 3934
rect 12363 3878 12431 3934
rect 12487 3878 12497 3934
rect 12297 3810 12497 3878
rect 12297 3754 12307 3810
rect 12363 3754 12431 3810
rect 12487 3754 12497 3810
rect 12297 3686 12497 3754
rect 12297 3630 12307 3686
rect 12363 3630 12431 3686
rect 12487 3630 12497 3686
rect 12297 3562 12497 3630
rect 12297 3506 12307 3562
rect 12363 3506 12431 3562
rect 12487 3506 12497 3562
rect 12297 3438 12497 3506
rect 12297 3382 12307 3438
rect 12363 3382 12431 3438
rect 12487 3382 12497 3438
rect 12297 3314 12497 3382
rect 12297 3258 12307 3314
rect 12363 3258 12431 3314
rect 12487 3258 12497 3314
rect 12297 3190 12497 3258
rect 12297 3134 12307 3190
rect 12363 3134 12431 3190
rect 12487 3134 12497 3190
rect 12297 3066 12497 3134
rect 12297 3010 12307 3066
rect 12363 3010 12431 3066
rect 12487 3010 12497 3066
rect 12297 2942 12497 3010
rect 12297 2886 12307 2942
rect 12363 2886 12431 2942
rect 12487 2886 12497 2942
rect 12297 2818 12497 2886
rect 12297 2762 12307 2818
rect 12363 2762 12431 2818
rect 12487 2762 12497 2818
rect 12297 2694 12497 2762
rect 12297 2638 12307 2694
rect 12363 2638 12431 2694
rect 12487 2638 12497 2694
rect 12297 2570 12497 2638
rect 12297 2514 12307 2570
rect 12363 2514 12431 2570
rect 12487 2514 12497 2570
rect 12297 2446 12497 2514
rect 12297 2390 12307 2446
rect 12363 2390 12431 2446
rect 12487 2390 12497 2446
rect 12297 2322 12497 2390
rect 12297 2266 12307 2322
rect 12363 2266 12431 2322
rect 12487 2266 12497 2322
rect 12297 2198 12497 2266
rect 12297 2142 12307 2198
rect 12363 2142 12431 2198
rect 12487 2142 12497 2198
rect 12297 2074 12497 2142
rect 12297 2018 12307 2074
rect 12363 2018 12431 2074
rect 12487 2018 12497 2074
rect 12297 1950 12497 2018
rect 12297 1894 12307 1950
rect 12363 1894 12431 1950
rect 12487 1894 12497 1950
rect 12297 1826 12497 1894
rect 12297 1770 12307 1826
rect 12363 1770 12431 1826
rect 12487 1770 12497 1826
rect 12297 1702 12497 1770
rect 12297 1646 12307 1702
rect 12363 1646 12431 1702
rect 12487 1646 12497 1702
rect 12297 1636 12497 1646
rect 261 0 2161 1190
rect 2741 0 4791 1190
rect 5111 0 7161 1190
rect 7817 0 9867 1190
rect 10187 0 12237 1190
rect 12817 0 14717 1190
<< via2 >>
rect 315 55692 371 55748
rect 439 55692 495 55748
rect 563 55692 619 55748
rect 687 55692 743 55748
rect 811 55692 867 55748
rect 935 55692 991 55748
rect 1059 55692 1115 55748
rect 1183 55692 1239 55748
rect 1307 55692 1363 55748
rect 1431 55692 1487 55748
rect 1555 55692 1611 55748
rect 1679 55692 1735 55748
rect 1803 55692 1859 55748
rect 1927 55692 1983 55748
rect 2051 55692 2107 55748
rect 315 55568 371 55624
rect 439 55568 495 55624
rect 563 55568 619 55624
rect 687 55568 743 55624
rect 811 55568 867 55624
rect 935 55568 991 55624
rect 1059 55568 1115 55624
rect 1183 55568 1239 55624
rect 1307 55568 1363 55624
rect 1431 55568 1487 55624
rect 1555 55568 1611 55624
rect 1679 55568 1735 55624
rect 1803 55568 1859 55624
rect 1927 55568 1983 55624
rect 2051 55568 2107 55624
rect 315 55444 371 55500
rect 439 55444 495 55500
rect 563 55444 619 55500
rect 687 55444 743 55500
rect 811 55444 867 55500
rect 935 55444 991 55500
rect 1059 55444 1115 55500
rect 1183 55444 1239 55500
rect 1307 55444 1363 55500
rect 1431 55444 1487 55500
rect 1555 55444 1611 55500
rect 1679 55444 1735 55500
rect 1803 55444 1859 55500
rect 1927 55444 1983 55500
rect 2051 55444 2107 55500
rect 315 55320 371 55376
rect 439 55320 495 55376
rect 563 55320 619 55376
rect 687 55320 743 55376
rect 811 55320 867 55376
rect 935 55320 991 55376
rect 1059 55320 1115 55376
rect 1183 55320 1239 55376
rect 1307 55320 1363 55376
rect 1431 55320 1487 55376
rect 1555 55320 1611 55376
rect 1679 55320 1735 55376
rect 1803 55320 1859 55376
rect 1927 55320 1983 55376
rect 2051 55320 2107 55376
rect 315 55196 371 55252
rect 439 55196 495 55252
rect 563 55196 619 55252
rect 687 55196 743 55252
rect 811 55196 867 55252
rect 935 55196 991 55252
rect 1059 55196 1115 55252
rect 1183 55196 1239 55252
rect 1307 55196 1363 55252
rect 1431 55196 1487 55252
rect 1555 55196 1611 55252
rect 1679 55196 1735 55252
rect 1803 55196 1859 55252
rect 1927 55196 1983 55252
rect 2051 55196 2107 55252
rect 315 55072 371 55128
rect 439 55072 495 55128
rect 563 55072 619 55128
rect 687 55072 743 55128
rect 811 55072 867 55128
rect 935 55072 991 55128
rect 1059 55072 1115 55128
rect 1183 55072 1239 55128
rect 1307 55072 1363 55128
rect 1431 55072 1487 55128
rect 1555 55072 1611 55128
rect 1679 55072 1735 55128
rect 1803 55072 1859 55128
rect 1927 55072 1983 55128
rect 2051 55072 2107 55128
rect 315 54948 371 55004
rect 439 54948 495 55004
rect 563 54948 619 55004
rect 687 54948 743 55004
rect 811 54948 867 55004
rect 935 54948 991 55004
rect 1059 54948 1115 55004
rect 1183 54948 1239 55004
rect 1307 54948 1363 55004
rect 1431 54948 1487 55004
rect 1555 54948 1611 55004
rect 1679 54948 1735 55004
rect 1803 54948 1859 55004
rect 1927 54948 1983 55004
rect 2051 54948 2107 55004
rect 315 54824 371 54880
rect 439 54824 495 54880
rect 563 54824 619 54880
rect 687 54824 743 54880
rect 811 54824 867 54880
rect 935 54824 991 54880
rect 1059 54824 1115 54880
rect 1183 54824 1239 54880
rect 1307 54824 1363 54880
rect 1431 54824 1487 54880
rect 1555 54824 1611 54880
rect 1679 54824 1735 54880
rect 1803 54824 1859 54880
rect 1927 54824 1983 54880
rect 2051 54824 2107 54880
rect 315 54700 371 54756
rect 439 54700 495 54756
rect 563 54700 619 54756
rect 687 54700 743 54756
rect 811 54700 867 54756
rect 935 54700 991 54756
rect 1059 54700 1115 54756
rect 1183 54700 1239 54756
rect 1307 54700 1363 54756
rect 1431 54700 1487 54756
rect 1555 54700 1611 54756
rect 1679 54700 1735 54756
rect 1803 54700 1859 54756
rect 1927 54700 1983 54756
rect 2051 54700 2107 54756
rect 315 54576 371 54632
rect 439 54576 495 54632
rect 563 54576 619 54632
rect 687 54576 743 54632
rect 811 54576 867 54632
rect 935 54576 991 54632
rect 1059 54576 1115 54632
rect 1183 54576 1239 54632
rect 1307 54576 1363 54632
rect 1431 54576 1487 54632
rect 1555 54576 1611 54632
rect 1679 54576 1735 54632
rect 1803 54576 1859 54632
rect 1927 54576 1983 54632
rect 2051 54576 2107 54632
rect 315 54452 371 54508
rect 439 54452 495 54508
rect 563 54452 619 54508
rect 687 54452 743 54508
rect 811 54452 867 54508
rect 935 54452 991 54508
rect 1059 54452 1115 54508
rect 1183 54452 1239 54508
rect 1307 54452 1363 54508
rect 1431 54452 1487 54508
rect 1555 54452 1611 54508
rect 1679 54452 1735 54508
rect 1803 54452 1859 54508
rect 1927 54452 1983 54508
rect 2051 54452 2107 54508
rect 20 52574 76 52576
rect 20 52522 22 52574
rect 22 52522 74 52574
rect 74 52522 76 52574
rect 20 52466 76 52522
rect 20 52414 22 52466
rect 22 52414 74 52466
rect 74 52414 76 52466
rect 20 52358 76 52414
rect 20 52306 22 52358
rect 22 52306 74 52358
rect 74 52306 76 52358
rect 20 52250 76 52306
rect 20 52198 22 52250
rect 22 52198 74 52250
rect 74 52198 76 52250
rect 20 52142 76 52198
rect 20 52090 22 52142
rect 22 52090 74 52142
rect 74 52090 76 52142
rect 20 52034 76 52090
rect 20 51982 22 52034
rect 22 51982 74 52034
rect 74 51982 76 52034
rect 20 51926 76 51982
rect 20 51874 22 51926
rect 22 51874 74 51926
rect 74 51874 76 51926
rect 20 51818 76 51874
rect 20 51766 22 51818
rect 22 51766 74 51818
rect 74 51766 76 51818
rect 20 51710 76 51766
rect 20 51658 22 51710
rect 22 51658 74 51710
rect 74 51658 76 51710
rect 20 51602 76 51658
rect 20 51550 22 51602
rect 22 51550 74 51602
rect 74 51550 76 51602
rect 20 51494 76 51550
rect 20 51442 22 51494
rect 22 51442 74 51494
rect 74 51442 76 51494
rect 20 51386 76 51442
rect 20 51334 22 51386
rect 22 51334 74 51386
rect 74 51334 76 51386
rect 20 51278 76 51334
rect 20 51226 22 51278
rect 22 51226 74 51278
rect 74 51226 76 51278
rect 20 51224 76 51226
rect 2491 57169 2547 57225
rect 2615 57169 2671 57225
rect 2491 57056 2501 57101
rect 2501 57056 2547 57101
rect 2615 57056 2661 57101
rect 2661 57056 2671 57101
rect 2491 57045 2547 57056
rect 2615 57045 2671 57056
rect 2491 56921 2547 56977
rect 2615 56921 2671 56977
rect 2491 56797 2547 56853
rect 2615 56797 2671 56853
rect 2491 56673 2547 56729
rect 2615 56673 2671 56729
rect 2491 56549 2547 56605
rect 2615 56549 2671 56605
rect 2491 56425 2547 56481
rect 2615 56425 2671 56481
rect 2491 56301 2547 56357
rect 2615 56301 2671 56357
rect 2491 56177 2547 56233
rect 2615 56177 2671 56233
rect 2491 56053 2547 56109
rect 2615 56053 2671 56109
rect 2491 54092 2547 54148
rect 2615 54092 2671 54148
rect 2491 53968 2547 54024
rect 2615 53968 2671 54024
rect 2491 53844 2547 53900
rect 2615 53844 2671 53900
rect 2491 53720 2547 53776
rect 2615 53720 2671 53776
rect 2491 53596 2547 53652
rect 2615 53596 2671 53652
rect 2491 53484 2547 53528
rect 2615 53484 2671 53528
rect 2491 53472 2501 53484
rect 2501 53472 2547 53484
rect 2615 53472 2661 53484
rect 2661 53472 2671 53484
rect 2491 53376 2547 53404
rect 2615 53376 2671 53404
rect 2491 53348 2501 53376
rect 2501 53348 2547 53376
rect 2615 53348 2661 53376
rect 2661 53348 2671 53376
rect 2491 53268 2547 53280
rect 2615 53268 2671 53280
rect 2491 53224 2501 53268
rect 2501 53224 2547 53268
rect 2615 53224 2661 53268
rect 2661 53224 2671 53268
rect 2491 53100 2547 53156
rect 2615 53100 2671 53156
rect 2491 52976 2547 53032
rect 2615 52976 2671 53032
rect 2491 52852 2547 52908
rect 2615 52852 2671 52908
rect 315 50892 371 50948
rect 439 50892 495 50948
rect 563 50892 619 50948
rect 687 50892 743 50948
rect 811 50892 867 50948
rect 935 50892 991 50948
rect 1059 50892 1115 50948
rect 1183 50892 1239 50948
rect 1307 50892 1363 50948
rect 1431 50892 1487 50948
rect 1555 50892 1611 50948
rect 1679 50892 1735 50948
rect 1803 50892 1859 50948
rect 1927 50892 1983 50948
rect 2051 50892 2107 50948
rect 315 50768 371 50824
rect 439 50768 495 50824
rect 563 50768 619 50824
rect 687 50768 743 50824
rect 811 50768 867 50824
rect 935 50768 991 50824
rect 1059 50768 1115 50824
rect 1183 50768 1239 50824
rect 1307 50768 1363 50824
rect 1431 50768 1487 50824
rect 1555 50768 1611 50824
rect 1679 50768 1735 50824
rect 1803 50768 1859 50824
rect 1927 50768 1983 50824
rect 2051 50768 2107 50824
rect 315 50644 371 50700
rect 439 50644 495 50700
rect 563 50644 619 50700
rect 687 50644 743 50700
rect 811 50644 867 50700
rect 935 50644 991 50700
rect 1059 50644 1115 50700
rect 1183 50644 1239 50700
rect 1307 50644 1363 50700
rect 1431 50644 1487 50700
rect 1555 50644 1611 50700
rect 1679 50644 1735 50700
rect 1803 50644 1859 50700
rect 1927 50644 1983 50700
rect 2051 50644 2107 50700
rect 315 50520 371 50576
rect 439 50520 495 50576
rect 563 50520 619 50576
rect 687 50520 743 50576
rect 811 50520 867 50576
rect 935 50520 991 50576
rect 1059 50520 1115 50576
rect 1183 50520 1239 50576
rect 1307 50520 1363 50576
rect 1431 50520 1487 50576
rect 1555 50520 1611 50576
rect 1679 50520 1735 50576
rect 1803 50520 1859 50576
rect 1927 50520 1983 50576
rect 2051 50520 2107 50576
rect 315 50396 371 50452
rect 439 50396 495 50452
rect 563 50396 619 50452
rect 687 50396 743 50452
rect 811 50396 867 50452
rect 935 50396 991 50452
rect 1059 50396 1115 50452
rect 1183 50396 1239 50452
rect 1307 50396 1363 50452
rect 1431 50396 1487 50452
rect 1555 50396 1611 50452
rect 1679 50396 1735 50452
rect 1803 50396 1859 50452
rect 1927 50396 1983 50452
rect 2051 50396 2107 50452
rect 315 50272 371 50328
rect 439 50272 495 50328
rect 563 50272 619 50328
rect 687 50272 743 50328
rect 811 50272 867 50328
rect 935 50272 991 50328
rect 1059 50272 1115 50328
rect 1183 50272 1239 50328
rect 1307 50272 1363 50328
rect 1431 50272 1487 50328
rect 1555 50272 1611 50328
rect 1679 50272 1735 50328
rect 1803 50272 1859 50328
rect 1927 50272 1983 50328
rect 2051 50272 2107 50328
rect 315 50148 371 50204
rect 439 50148 495 50204
rect 563 50148 619 50204
rect 687 50148 743 50204
rect 811 50148 867 50204
rect 935 50148 991 50204
rect 1059 50148 1115 50204
rect 1183 50148 1239 50204
rect 1307 50148 1363 50204
rect 1431 50148 1487 50204
rect 1555 50148 1611 50204
rect 1679 50148 1735 50204
rect 1803 50148 1859 50204
rect 1927 50148 1983 50204
rect 2051 50148 2107 50204
rect 315 50024 371 50080
rect 439 50024 495 50080
rect 563 50024 619 50080
rect 687 50024 743 50080
rect 811 50024 867 50080
rect 935 50024 991 50080
rect 1059 50024 1115 50080
rect 1183 50024 1239 50080
rect 1307 50024 1363 50080
rect 1431 50024 1487 50080
rect 1555 50024 1611 50080
rect 1679 50024 1735 50080
rect 1803 50024 1859 50080
rect 1927 50024 1983 50080
rect 2051 50024 2107 50080
rect 315 49900 371 49956
rect 439 49900 495 49956
rect 563 49900 619 49956
rect 687 49900 743 49956
rect 811 49900 867 49956
rect 935 49900 991 49956
rect 1059 49900 1115 49956
rect 1183 49900 1239 49956
rect 1307 49900 1363 49956
rect 1431 49900 1487 49956
rect 1555 49900 1611 49956
rect 1679 49900 1735 49956
rect 1803 49900 1859 49956
rect 1927 49900 1983 49956
rect 2051 49900 2107 49956
rect 315 49776 371 49832
rect 439 49776 495 49832
rect 563 49776 619 49832
rect 687 49776 743 49832
rect 811 49776 867 49832
rect 935 49776 991 49832
rect 1059 49776 1115 49832
rect 1183 49776 1239 49832
rect 1307 49776 1363 49832
rect 1431 49776 1487 49832
rect 1555 49776 1611 49832
rect 1679 49776 1735 49832
rect 1803 49776 1859 49832
rect 1927 49776 1983 49832
rect 2051 49776 2107 49832
rect 315 49652 371 49708
rect 439 49652 495 49708
rect 563 49652 619 49708
rect 687 49652 743 49708
rect 811 49652 867 49708
rect 935 49652 991 49708
rect 1059 49652 1115 49708
rect 1183 49652 1239 49708
rect 1307 49652 1363 49708
rect 1431 49652 1487 49708
rect 1555 49652 1611 49708
rect 1679 49652 1735 49708
rect 1803 49652 1859 49708
rect 1927 49652 1983 49708
rect 2051 49652 2107 49708
rect 315 47692 371 47748
rect 439 47692 495 47748
rect 563 47692 619 47748
rect 687 47692 743 47748
rect 811 47692 867 47748
rect 935 47692 991 47748
rect 1059 47692 1115 47748
rect 1183 47692 1239 47748
rect 1307 47692 1363 47748
rect 1431 47692 1487 47748
rect 1555 47692 1611 47748
rect 1679 47692 1735 47748
rect 1803 47692 1859 47748
rect 1927 47692 1983 47748
rect 2051 47692 2107 47748
rect 315 47568 371 47624
rect 439 47568 495 47624
rect 563 47568 619 47624
rect 687 47568 743 47624
rect 811 47568 867 47624
rect 935 47568 991 47624
rect 1059 47568 1115 47624
rect 1183 47568 1239 47624
rect 1307 47568 1363 47624
rect 1431 47568 1487 47624
rect 1555 47568 1611 47624
rect 1679 47568 1735 47624
rect 1803 47568 1859 47624
rect 1927 47568 1983 47624
rect 2051 47568 2107 47624
rect 315 47444 371 47500
rect 439 47444 495 47500
rect 563 47444 619 47500
rect 687 47444 743 47500
rect 811 47444 867 47500
rect 935 47444 991 47500
rect 1059 47444 1115 47500
rect 1183 47444 1239 47500
rect 1307 47444 1363 47500
rect 1431 47444 1487 47500
rect 1555 47444 1611 47500
rect 1679 47444 1735 47500
rect 1803 47444 1859 47500
rect 1927 47444 1983 47500
rect 2051 47444 2107 47500
rect 315 47320 371 47376
rect 439 47320 495 47376
rect 563 47320 619 47376
rect 687 47320 743 47376
rect 811 47320 867 47376
rect 935 47320 991 47376
rect 1059 47320 1115 47376
rect 1183 47320 1239 47376
rect 1307 47320 1363 47376
rect 1431 47320 1487 47376
rect 1555 47320 1611 47376
rect 1679 47320 1735 47376
rect 1803 47320 1859 47376
rect 1927 47320 1983 47376
rect 2051 47320 2107 47376
rect 2289 52465 2345 52521
rect 2289 52333 2345 52389
rect 2289 52201 2345 52257
rect 2289 52069 2345 52125
rect 2289 51937 2345 51993
rect 2289 51805 2345 51861
rect 2289 51673 2345 51729
rect 2289 51541 2345 51597
rect 2289 51409 2345 51465
rect 2289 51277 2345 51333
rect 315 47196 371 47252
rect 439 47196 495 47252
rect 563 47196 619 47252
rect 687 47196 743 47252
rect 811 47196 867 47252
rect 935 47196 991 47252
rect 1059 47196 1115 47252
rect 1183 47196 1239 47252
rect 1307 47196 1363 47252
rect 1431 47196 1487 47252
rect 1555 47196 1611 47252
rect 1679 47196 1735 47252
rect 1803 47196 1859 47252
rect 1927 47196 1983 47252
rect 2051 47196 2107 47252
rect 315 47072 371 47128
rect 439 47072 495 47128
rect 563 47072 619 47128
rect 687 47072 743 47128
rect 811 47072 867 47128
rect 935 47072 991 47128
rect 1059 47072 1115 47128
rect 1183 47072 1239 47128
rect 1307 47072 1363 47128
rect 1431 47072 1487 47128
rect 1555 47072 1611 47128
rect 1679 47072 1735 47128
rect 1803 47072 1859 47128
rect 1927 47072 1983 47128
rect 2051 47072 2107 47128
rect 315 46948 371 47004
rect 439 46948 495 47004
rect 563 46948 619 47004
rect 687 46948 743 47004
rect 811 46948 867 47004
rect 935 46948 991 47004
rect 1059 46948 1115 47004
rect 1183 46948 1239 47004
rect 1307 46948 1363 47004
rect 1431 46948 1487 47004
rect 1555 46948 1611 47004
rect 1679 46948 1735 47004
rect 1803 46948 1859 47004
rect 1927 46948 1983 47004
rect 2051 46948 2107 47004
rect 315 46824 371 46880
rect 439 46824 495 46880
rect 563 46824 619 46880
rect 687 46824 743 46880
rect 811 46824 867 46880
rect 935 46824 991 46880
rect 1059 46824 1115 46880
rect 1183 46824 1239 46880
rect 1307 46824 1363 46880
rect 1431 46824 1487 46880
rect 1555 46824 1611 46880
rect 1679 46824 1735 46880
rect 1803 46824 1859 46880
rect 1927 46824 1983 46880
rect 2051 46824 2107 46880
rect 315 46700 371 46756
rect 439 46700 495 46756
rect 563 46700 619 46756
rect 687 46700 743 46756
rect 811 46700 867 46756
rect 935 46700 991 46756
rect 1059 46700 1115 46756
rect 1183 46700 1239 46756
rect 1307 46700 1363 46756
rect 1431 46700 1487 46756
rect 1555 46700 1611 46756
rect 1679 46700 1735 46756
rect 1803 46700 1859 46756
rect 1927 46700 1983 46756
rect 2051 46700 2107 46756
rect 315 46576 371 46632
rect 439 46576 495 46632
rect 563 46576 619 46632
rect 687 46576 743 46632
rect 811 46576 867 46632
rect 935 46576 991 46632
rect 1059 46576 1115 46632
rect 1183 46576 1239 46632
rect 1307 46576 1363 46632
rect 1431 46576 1487 46632
rect 1555 46576 1611 46632
rect 1679 46576 1735 46632
rect 1803 46576 1859 46632
rect 1927 46576 1983 46632
rect 2051 46576 2107 46632
rect 315 46452 371 46508
rect 439 46452 495 46508
rect 563 46452 619 46508
rect 687 46452 743 46508
rect 811 46452 867 46508
rect 935 46452 991 46508
rect 1059 46452 1115 46508
rect 1183 46452 1239 46508
rect 1307 46452 1363 46508
rect 1431 46452 1487 46508
rect 1555 46452 1611 46508
rect 1679 46452 1735 46508
rect 1803 46452 1859 46508
rect 1927 46452 1983 46508
rect 2051 46452 2107 46508
rect 315 44492 371 44548
rect 439 44492 495 44548
rect 563 44492 619 44548
rect 687 44492 743 44548
rect 811 44492 867 44548
rect 935 44492 991 44548
rect 1059 44492 1115 44548
rect 1183 44492 1239 44548
rect 1307 44492 1363 44548
rect 1431 44492 1487 44548
rect 1555 44492 1611 44548
rect 1679 44492 1735 44548
rect 1803 44492 1859 44548
rect 1927 44492 1983 44548
rect 2051 44492 2107 44548
rect 315 44368 371 44424
rect 439 44368 495 44424
rect 563 44368 619 44424
rect 687 44368 743 44424
rect 811 44368 867 44424
rect 935 44368 991 44424
rect 1059 44368 1115 44424
rect 1183 44368 1239 44424
rect 1307 44368 1363 44424
rect 1431 44368 1487 44424
rect 1555 44368 1611 44424
rect 1679 44368 1735 44424
rect 1803 44368 1859 44424
rect 1927 44368 1983 44424
rect 2051 44368 2107 44424
rect 315 44244 371 44300
rect 439 44244 495 44300
rect 563 44244 619 44300
rect 687 44244 743 44300
rect 811 44244 867 44300
rect 935 44244 991 44300
rect 1059 44244 1115 44300
rect 1183 44244 1239 44300
rect 1307 44244 1363 44300
rect 1431 44244 1487 44300
rect 1555 44244 1611 44300
rect 1679 44244 1735 44300
rect 1803 44244 1859 44300
rect 1927 44244 1983 44300
rect 2051 44244 2107 44300
rect 315 44120 371 44176
rect 439 44120 495 44176
rect 563 44120 619 44176
rect 687 44120 743 44176
rect 811 44120 867 44176
rect 935 44120 991 44176
rect 1059 44120 1115 44176
rect 1183 44120 1239 44176
rect 1307 44120 1363 44176
rect 1431 44120 1487 44176
rect 1555 44120 1611 44176
rect 1679 44120 1735 44176
rect 1803 44120 1859 44176
rect 1927 44120 1983 44176
rect 2051 44120 2107 44176
rect 315 43996 371 44052
rect 439 43996 495 44052
rect 563 43996 619 44052
rect 687 43996 743 44052
rect 811 43996 867 44052
rect 935 43996 991 44052
rect 1059 43996 1115 44052
rect 1183 43996 1239 44052
rect 1307 43996 1363 44052
rect 1431 43996 1487 44052
rect 1555 43996 1611 44052
rect 1679 43996 1735 44052
rect 1803 43996 1859 44052
rect 1927 43996 1983 44052
rect 2051 43996 2107 44052
rect 315 43872 371 43928
rect 439 43872 495 43928
rect 563 43872 619 43928
rect 687 43872 743 43928
rect 811 43872 867 43928
rect 935 43872 991 43928
rect 1059 43872 1115 43928
rect 1183 43872 1239 43928
rect 1307 43872 1363 43928
rect 1431 43872 1487 43928
rect 1555 43872 1611 43928
rect 1679 43872 1735 43928
rect 1803 43872 1859 43928
rect 1927 43872 1983 43928
rect 2051 43872 2107 43928
rect 315 43748 371 43804
rect 439 43748 495 43804
rect 563 43748 619 43804
rect 687 43748 743 43804
rect 811 43748 867 43804
rect 935 43748 991 43804
rect 1059 43748 1115 43804
rect 1183 43748 1239 43804
rect 1307 43748 1363 43804
rect 1431 43748 1487 43804
rect 1555 43748 1611 43804
rect 1679 43748 1735 43804
rect 1803 43748 1859 43804
rect 1927 43748 1983 43804
rect 2051 43748 2107 43804
rect 315 43624 371 43680
rect 439 43624 495 43680
rect 563 43624 619 43680
rect 687 43624 743 43680
rect 811 43624 867 43680
rect 935 43624 991 43680
rect 1059 43624 1115 43680
rect 1183 43624 1239 43680
rect 1307 43624 1363 43680
rect 1431 43624 1487 43680
rect 1555 43624 1611 43680
rect 1679 43624 1735 43680
rect 1803 43624 1859 43680
rect 1927 43624 1983 43680
rect 2051 43624 2107 43680
rect 315 43500 371 43556
rect 439 43500 495 43556
rect 563 43500 619 43556
rect 687 43500 743 43556
rect 811 43500 867 43556
rect 935 43500 991 43556
rect 1059 43500 1115 43556
rect 1183 43500 1239 43556
rect 1307 43500 1363 43556
rect 1431 43500 1487 43556
rect 1555 43500 1611 43556
rect 1679 43500 1735 43556
rect 1803 43500 1859 43556
rect 1927 43500 1983 43556
rect 2051 43500 2107 43556
rect 315 43376 371 43432
rect 439 43376 495 43432
rect 563 43376 619 43432
rect 687 43376 743 43432
rect 811 43376 867 43432
rect 935 43376 991 43432
rect 1059 43376 1115 43432
rect 1183 43376 1239 43432
rect 1307 43376 1363 43432
rect 1431 43376 1487 43432
rect 1555 43376 1611 43432
rect 1679 43376 1735 43432
rect 1803 43376 1859 43432
rect 1927 43376 1983 43432
rect 2051 43376 2107 43432
rect 315 43252 371 43308
rect 439 43252 495 43308
rect 563 43252 619 43308
rect 687 43252 743 43308
rect 811 43252 867 43308
rect 935 43252 991 43308
rect 1059 43252 1115 43308
rect 1183 43252 1239 43308
rect 1307 43252 1363 43308
rect 1431 43252 1487 43308
rect 1555 43252 1611 43308
rect 1679 43252 1735 43308
rect 1803 43252 1859 43308
rect 1927 43252 1983 43308
rect 2051 43252 2107 43308
rect 315 42892 371 42948
rect 439 42892 495 42948
rect 563 42892 619 42948
rect 687 42892 743 42948
rect 811 42892 867 42948
rect 935 42892 991 42948
rect 1059 42892 1115 42948
rect 1183 42892 1239 42948
rect 1307 42892 1363 42948
rect 1431 42892 1487 42948
rect 1555 42892 1611 42948
rect 1679 42892 1735 42948
rect 1803 42892 1859 42948
rect 1927 42892 1983 42948
rect 2051 42892 2107 42948
rect 315 42768 371 42824
rect 439 42768 495 42824
rect 563 42768 619 42824
rect 687 42768 743 42824
rect 811 42768 867 42824
rect 935 42768 991 42824
rect 1059 42768 1115 42824
rect 1183 42768 1239 42824
rect 1307 42768 1363 42824
rect 1431 42768 1487 42824
rect 1555 42768 1611 42824
rect 1679 42768 1735 42824
rect 1803 42768 1859 42824
rect 1927 42768 1983 42824
rect 2051 42768 2107 42824
rect 315 42644 371 42700
rect 439 42644 495 42700
rect 563 42644 619 42700
rect 687 42644 743 42700
rect 811 42644 867 42700
rect 935 42644 991 42700
rect 1059 42644 1115 42700
rect 1183 42644 1239 42700
rect 1307 42644 1363 42700
rect 1431 42644 1487 42700
rect 1555 42644 1611 42700
rect 1679 42644 1735 42700
rect 1803 42644 1859 42700
rect 1927 42644 1983 42700
rect 2051 42644 2107 42700
rect 315 42520 371 42576
rect 439 42520 495 42576
rect 563 42520 619 42576
rect 687 42520 743 42576
rect 811 42520 867 42576
rect 935 42520 991 42576
rect 1059 42520 1115 42576
rect 1183 42520 1239 42576
rect 1307 42520 1363 42576
rect 1431 42520 1487 42576
rect 1555 42520 1611 42576
rect 1679 42520 1735 42576
rect 1803 42520 1859 42576
rect 1927 42520 1983 42576
rect 2051 42520 2107 42576
rect 315 42396 371 42452
rect 439 42396 495 42452
rect 563 42396 619 42452
rect 687 42396 743 42452
rect 811 42396 867 42452
rect 935 42396 991 42452
rect 1059 42396 1115 42452
rect 1183 42396 1239 42452
rect 1307 42396 1363 42452
rect 1431 42396 1487 42452
rect 1555 42396 1611 42452
rect 1679 42396 1735 42452
rect 1803 42396 1859 42452
rect 1927 42396 1983 42452
rect 2051 42396 2107 42452
rect 315 42272 371 42328
rect 439 42272 495 42328
rect 563 42272 619 42328
rect 687 42272 743 42328
rect 811 42272 867 42328
rect 935 42272 991 42328
rect 1059 42272 1115 42328
rect 1183 42272 1239 42328
rect 1307 42272 1363 42328
rect 1431 42272 1487 42328
rect 1555 42272 1611 42328
rect 1679 42272 1735 42328
rect 1803 42272 1859 42328
rect 1927 42272 1983 42328
rect 2051 42272 2107 42328
rect 315 42148 371 42204
rect 439 42148 495 42204
rect 563 42148 619 42204
rect 687 42148 743 42204
rect 811 42148 867 42204
rect 935 42148 991 42204
rect 1059 42148 1115 42204
rect 1183 42148 1239 42204
rect 1307 42148 1363 42204
rect 1431 42148 1487 42204
rect 1555 42148 1611 42204
rect 1679 42148 1735 42204
rect 1803 42148 1859 42204
rect 1927 42148 1983 42204
rect 2051 42148 2107 42204
rect 315 42024 371 42080
rect 439 42024 495 42080
rect 563 42024 619 42080
rect 687 42024 743 42080
rect 811 42024 867 42080
rect 935 42024 991 42080
rect 1059 42024 1115 42080
rect 1183 42024 1239 42080
rect 1307 42024 1363 42080
rect 1431 42024 1487 42080
rect 1555 42024 1611 42080
rect 1679 42024 1735 42080
rect 1803 42024 1859 42080
rect 1927 42024 1983 42080
rect 2051 42024 2107 42080
rect 315 41900 371 41956
rect 439 41900 495 41956
rect 563 41900 619 41956
rect 687 41900 743 41956
rect 811 41900 867 41956
rect 935 41900 991 41956
rect 1059 41900 1115 41956
rect 1183 41900 1239 41956
rect 1307 41900 1363 41956
rect 1431 41900 1487 41956
rect 1555 41900 1611 41956
rect 1679 41900 1735 41956
rect 1803 41900 1859 41956
rect 1927 41900 1983 41956
rect 2051 41900 2107 41956
rect 315 41776 371 41832
rect 439 41776 495 41832
rect 563 41776 619 41832
rect 687 41776 743 41832
rect 811 41776 867 41832
rect 935 41776 991 41832
rect 1059 41776 1115 41832
rect 1183 41776 1239 41832
rect 1307 41776 1363 41832
rect 1431 41776 1487 41832
rect 1555 41776 1611 41832
rect 1679 41776 1735 41832
rect 1803 41776 1859 41832
rect 1927 41776 1983 41832
rect 2051 41776 2107 41832
rect 315 41652 371 41708
rect 439 41652 495 41708
rect 563 41652 619 41708
rect 687 41652 743 41708
rect 811 41652 867 41708
rect 935 41652 991 41708
rect 1059 41652 1115 41708
rect 1183 41652 1239 41708
rect 1307 41652 1363 41708
rect 1431 41652 1487 41708
rect 1555 41652 1611 41708
rect 1679 41652 1735 41708
rect 1803 41652 1859 41708
rect 1927 41652 1983 41708
rect 2051 41652 2107 41708
rect 315 41292 371 41348
rect 439 41292 495 41348
rect 563 41292 619 41348
rect 687 41292 743 41348
rect 811 41292 867 41348
rect 935 41292 991 41348
rect 1059 41292 1115 41348
rect 1183 41292 1239 41348
rect 1307 41292 1363 41348
rect 1431 41292 1487 41348
rect 1555 41292 1611 41348
rect 1679 41292 1735 41348
rect 1803 41292 1859 41348
rect 1927 41292 1983 41348
rect 2051 41292 2107 41348
rect 315 41168 371 41224
rect 439 41168 495 41224
rect 563 41168 619 41224
rect 687 41168 743 41224
rect 811 41168 867 41224
rect 935 41168 991 41224
rect 1059 41168 1115 41224
rect 1183 41168 1239 41224
rect 1307 41168 1363 41224
rect 1431 41168 1487 41224
rect 1555 41168 1611 41224
rect 1679 41168 1735 41224
rect 1803 41168 1859 41224
rect 1927 41168 1983 41224
rect 2051 41168 2107 41224
rect 315 41044 371 41100
rect 439 41044 495 41100
rect 563 41044 619 41100
rect 687 41044 743 41100
rect 811 41044 867 41100
rect 935 41044 991 41100
rect 1059 41044 1115 41100
rect 1183 41044 1239 41100
rect 1307 41044 1363 41100
rect 1431 41044 1487 41100
rect 1555 41044 1611 41100
rect 1679 41044 1735 41100
rect 1803 41044 1859 41100
rect 1927 41044 1983 41100
rect 2051 41044 2107 41100
rect 315 40920 371 40976
rect 439 40920 495 40976
rect 563 40920 619 40976
rect 687 40920 743 40976
rect 811 40920 867 40976
rect 935 40920 991 40976
rect 1059 40920 1115 40976
rect 1183 40920 1239 40976
rect 1307 40920 1363 40976
rect 1431 40920 1487 40976
rect 1555 40920 1611 40976
rect 1679 40920 1735 40976
rect 1803 40920 1859 40976
rect 1927 40920 1983 40976
rect 2051 40920 2107 40976
rect 315 40796 371 40852
rect 439 40796 495 40852
rect 563 40796 619 40852
rect 687 40796 743 40852
rect 811 40796 867 40852
rect 935 40796 991 40852
rect 1059 40796 1115 40852
rect 1183 40796 1239 40852
rect 1307 40796 1363 40852
rect 1431 40796 1487 40852
rect 1555 40796 1611 40852
rect 1679 40796 1735 40852
rect 1803 40796 1859 40852
rect 1927 40796 1983 40852
rect 2051 40796 2107 40852
rect 315 40672 371 40728
rect 439 40672 495 40728
rect 563 40672 619 40728
rect 687 40672 743 40728
rect 811 40672 867 40728
rect 935 40672 991 40728
rect 1059 40672 1115 40728
rect 1183 40672 1239 40728
rect 1307 40672 1363 40728
rect 1431 40672 1487 40728
rect 1555 40672 1611 40728
rect 1679 40672 1735 40728
rect 1803 40672 1859 40728
rect 1927 40672 1983 40728
rect 2051 40672 2107 40728
rect 315 40548 371 40604
rect 439 40548 495 40604
rect 563 40548 619 40604
rect 687 40548 743 40604
rect 811 40548 867 40604
rect 935 40548 991 40604
rect 1059 40548 1115 40604
rect 1183 40548 1239 40604
rect 1307 40548 1363 40604
rect 1431 40548 1487 40604
rect 1555 40548 1611 40604
rect 1679 40548 1735 40604
rect 1803 40548 1859 40604
rect 1927 40548 1983 40604
rect 2051 40548 2107 40604
rect 315 40424 371 40480
rect 439 40424 495 40480
rect 563 40424 619 40480
rect 687 40424 743 40480
rect 811 40424 867 40480
rect 935 40424 991 40480
rect 1059 40424 1115 40480
rect 1183 40424 1239 40480
rect 1307 40424 1363 40480
rect 1431 40424 1487 40480
rect 1555 40424 1611 40480
rect 1679 40424 1735 40480
rect 1803 40424 1859 40480
rect 1927 40424 1983 40480
rect 2051 40424 2107 40480
rect 315 40300 371 40356
rect 439 40300 495 40356
rect 563 40300 619 40356
rect 687 40300 743 40356
rect 811 40300 867 40356
rect 935 40300 991 40356
rect 1059 40300 1115 40356
rect 1183 40300 1239 40356
rect 1307 40300 1363 40356
rect 1431 40300 1487 40356
rect 1555 40300 1611 40356
rect 1679 40300 1735 40356
rect 1803 40300 1859 40356
rect 1927 40300 1983 40356
rect 2051 40300 2107 40356
rect 315 40176 371 40232
rect 439 40176 495 40232
rect 563 40176 619 40232
rect 687 40176 743 40232
rect 811 40176 867 40232
rect 935 40176 991 40232
rect 1059 40176 1115 40232
rect 1183 40176 1239 40232
rect 1307 40176 1363 40232
rect 1431 40176 1487 40232
rect 1555 40176 1611 40232
rect 1679 40176 1735 40232
rect 1803 40176 1859 40232
rect 1927 40176 1983 40232
rect 2051 40176 2107 40232
rect 315 40052 371 40108
rect 439 40052 495 40108
rect 563 40052 619 40108
rect 687 40052 743 40108
rect 811 40052 867 40108
rect 935 40052 991 40108
rect 1059 40052 1115 40108
rect 1183 40052 1239 40108
rect 1307 40052 1363 40108
rect 1431 40052 1487 40108
rect 1555 40052 1611 40108
rect 1679 40052 1735 40108
rect 1803 40052 1859 40108
rect 1927 40052 1983 40108
rect 2051 40052 2107 40108
rect 315 39692 371 39748
rect 439 39692 495 39748
rect 563 39692 619 39748
rect 687 39692 743 39748
rect 811 39692 867 39748
rect 935 39692 991 39748
rect 1059 39692 1115 39748
rect 1183 39692 1239 39748
rect 1307 39692 1363 39748
rect 1431 39692 1487 39748
rect 1555 39692 1611 39748
rect 1679 39692 1735 39748
rect 1803 39692 1859 39748
rect 1927 39692 1983 39748
rect 2051 39692 2107 39748
rect 315 39568 371 39624
rect 439 39568 495 39624
rect 563 39568 619 39624
rect 687 39568 743 39624
rect 811 39568 867 39624
rect 935 39568 991 39624
rect 1059 39568 1115 39624
rect 1183 39568 1239 39624
rect 1307 39568 1363 39624
rect 1431 39568 1487 39624
rect 1555 39568 1611 39624
rect 1679 39568 1735 39624
rect 1803 39568 1859 39624
rect 1927 39568 1983 39624
rect 2051 39568 2107 39624
rect 315 39444 371 39500
rect 439 39444 495 39500
rect 563 39444 619 39500
rect 687 39444 743 39500
rect 811 39444 867 39500
rect 935 39444 991 39500
rect 1059 39444 1115 39500
rect 1183 39444 1239 39500
rect 1307 39444 1363 39500
rect 1431 39444 1487 39500
rect 1555 39444 1611 39500
rect 1679 39444 1735 39500
rect 1803 39444 1859 39500
rect 1927 39444 1983 39500
rect 2051 39444 2107 39500
rect 315 39320 371 39376
rect 439 39320 495 39376
rect 563 39320 619 39376
rect 687 39320 743 39376
rect 811 39320 867 39376
rect 935 39320 991 39376
rect 1059 39320 1115 39376
rect 1183 39320 1239 39376
rect 1307 39320 1363 39376
rect 1431 39320 1487 39376
rect 1555 39320 1611 39376
rect 1679 39320 1735 39376
rect 1803 39320 1859 39376
rect 1927 39320 1983 39376
rect 2051 39320 2107 39376
rect 315 39196 371 39252
rect 439 39196 495 39252
rect 563 39196 619 39252
rect 687 39196 743 39252
rect 811 39196 867 39252
rect 935 39196 991 39252
rect 1059 39196 1115 39252
rect 1183 39196 1239 39252
rect 1307 39196 1363 39252
rect 1431 39196 1487 39252
rect 1555 39196 1611 39252
rect 1679 39196 1735 39252
rect 1803 39196 1859 39252
rect 1927 39196 1983 39252
rect 2051 39196 2107 39252
rect 315 39072 371 39128
rect 439 39072 495 39128
rect 563 39072 619 39128
rect 687 39072 743 39128
rect 811 39072 867 39128
rect 935 39072 991 39128
rect 1059 39072 1115 39128
rect 1183 39072 1239 39128
rect 1307 39072 1363 39128
rect 1431 39072 1487 39128
rect 1555 39072 1611 39128
rect 1679 39072 1735 39128
rect 1803 39072 1859 39128
rect 1927 39072 1983 39128
rect 2051 39072 2107 39128
rect 315 38948 371 39004
rect 439 38948 495 39004
rect 563 38948 619 39004
rect 687 38948 743 39004
rect 811 38948 867 39004
rect 935 38948 991 39004
rect 1059 38948 1115 39004
rect 1183 38948 1239 39004
rect 1307 38948 1363 39004
rect 1431 38948 1487 39004
rect 1555 38948 1611 39004
rect 1679 38948 1735 39004
rect 1803 38948 1859 39004
rect 1927 38948 1983 39004
rect 2051 38948 2107 39004
rect 315 38824 371 38880
rect 439 38824 495 38880
rect 563 38824 619 38880
rect 687 38824 743 38880
rect 811 38824 867 38880
rect 935 38824 991 38880
rect 1059 38824 1115 38880
rect 1183 38824 1239 38880
rect 1307 38824 1363 38880
rect 1431 38824 1487 38880
rect 1555 38824 1611 38880
rect 1679 38824 1735 38880
rect 1803 38824 1859 38880
rect 1927 38824 1983 38880
rect 2051 38824 2107 38880
rect 315 38700 371 38756
rect 439 38700 495 38756
rect 563 38700 619 38756
rect 687 38700 743 38756
rect 811 38700 867 38756
rect 935 38700 991 38756
rect 1059 38700 1115 38756
rect 1183 38700 1239 38756
rect 1307 38700 1363 38756
rect 1431 38700 1487 38756
rect 1555 38700 1611 38756
rect 1679 38700 1735 38756
rect 1803 38700 1859 38756
rect 1927 38700 1983 38756
rect 2051 38700 2107 38756
rect 315 38576 371 38632
rect 439 38576 495 38632
rect 563 38576 619 38632
rect 687 38576 743 38632
rect 811 38576 867 38632
rect 935 38576 991 38632
rect 1059 38576 1115 38632
rect 1183 38576 1239 38632
rect 1307 38576 1363 38632
rect 1431 38576 1487 38632
rect 1555 38576 1611 38632
rect 1679 38576 1735 38632
rect 1803 38576 1859 38632
rect 1927 38576 1983 38632
rect 2051 38576 2107 38632
rect 315 38452 371 38508
rect 439 38452 495 38508
rect 563 38452 619 38508
rect 687 38452 743 38508
rect 811 38452 867 38508
rect 935 38452 991 38508
rect 1059 38452 1115 38508
rect 1183 38452 1239 38508
rect 1307 38452 1363 38508
rect 1431 38452 1487 38508
rect 1555 38452 1611 38508
rect 1679 38452 1735 38508
rect 1803 38452 1859 38508
rect 1927 38452 1983 38508
rect 2051 38452 2107 38508
rect 20 38174 76 38176
rect 20 38122 22 38174
rect 22 38122 74 38174
rect 74 38122 76 38174
rect 20 38066 76 38122
rect 20 38014 22 38066
rect 22 38014 74 38066
rect 74 38014 76 38066
rect 20 37958 76 38014
rect 20 37906 22 37958
rect 22 37906 74 37958
rect 74 37906 76 37958
rect 20 37850 76 37906
rect 20 37798 22 37850
rect 22 37798 74 37850
rect 74 37798 76 37850
rect 20 37742 76 37798
rect 20 37690 22 37742
rect 22 37690 74 37742
rect 74 37690 76 37742
rect 20 37634 76 37690
rect 20 37582 22 37634
rect 22 37582 74 37634
rect 74 37582 76 37634
rect 20 37526 76 37582
rect 20 37474 22 37526
rect 22 37474 74 37526
rect 74 37474 76 37526
rect 20 37418 76 37474
rect 20 37366 22 37418
rect 22 37366 74 37418
rect 74 37366 76 37418
rect 20 37310 76 37366
rect 20 37258 22 37310
rect 22 37258 74 37310
rect 74 37258 76 37310
rect 20 37202 76 37258
rect 20 37150 22 37202
rect 22 37150 74 37202
rect 74 37150 76 37202
rect 20 37094 76 37150
rect 20 37042 22 37094
rect 22 37042 74 37094
rect 74 37042 76 37094
rect 20 36986 76 37042
rect 20 36934 22 36986
rect 22 36934 74 36986
rect 74 36934 76 36986
rect 20 36878 76 36934
rect 20 36826 22 36878
rect 22 36826 74 36878
rect 74 36826 76 36878
rect 20 36824 76 36826
rect 2491 49292 2547 49348
rect 2615 49292 2671 49348
rect 2491 49168 2547 49224
rect 2615 49168 2671 49224
rect 2491 49044 2547 49100
rect 2615 49044 2671 49100
rect 2491 48920 2547 48976
rect 2615 48920 2671 48976
rect 2491 48796 2547 48852
rect 2615 48796 2671 48852
rect 2491 48672 2547 48728
rect 2615 48672 2671 48728
rect 2491 48548 2547 48604
rect 2615 48548 2671 48604
rect 2491 48424 2547 48480
rect 2615 48424 2671 48480
rect 2491 48300 2547 48356
rect 2615 48300 2671 48356
rect 2491 48176 2547 48232
rect 2615 48176 2671 48232
rect 2491 48052 2547 48108
rect 2615 48052 2671 48108
rect 2808 55692 2864 55748
rect 2932 55692 2988 55748
rect 3056 55692 3112 55748
rect 3180 55692 3236 55748
rect 3304 55692 3360 55748
rect 3428 55692 3484 55748
rect 3552 55692 3608 55748
rect 3676 55692 3732 55748
rect 3800 55692 3856 55748
rect 3924 55692 3980 55748
rect 4048 55692 4104 55748
rect 4172 55692 4228 55748
rect 4296 55692 4352 55748
rect 4420 55692 4476 55748
rect 4544 55692 4600 55748
rect 4668 55692 4724 55748
rect 2808 55568 2864 55624
rect 2932 55568 2988 55624
rect 3056 55568 3112 55624
rect 3180 55568 3236 55624
rect 3304 55568 3360 55624
rect 3428 55568 3484 55624
rect 3552 55568 3608 55624
rect 3676 55568 3732 55624
rect 3800 55568 3856 55624
rect 3924 55568 3980 55624
rect 4048 55568 4104 55624
rect 4172 55568 4228 55624
rect 4296 55568 4352 55624
rect 4420 55568 4476 55624
rect 4544 55568 4600 55624
rect 4668 55568 4724 55624
rect 2808 55444 2864 55500
rect 2932 55444 2988 55500
rect 3056 55444 3112 55500
rect 3180 55444 3236 55500
rect 3304 55444 3360 55500
rect 3428 55444 3484 55500
rect 3552 55444 3608 55500
rect 3676 55444 3732 55500
rect 3800 55444 3856 55500
rect 3924 55444 3980 55500
rect 4048 55444 4104 55500
rect 4172 55444 4228 55500
rect 4296 55444 4352 55500
rect 4420 55444 4476 55500
rect 4544 55444 4600 55500
rect 4668 55444 4724 55500
rect 2808 55320 2864 55376
rect 2932 55320 2988 55376
rect 3056 55320 3112 55376
rect 3180 55320 3236 55376
rect 3304 55320 3360 55376
rect 3428 55320 3484 55376
rect 3552 55320 3608 55376
rect 3676 55320 3732 55376
rect 3800 55320 3856 55376
rect 3924 55320 3980 55376
rect 4048 55320 4104 55376
rect 4172 55320 4228 55376
rect 4296 55320 4352 55376
rect 4420 55320 4476 55376
rect 4544 55320 4600 55376
rect 4668 55320 4724 55376
rect 2808 55196 2864 55252
rect 2932 55196 2988 55252
rect 3056 55196 3112 55252
rect 3180 55196 3236 55252
rect 3304 55196 3360 55252
rect 3428 55196 3484 55252
rect 3552 55196 3608 55252
rect 3676 55196 3732 55252
rect 3800 55196 3856 55252
rect 3924 55196 3980 55252
rect 4048 55196 4104 55252
rect 4172 55196 4228 55252
rect 4296 55196 4352 55252
rect 4420 55196 4476 55252
rect 4544 55196 4600 55252
rect 4668 55196 4724 55252
rect 2808 55072 2864 55128
rect 2932 55072 2988 55128
rect 3056 55072 3112 55128
rect 3180 55072 3236 55128
rect 3304 55072 3360 55128
rect 3428 55072 3484 55128
rect 3552 55072 3608 55128
rect 3676 55072 3732 55128
rect 3800 55072 3856 55128
rect 3924 55072 3980 55128
rect 4048 55072 4104 55128
rect 4172 55072 4228 55128
rect 4296 55072 4352 55128
rect 4420 55072 4476 55128
rect 4544 55072 4600 55128
rect 4668 55072 4724 55128
rect 2808 54948 2864 55004
rect 2932 54948 2988 55004
rect 3056 54948 3112 55004
rect 3180 54948 3236 55004
rect 3304 54948 3360 55004
rect 3428 54948 3484 55004
rect 3552 54948 3608 55004
rect 3676 54948 3732 55004
rect 3800 54948 3856 55004
rect 3924 54948 3980 55004
rect 4048 54948 4104 55004
rect 4172 54948 4228 55004
rect 4296 54948 4352 55004
rect 4420 54948 4476 55004
rect 4544 54948 4600 55004
rect 4668 54948 4724 55004
rect 2808 54824 2864 54880
rect 2932 54824 2988 54880
rect 3056 54824 3112 54880
rect 3180 54824 3236 54880
rect 3304 54824 3360 54880
rect 3428 54824 3484 54880
rect 3552 54824 3608 54880
rect 3676 54824 3732 54880
rect 3800 54824 3856 54880
rect 3924 54824 3980 54880
rect 4048 54824 4104 54880
rect 4172 54824 4228 54880
rect 4296 54824 4352 54880
rect 4420 54824 4476 54880
rect 4544 54824 4600 54880
rect 4668 54824 4724 54880
rect 2808 54700 2864 54756
rect 2932 54700 2988 54756
rect 3056 54700 3112 54756
rect 3180 54700 3236 54756
rect 3304 54700 3360 54756
rect 3428 54700 3484 54756
rect 3552 54700 3608 54756
rect 3676 54700 3732 54756
rect 3800 54700 3856 54756
rect 3924 54700 3980 54756
rect 4048 54700 4104 54756
rect 4172 54700 4228 54756
rect 4296 54700 4352 54756
rect 4420 54700 4476 54756
rect 4544 54700 4600 54756
rect 4668 54700 4724 54756
rect 2808 54576 2864 54632
rect 2932 54576 2988 54632
rect 3056 54576 3112 54632
rect 3180 54576 3236 54632
rect 3304 54576 3360 54632
rect 3428 54576 3484 54632
rect 3552 54576 3608 54632
rect 3676 54576 3732 54632
rect 3800 54576 3856 54632
rect 3924 54576 3980 54632
rect 4048 54576 4104 54632
rect 4172 54576 4228 54632
rect 4296 54576 4352 54632
rect 4420 54576 4476 54632
rect 4544 54576 4600 54632
rect 4668 54576 4724 54632
rect 2808 54452 2864 54508
rect 2932 54452 2988 54508
rect 3056 54452 3112 54508
rect 3180 54452 3236 54508
rect 3304 54452 3360 54508
rect 3428 54452 3484 54508
rect 3552 54452 3608 54508
rect 3676 54452 3732 54508
rect 3800 54452 3856 54508
rect 3924 54452 3980 54508
rect 4048 54452 4104 54508
rect 4172 54452 4228 54508
rect 4296 54452 4352 54508
rect 4420 54452 4476 54508
rect 4544 54452 4600 54508
rect 4668 54452 4724 54508
rect 2808 50892 2864 50948
rect 2932 50892 2988 50948
rect 3056 50892 3112 50948
rect 3180 50892 3236 50948
rect 3304 50892 3360 50948
rect 3428 50892 3484 50948
rect 3552 50892 3608 50948
rect 3676 50892 3732 50948
rect 3800 50892 3856 50948
rect 3924 50892 3980 50948
rect 4048 50892 4104 50948
rect 4172 50892 4228 50948
rect 4296 50892 4352 50948
rect 4420 50892 4476 50948
rect 4544 50892 4600 50948
rect 4668 50892 4724 50948
rect 2808 50768 2864 50824
rect 2932 50768 2988 50824
rect 3056 50768 3112 50824
rect 3180 50768 3236 50824
rect 3304 50768 3360 50824
rect 3428 50768 3484 50824
rect 3552 50768 3608 50824
rect 3676 50768 3732 50824
rect 3800 50768 3856 50824
rect 3924 50768 3980 50824
rect 4048 50768 4104 50824
rect 4172 50768 4228 50824
rect 4296 50768 4352 50824
rect 4420 50768 4476 50824
rect 4544 50768 4600 50824
rect 4668 50768 4724 50824
rect 2808 50644 2864 50700
rect 2932 50644 2988 50700
rect 3056 50644 3112 50700
rect 3180 50644 3236 50700
rect 3304 50644 3360 50700
rect 3428 50644 3484 50700
rect 3552 50693 3608 50700
rect 3676 50693 3732 50700
rect 3800 50693 3856 50700
rect 3924 50693 3980 50700
rect 4048 50693 4104 50700
rect 4172 50693 4228 50700
rect 4296 50693 4352 50700
rect 4420 50693 4476 50700
rect 4544 50693 4600 50700
rect 4668 50693 4724 50700
rect 3552 50644 3559 50693
rect 3559 50644 3608 50693
rect 3676 50644 3683 50693
rect 3683 50644 3732 50693
rect 3800 50644 3807 50693
rect 3807 50644 3856 50693
rect 3924 50644 3931 50693
rect 3931 50644 3980 50693
rect 4048 50644 4055 50693
rect 4055 50644 4104 50693
rect 4172 50644 4179 50693
rect 4179 50644 4228 50693
rect 4296 50644 4303 50693
rect 4303 50644 4352 50693
rect 4420 50644 4427 50693
rect 4427 50644 4476 50693
rect 4544 50644 4551 50693
rect 4551 50644 4600 50693
rect 4668 50644 4675 50693
rect 4675 50644 4724 50693
rect 2808 50520 2864 50576
rect 2932 50520 2988 50576
rect 3056 50520 3112 50576
rect 3180 50520 3236 50576
rect 3304 50520 3360 50576
rect 3428 50520 3484 50576
rect 3552 50569 3608 50576
rect 3676 50569 3732 50576
rect 3800 50569 3856 50576
rect 3924 50569 3980 50576
rect 4048 50569 4104 50576
rect 4172 50569 4228 50576
rect 4296 50569 4352 50576
rect 4420 50569 4476 50576
rect 4544 50569 4600 50576
rect 4668 50569 4724 50576
rect 3552 50520 3559 50569
rect 3559 50520 3608 50569
rect 3676 50520 3683 50569
rect 3683 50520 3732 50569
rect 3800 50520 3807 50569
rect 3807 50520 3856 50569
rect 3924 50520 3931 50569
rect 3931 50520 3980 50569
rect 4048 50520 4055 50569
rect 4055 50520 4104 50569
rect 4172 50520 4179 50569
rect 4179 50520 4228 50569
rect 4296 50520 4303 50569
rect 4303 50520 4352 50569
rect 4420 50520 4427 50569
rect 4427 50520 4476 50569
rect 4544 50520 4551 50569
rect 4551 50520 4600 50569
rect 4668 50520 4675 50569
rect 4675 50520 4724 50569
rect 2808 50396 2864 50452
rect 2932 50396 2988 50452
rect 3056 50396 3112 50452
rect 3180 50396 3236 50452
rect 3304 50396 3360 50452
rect 3428 50396 3484 50452
rect 3552 50396 3608 50452
rect 3676 50396 3732 50452
rect 3800 50396 3856 50452
rect 3924 50396 3980 50452
rect 4048 50396 4104 50452
rect 4172 50396 4228 50452
rect 4296 50396 4352 50452
rect 4420 50396 4476 50452
rect 4544 50396 4600 50452
rect 4668 50396 4724 50452
rect 2808 50272 2864 50328
rect 2932 50272 2988 50328
rect 3056 50272 3112 50328
rect 3180 50272 3236 50328
rect 3304 50272 3360 50328
rect 3428 50272 3484 50328
rect 3552 50272 3608 50328
rect 3676 50272 3732 50328
rect 3800 50272 3856 50328
rect 3924 50272 3980 50328
rect 4048 50272 4104 50328
rect 4172 50272 4228 50328
rect 4296 50272 4352 50328
rect 4420 50272 4476 50328
rect 4544 50272 4600 50328
rect 4668 50272 4724 50328
rect 2808 50148 2864 50204
rect 2932 50148 2988 50204
rect 3056 50148 3112 50204
rect 3180 50148 3236 50204
rect 3304 50148 3360 50204
rect 3428 50148 3484 50204
rect 3552 50148 3608 50204
rect 3676 50148 3732 50204
rect 3800 50148 3856 50204
rect 3924 50148 3980 50204
rect 4048 50148 4104 50204
rect 4172 50148 4228 50204
rect 4296 50148 4352 50204
rect 4420 50148 4476 50204
rect 4544 50148 4600 50204
rect 4668 50148 4724 50204
rect 2808 50024 2864 50080
rect 2932 50024 2988 50080
rect 3056 50024 3112 50080
rect 3180 50024 3236 50080
rect 3304 50024 3360 50080
rect 3428 50024 3484 50080
rect 3552 50024 3608 50080
rect 3676 50024 3732 50080
rect 3800 50024 3856 50080
rect 3924 50024 3980 50080
rect 4048 50024 4104 50080
rect 4172 50024 4228 50080
rect 4296 50024 4352 50080
rect 4420 50024 4476 50080
rect 4544 50024 4600 50080
rect 4668 50024 4724 50080
rect 2808 49900 2864 49956
rect 2932 49900 2988 49956
rect 3056 49900 3112 49956
rect 3180 49900 3236 49956
rect 3304 49900 3360 49956
rect 3428 49900 3484 49956
rect 3552 49900 3608 49956
rect 3676 49900 3732 49956
rect 3800 49900 3856 49956
rect 3924 49900 3980 49956
rect 4048 49900 4104 49956
rect 4172 49900 4228 49956
rect 4296 49900 4352 49956
rect 4420 49900 4476 49956
rect 4544 49900 4600 49956
rect 4668 49900 4724 49956
rect 2808 49776 2864 49832
rect 2932 49776 2988 49832
rect 3056 49776 3112 49832
rect 3180 49776 3236 49832
rect 3304 49776 3360 49832
rect 3428 49776 3484 49832
rect 3552 49776 3608 49832
rect 3676 49776 3732 49832
rect 3800 49776 3856 49832
rect 3924 49776 3980 49832
rect 4048 49776 4104 49832
rect 4172 49776 4228 49832
rect 4296 49776 4352 49832
rect 4420 49776 4476 49832
rect 4544 49776 4600 49832
rect 4668 49776 4724 49832
rect 2808 49652 2864 49708
rect 2932 49652 2988 49708
rect 3056 49652 3112 49708
rect 3180 49652 3236 49708
rect 3304 49652 3360 49708
rect 3428 49652 3484 49708
rect 3552 49707 3559 49708
rect 3559 49707 3608 49708
rect 3676 49707 3683 49708
rect 3683 49707 3732 49708
rect 3800 49707 3807 49708
rect 3807 49707 3856 49708
rect 3924 49707 3931 49708
rect 3931 49707 3980 49708
rect 4048 49707 4055 49708
rect 4055 49707 4104 49708
rect 4172 49707 4179 49708
rect 4179 49707 4228 49708
rect 4296 49707 4303 49708
rect 4303 49707 4352 49708
rect 4420 49707 4427 49708
rect 4427 49707 4476 49708
rect 4544 49707 4551 49708
rect 4551 49707 4600 49708
rect 4668 49707 4675 49708
rect 4675 49707 4724 49708
rect 3552 49652 3608 49707
rect 3676 49652 3732 49707
rect 3800 49652 3856 49707
rect 3924 49652 3980 49707
rect 4048 49652 4104 49707
rect 4172 49652 4228 49707
rect 4296 49652 4352 49707
rect 4420 49652 4476 49707
rect 4544 49652 4600 49707
rect 4668 49652 4724 49707
rect 2808 47740 2864 47748
rect 2808 47692 2810 47740
rect 2810 47692 2862 47740
rect 2862 47692 2864 47740
rect 2932 47740 2988 47748
rect 2932 47692 2934 47740
rect 2934 47692 2986 47740
rect 2986 47692 2988 47740
rect 3056 47740 3112 47748
rect 3056 47692 3058 47740
rect 3058 47692 3110 47740
rect 3110 47692 3112 47740
rect 3180 47740 3236 47748
rect 3180 47692 3182 47740
rect 3182 47692 3234 47740
rect 3234 47692 3236 47740
rect 3304 47740 3360 47748
rect 3304 47692 3306 47740
rect 3306 47692 3358 47740
rect 3358 47692 3360 47740
rect 3428 47740 3484 47748
rect 3428 47692 3430 47740
rect 3430 47692 3482 47740
rect 3482 47692 3484 47740
rect 3552 47740 3608 47748
rect 3552 47692 3554 47740
rect 3554 47692 3606 47740
rect 3606 47692 3608 47740
rect 3676 47740 3732 47748
rect 3676 47692 3678 47740
rect 3678 47692 3730 47740
rect 3730 47692 3732 47740
rect 3800 47740 3856 47748
rect 3800 47692 3802 47740
rect 3802 47692 3854 47740
rect 3854 47692 3856 47740
rect 3924 47740 3980 47748
rect 3924 47692 3926 47740
rect 3926 47692 3978 47740
rect 3978 47692 3980 47740
rect 4048 47740 4104 47748
rect 4048 47692 4050 47740
rect 4050 47692 4102 47740
rect 4102 47692 4104 47740
rect 4172 47740 4228 47748
rect 4172 47692 4174 47740
rect 4174 47692 4226 47740
rect 4226 47692 4228 47740
rect 4296 47740 4352 47748
rect 4296 47692 4298 47740
rect 4298 47692 4350 47740
rect 4350 47692 4352 47740
rect 4420 47740 4476 47748
rect 4420 47692 4422 47740
rect 4422 47692 4474 47740
rect 4474 47692 4476 47740
rect 4544 47740 4600 47748
rect 4544 47692 4546 47740
rect 4546 47692 4598 47740
rect 4598 47692 4600 47740
rect 4668 47740 4724 47748
rect 4668 47692 4670 47740
rect 4670 47692 4722 47740
rect 4722 47692 4724 47740
rect 2808 47568 2864 47624
rect 2932 47568 2988 47624
rect 3056 47568 3112 47624
rect 3180 47568 3236 47624
rect 3304 47568 3360 47624
rect 3428 47568 3484 47624
rect 3552 47568 3608 47624
rect 3676 47568 3732 47624
rect 3800 47568 3856 47624
rect 3924 47568 3980 47624
rect 4048 47568 4104 47624
rect 4172 47568 4228 47624
rect 4296 47568 4352 47624
rect 4420 47568 4476 47624
rect 4544 47568 4600 47624
rect 4668 47568 4724 47624
rect 2808 47444 2864 47500
rect 2932 47444 2988 47500
rect 3056 47444 3112 47500
rect 3180 47444 3236 47500
rect 3304 47444 3360 47500
rect 3428 47444 3484 47500
rect 3552 47444 3608 47500
rect 3676 47444 3732 47500
rect 3800 47444 3856 47500
rect 3924 47444 3980 47500
rect 4048 47444 4104 47500
rect 4172 47444 4228 47500
rect 4296 47444 4352 47500
rect 4420 47444 4476 47500
rect 4544 47444 4600 47500
rect 4668 47444 4724 47500
rect 2808 47320 2864 47376
rect 2932 47320 2988 47376
rect 3056 47320 3112 47376
rect 3180 47320 3236 47376
rect 3304 47320 3360 47376
rect 3428 47320 3484 47376
rect 3552 47320 3608 47376
rect 3676 47320 3732 47376
rect 3800 47320 3856 47376
rect 3924 47320 3980 47376
rect 4048 47320 4104 47376
rect 4172 47320 4228 47376
rect 4296 47320 4352 47376
rect 4420 47320 4476 47376
rect 4544 47320 4600 47376
rect 4668 47320 4724 47376
rect 4861 57169 4917 57225
rect 4985 57169 5041 57225
rect 4861 57056 4871 57101
rect 4871 57056 4917 57101
rect 4985 57056 5031 57101
rect 5031 57056 5041 57101
rect 4861 57045 4917 57056
rect 4985 57045 5041 57056
rect 4861 56921 4917 56977
rect 4985 56921 5041 56977
rect 4861 56797 4917 56853
rect 4985 56797 5041 56853
rect 4861 56673 4917 56729
rect 4985 56673 5041 56729
rect 4861 56549 4917 56605
rect 4985 56549 5041 56605
rect 4861 56425 4917 56481
rect 4985 56425 5041 56481
rect 4861 56301 4917 56357
rect 4985 56301 5041 56357
rect 4861 56177 4917 56233
rect 4985 56177 5041 56233
rect 4861 56053 4917 56109
rect 4985 56053 5041 56109
rect 4861 54092 4917 54148
rect 4985 54092 5041 54148
rect 4861 53968 4917 54024
rect 4985 53968 5041 54024
rect 4861 53844 4917 53900
rect 4985 53844 5041 53900
rect 4861 53720 4917 53776
rect 4985 53720 5041 53776
rect 4861 53596 4917 53652
rect 4985 53596 5041 53652
rect 4861 53484 4917 53528
rect 4985 53484 5041 53528
rect 4861 53472 4871 53484
rect 4871 53472 4917 53484
rect 4985 53472 5031 53484
rect 5031 53472 5041 53484
rect 4861 53376 4917 53404
rect 4985 53376 5041 53404
rect 4861 53348 4871 53376
rect 4871 53348 4917 53376
rect 4985 53348 5031 53376
rect 5031 53348 5041 53376
rect 4861 53268 4917 53280
rect 4985 53268 5041 53280
rect 4861 53224 4871 53268
rect 4871 53224 4917 53268
rect 4985 53224 5031 53268
rect 5031 53224 5041 53268
rect 4861 53100 4917 53156
rect 4985 53100 5041 53156
rect 4861 52976 4917 53032
rect 4985 52976 5041 53032
rect 4861 52852 4917 52908
rect 4985 52852 5041 52908
rect 4861 49302 4863 49348
rect 4863 49302 4915 49348
rect 4915 49302 4917 49348
rect 4861 49292 4917 49302
rect 4985 49302 4987 49348
rect 4987 49302 5039 49348
rect 5039 49302 5041 49348
rect 4985 49292 5041 49302
rect 4861 49178 4863 49224
rect 4863 49178 4915 49224
rect 4915 49178 4917 49224
rect 4861 49168 4917 49178
rect 4985 49178 4987 49224
rect 4987 49178 5039 49224
rect 5039 49178 5041 49224
rect 4985 49168 5041 49178
rect 4861 49054 4863 49100
rect 4863 49054 4915 49100
rect 4915 49054 4917 49100
rect 4861 49044 4917 49054
rect 4985 49054 4987 49100
rect 4987 49054 5039 49100
rect 5039 49054 5041 49100
rect 4985 49044 5041 49054
rect 4861 48920 4917 48976
rect 4985 48920 5041 48976
rect 4861 48796 4917 48852
rect 4985 48796 5041 48852
rect 4861 48672 4917 48728
rect 4985 48672 5041 48728
rect 4861 48548 4917 48604
rect 4985 48548 5041 48604
rect 4861 48435 4917 48480
rect 4861 48424 4863 48435
rect 4863 48424 4915 48435
rect 4915 48424 4917 48435
rect 4985 48435 5041 48480
rect 4985 48424 4987 48435
rect 4987 48424 5039 48435
rect 5039 48424 5041 48435
rect 4861 48311 4917 48356
rect 4861 48300 4863 48311
rect 4863 48300 4915 48311
rect 4915 48300 4917 48311
rect 4985 48311 5041 48356
rect 4985 48300 4987 48311
rect 4987 48300 5039 48311
rect 5039 48300 5041 48311
rect 4861 48176 4917 48232
rect 4985 48176 5041 48232
rect 4861 48052 4917 48108
rect 4985 48052 5041 48108
rect 5178 55692 5234 55748
rect 5302 55692 5358 55748
rect 5426 55692 5482 55748
rect 5550 55692 5606 55748
rect 5674 55692 5730 55748
rect 5798 55692 5854 55748
rect 5922 55692 5978 55748
rect 6046 55692 6102 55748
rect 6170 55692 6226 55748
rect 6294 55692 6350 55748
rect 6418 55692 6474 55748
rect 6542 55692 6598 55748
rect 6666 55692 6722 55748
rect 6790 55692 6846 55748
rect 6914 55692 6970 55748
rect 7038 55692 7094 55748
rect 5178 55568 5234 55624
rect 5302 55568 5358 55624
rect 5426 55568 5482 55624
rect 5550 55568 5606 55624
rect 5674 55568 5730 55624
rect 5798 55568 5854 55624
rect 5922 55568 5978 55624
rect 6046 55568 6102 55624
rect 6170 55568 6226 55624
rect 6294 55568 6350 55624
rect 6418 55568 6474 55624
rect 6542 55568 6598 55624
rect 6666 55568 6722 55624
rect 6790 55568 6846 55624
rect 6914 55568 6970 55624
rect 7038 55568 7094 55624
rect 5178 55444 5234 55500
rect 5302 55444 5358 55500
rect 5426 55444 5482 55500
rect 5550 55444 5606 55500
rect 5674 55444 5730 55500
rect 5798 55444 5854 55500
rect 5922 55444 5978 55500
rect 6046 55444 6102 55500
rect 6170 55444 6226 55500
rect 6294 55444 6350 55500
rect 6418 55444 6474 55500
rect 6542 55444 6598 55500
rect 6666 55444 6722 55500
rect 6790 55444 6846 55500
rect 6914 55444 6970 55500
rect 7038 55444 7094 55500
rect 5178 55320 5234 55376
rect 5302 55320 5358 55376
rect 5426 55320 5482 55376
rect 5550 55320 5606 55376
rect 5674 55320 5730 55376
rect 5798 55320 5854 55376
rect 5922 55320 5978 55376
rect 6046 55320 6102 55376
rect 6170 55320 6226 55376
rect 6294 55320 6350 55376
rect 6418 55320 6474 55376
rect 6542 55320 6598 55376
rect 6666 55320 6722 55376
rect 6790 55320 6846 55376
rect 6914 55320 6970 55376
rect 7038 55320 7094 55376
rect 5178 55196 5234 55252
rect 5302 55196 5358 55252
rect 5426 55196 5482 55252
rect 5550 55196 5606 55252
rect 5674 55196 5730 55252
rect 5798 55196 5854 55252
rect 5922 55196 5978 55252
rect 6046 55196 6102 55252
rect 6170 55196 6226 55252
rect 6294 55196 6350 55252
rect 6418 55196 6474 55252
rect 6542 55196 6598 55252
rect 6666 55196 6722 55252
rect 6790 55196 6846 55252
rect 6914 55196 6970 55252
rect 7038 55196 7094 55252
rect 5178 55072 5234 55128
rect 5302 55072 5358 55128
rect 5426 55072 5482 55128
rect 5550 55072 5606 55128
rect 5674 55072 5730 55128
rect 5798 55072 5854 55128
rect 5922 55072 5978 55128
rect 6046 55072 6102 55128
rect 6170 55072 6226 55128
rect 6294 55072 6350 55128
rect 6418 55072 6474 55128
rect 6542 55072 6598 55128
rect 6666 55072 6722 55128
rect 6790 55072 6846 55128
rect 6914 55072 6970 55128
rect 7038 55072 7094 55128
rect 5178 54948 5234 55004
rect 5302 54948 5358 55004
rect 5426 54948 5482 55004
rect 5550 54948 5606 55004
rect 5674 54948 5730 55004
rect 5798 54948 5854 55004
rect 5922 54948 5978 55004
rect 6046 54948 6102 55004
rect 6170 54948 6226 55004
rect 6294 54948 6350 55004
rect 6418 54948 6474 55004
rect 6542 54948 6598 55004
rect 6666 54948 6722 55004
rect 6790 54948 6846 55004
rect 6914 54948 6970 55004
rect 7038 54948 7094 55004
rect 5178 54824 5234 54880
rect 5302 54824 5358 54880
rect 5426 54824 5482 54880
rect 5550 54824 5606 54880
rect 5674 54824 5730 54880
rect 5798 54824 5854 54880
rect 5922 54824 5978 54880
rect 6046 54824 6102 54880
rect 6170 54824 6226 54880
rect 6294 54824 6350 54880
rect 6418 54824 6474 54880
rect 6542 54824 6598 54880
rect 6666 54824 6722 54880
rect 6790 54824 6846 54880
rect 6914 54824 6970 54880
rect 7038 54824 7094 54880
rect 5178 54700 5234 54756
rect 5302 54700 5358 54756
rect 5426 54700 5482 54756
rect 5550 54700 5606 54756
rect 5674 54700 5730 54756
rect 5798 54700 5854 54756
rect 5922 54700 5978 54756
rect 6046 54700 6102 54756
rect 6170 54700 6226 54756
rect 6294 54700 6350 54756
rect 6418 54700 6474 54756
rect 6542 54700 6598 54756
rect 6666 54700 6722 54756
rect 6790 54700 6846 54756
rect 6914 54700 6970 54756
rect 7038 54700 7094 54756
rect 5178 54576 5234 54632
rect 5302 54576 5358 54632
rect 5426 54576 5482 54632
rect 5550 54576 5606 54632
rect 5674 54576 5730 54632
rect 5798 54576 5854 54632
rect 5922 54576 5978 54632
rect 6046 54576 6102 54632
rect 6170 54576 6226 54632
rect 6294 54576 6350 54632
rect 6418 54576 6474 54632
rect 6542 54576 6598 54632
rect 6666 54576 6722 54632
rect 6790 54576 6846 54632
rect 6914 54576 6970 54632
rect 7038 54576 7094 54632
rect 5178 54452 5234 54508
rect 5302 54452 5358 54508
rect 5426 54452 5482 54508
rect 5550 54452 5606 54508
rect 5674 54452 5730 54508
rect 5798 54452 5854 54508
rect 5922 54452 5978 54508
rect 6046 54452 6102 54508
rect 6170 54452 6226 54508
rect 6294 54452 6350 54508
rect 6418 54452 6474 54508
rect 6542 54452 6598 54508
rect 6666 54452 6722 54508
rect 6790 54452 6846 54508
rect 6914 54452 6970 54508
rect 7038 54452 7094 54508
rect 5178 50892 5234 50948
rect 5302 50892 5358 50948
rect 5426 50892 5482 50948
rect 5550 50892 5606 50948
rect 5674 50892 5730 50948
rect 5798 50892 5854 50948
rect 5922 50892 5978 50948
rect 6046 50892 6102 50948
rect 6170 50892 6226 50948
rect 6294 50892 6350 50948
rect 6418 50892 6474 50948
rect 6542 50892 6598 50948
rect 6666 50892 6722 50948
rect 6790 50892 6846 50948
rect 6914 50892 6970 50948
rect 7038 50892 7094 50948
rect 5178 50768 5234 50824
rect 5302 50768 5358 50824
rect 5426 50768 5482 50824
rect 5550 50768 5606 50824
rect 5674 50768 5730 50824
rect 5798 50768 5854 50824
rect 5922 50768 5978 50824
rect 6046 50768 6102 50824
rect 6170 50768 6226 50824
rect 6294 50768 6350 50824
rect 6418 50768 6474 50824
rect 6542 50768 6598 50824
rect 6666 50768 6722 50824
rect 6790 50768 6846 50824
rect 6914 50768 6970 50824
rect 7038 50768 7094 50824
rect 5178 50693 5234 50700
rect 5178 50644 5180 50693
rect 5180 50644 5232 50693
rect 5232 50644 5234 50693
rect 5302 50693 5358 50700
rect 5302 50644 5304 50693
rect 5304 50644 5356 50693
rect 5356 50644 5358 50693
rect 5426 50693 5482 50700
rect 5426 50644 5428 50693
rect 5428 50644 5480 50693
rect 5480 50644 5482 50693
rect 5550 50693 5606 50700
rect 5550 50644 5552 50693
rect 5552 50644 5604 50693
rect 5604 50644 5606 50693
rect 5674 50693 5730 50700
rect 5674 50644 5676 50693
rect 5676 50644 5728 50693
rect 5728 50644 5730 50693
rect 5798 50693 5854 50700
rect 5798 50644 5800 50693
rect 5800 50644 5852 50693
rect 5852 50644 5854 50693
rect 5922 50693 5978 50700
rect 5922 50644 5924 50693
rect 5924 50644 5976 50693
rect 5976 50644 5978 50693
rect 6046 50693 6102 50700
rect 6046 50644 6048 50693
rect 6048 50644 6100 50693
rect 6100 50644 6102 50693
rect 6170 50693 6226 50700
rect 6170 50644 6172 50693
rect 6172 50644 6224 50693
rect 6224 50644 6226 50693
rect 6294 50693 6350 50700
rect 6294 50644 6296 50693
rect 6296 50644 6348 50693
rect 6348 50644 6350 50693
rect 6418 50693 6474 50700
rect 6418 50644 6420 50693
rect 6420 50644 6472 50693
rect 6472 50644 6474 50693
rect 6542 50693 6598 50700
rect 6542 50644 6544 50693
rect 6544 50644 6596 50693
rect 6596 50644 6598 50693
rect 6666 50693 6722 50700
rect 6666 50644 6668 50693
rect 6668 50644 6720 50693
rect 6720 50644 6722 50693
rect 6790 50693 6846 50700
rect 6790 50644 6792 50693
rect 6792 50644 6844 50693
rect 6844 50644 6846 50693
rect 6914 50693 6970 50700
rect 6914 50644 6916 50693
rect 6916 50644 6968 50693
rect 6968 50644 6970 50693
rect 7038 50693 7094 50700
rect 7038 50644 7040 50693
rect 7040 50644 7092 50693
rect 7092 50644 7094 50693
rect 5178 50569 5234 50576
rect 5178 50520 5180 50569
rect 5180 50520 5232 50569
rect 5232 50520 5234 50569
rect 5302 50569 5358 50576
rect 5302 50520 5304 50569
rect 5304 50520 5356 50569
rect 5356 50520 5358 50569
rect 5426 50569 5482 50576
rect 5426 50520 5428 50569
rect 5428 50520 5480 50569
rect 5480 50520 5482 50569
rect 5550 50569 5606 50576
rect 5550 50520 5552 50569
rect 5552 50520 5604 50569
rect 5604 50520 5606 50569
rect 5674 50569 5730 50576
rect 5674 50520 5676 50569
rect 5676 50520 5728 50569
rect 5728 50520 5730 50569
rect 5798 50569 5854 50576
rect 5798 50520 5800 50569
rect 5800 50520 5852 50569
rect 5852 50520 5854 50569
rect 5922 50569 5978 50576
rect 5922 50520 5924 50569
rect 5924 50520 5976 50569
rect 5976 50520 5978 50569
rect 6046 50569 6102 50576
rect 6046 50520 6048 50569
rect 6048 50520 6100 50569
rect 6100 50520 6102 50569
rect 6170 50569 6226 50576
rect 6170 50520 6172 50569
rect 6172 50520 6224 50569
rect 6224 50520 6226 50569
rect 6294 50569 6350 50576
rect 6294 50520 6296 50569
rect 6296 50520 6348 50569
rect 6348 50520 6350 50569
rect 6418 50569 6474 50576
rect 6418 50520 6420 50569
rect 6420 50520 6472 50569
rect 6472 50520 6474 50569
rect 6542 50569 6598 50576
rect 6542 50520 6544 50569
rect 6544 50520 6596 50569
rect 6596 50520 6598 50569
rect 6666 50569 6722 50576
rect 6666 50520 6668 50569
rect 6668 50520 6720 50569
rect 6720 50520 6722 50569
rect 6790 50569 6846 50576
rect 6790 50520 6792 50569
rect 6792 50520 6844 50569
rect 6844 50520 6846 50569
rect 6914 50569 6970 50576
rect 6914 50520 6916 50569
rect 6916 50520 6968 50569
rect 6968 50520 6970 50569
rect 7038 50569 7094 50576
rect 7038 50520 7040 50569
rect 7040 50520 7092 50569
rect 7092 50520 7094 50569
rect 5178 50396 5234 50452
rect 5302 50396 5358 50452
rect 5426 50396 5482 50452
rect 5550 50396 5606 50452
rect 5674 50396 5730 50452
rect 5798 50396 5854 50452
rect 5922 50396 5978 50452
rect 6046 50396 6102 50452
rect 6170 50396 6226 50452
rect 6294 50396 6350 50452
rect 6418 50396 6474 50452
rect 6542 50396 6598 50452
rect 6666 50396 6722 50452
rect 6790 50396 6846 50452
rect 6914 50396 6970 50452
rect 7038 50396 7094 50452
rect 5178 50272 5234 50328
rect 5302 50272 5358 50328
rect 5426 50272 5482 50328
rect 5550 50272 5606 50328
rect 5674 50272 5730 50328
rect 5798 50272 5854 50328
rect 5922 50272 5978 50328
rect 6046 50272 6102 50328
rect 6170 50272 6226 50328
rect 6294 50272 6350 50328
rect 6418 50272 6474 50328
rect 6542 50272 6598 50328
rect 6666 50272 6722 50328
rect 6790 50272 6846 50328
rect 6914 50272 6970 50328
rect 7038 50272 7094 50328
rect 5178 50148 5234 50204
rect 5302 50148 5358 50204
rect 5426 50148 5482 50204
rect 5550 50148 5606 50204
rect 5674 50148 5730 50204
rect 5798 50148 5854 50204
rect 5922 50148 5978 50204
rect 6046 50148 6102 50204
rect 6170 50148 6226 50204
rect 6294 50148 6350 50204
rect 6418 50148 6474 50204
rect 6542 50148 6598 50204
rect 6666 50148 6722 50204
rect 6790 50148 6846 50204
rect 6914 50148 6970 50204
rect 7038 50148 7094 50204
rect 5178 50024 5234 50080
rect 5302 50024 5358 50080
rect 5426 50024 5482 50080
rect 5550 50024 5606 50080
rect 5674 50024 5730 50080
rect 5798 50024 5854 50080
rect 5922 50024 5978 50080
rect 6046 50024 6102 50080
rect 6170 50024 6226 50080
rect 6294 50024 6350 50080
rect 6418 50024 6474 50080
rect 6542 50024 6598 50080
rect 6666 50024 6722 50080
rect 6790 50024 6846 50080
rect 6914 50024 6970 50080
rect 7038 50024 7094 50080
rect 5178 49900 5234 49956
rect 5302 49900 5358 49956
rect 5426 49900 5482 49956
rect 5550 49900 5606 49956
rect 5674 49900 5730 49956
rect 5798 49900 5854 49956
rect 5922 49900 5978 49956
rect 6046 49900 6102 49956
rect 6170 49900 6226 49956
rect 6294 49900 6350 49956
rect 6418 49900 6474 49956
rect 6542 49900 6598 49956
rect 6666 49900 6722 49956
rect 6790 49900 6846 49956
rect 6914 49900 6970 49956
rect 7038 49900 7094 49956
rect 5178 49776 5234 49832
rect 5302 49776 5358 49832
rect 5426 49776 5482 49832
rect 5550 49776 5606 49832
rect 5674 49776 5730 49832
rect 5798 49776 5854 49832
rect 5922 49776 5978 49832
rect 6046 49776 6102 49832
rect 6170 49776 6226 49832
rect 6294 49776 6350 49832
rect 6418 49776 6474 49832
rect 6542 49776 6598 49832
rect 6666 49776 6722 49832
rect 6790 49776 6846 49832
rect 6914 49776 6970 49832
rect 7038 49776 7094 49832
rect 5178 49707 5180 49708
rect 5180 49707 5232 49708
rect 5232 49707 5234 49708
rect 5178 49652 5234 49707
rect 5302 49707 5304 49708
rect 5304 49707 5356 49708
rect 5356 49707 5358 49708
rect 5302 49652 5358 49707
rect 5426 49707 5428 49708
rect 5428 49707 5480 49708
rect 5480 49707 5482 49708
rect 5426 49652 5482 49707
rect 5550 49707 5552 49708
rect 5552 49707 5604 49708
rect 5604 49707 5606 49708
rect 5550 49652 5606 49707
rect 5674 49707 5676 49708
rect 5676 49707 5728 49708
rect 5728 49707 5730 49708
rect 5674 49652 5730 49707
rect 5798 49707 5800 49708
rect 5800 49707 5852 49708
rect 5852 49707 5854 49708
rect 5798 49652 5854 49707
rect 5922 49707 5924 49708
rect 5924 49707 5976 49708
rect 5976 49707 5978 49708
rect 5922 49652 5978 49707
rect 6046 49707 6048 49708
rect 6048 49707 6100 49708
rect 6100 49707 6102 49708
rect 6046 49652 6102 49707
rect 6170 49707 6172 49708
rect 6172 49707 6224 49708
rect 6224 49707 6226 49708
rect 6170 49652 6226 49707
rect 6294 49707 6296 49708
rect 6296 49707 6348 49708
rect 6348 49707 6350 49708
rect 6294 49652 6350 49707
rect 6418 49707 6420 49708
rect 6420 49707 6472 49708
rect 6472 49707 6474 49708
rect 6418 49652 6474 49707
rect 6542 49707 6544 49708
rect 6544 49707 6596 49708
rect 6596 49707 6598 49708
rect 6542 49652 6598 49707
rect 6666 49707 6668 49708
rect 6668 49707 6720 49708
rect 6720 49707 6722 49708
rect 6666 49652 6722 49707
rect 6790 49707 6792 49708
rect 6792 49707 6844 49708
rect 6844 49707 6846 49708
rect 6790 49652 6846 49707
rect 6914 49707 6916 49708
rect 6916 49707 6968 49708
rect 6968 49707 6970 49708
rect 6914 49652 6970 49707
rect 7038 49707 7040 49708
rect 7040 49707 7092 49708
rect 7092 49707 7094 49708
rect 7038 49652 7094 49707
rect 5178 47740 5234 47748
rect 5178 47692 5180 47740
rect 5180 47692 5232 47740
rect 5232 47692 5234 47740
rect 5302 47740 5358 47748
rect 5302 47692 5304 47740
rect 5304 47692 5356 47740
rect 5356 47692 5358 47740
rect 5426 47740 5482 47748
rect 5426 47692 5428 47740
rect 5428 47692 5480 47740
rect 5480 47692 5482 47740
rect 5550 47740 5606 47748
rect 5550 47692 5552 47740
rect 5552 47692 5604 47740
rect 5604 47692 5606 47740
rect 5674 47740 5730 47748
rect 5674 47692 5676 47740
rect 5676 47692 5728 47740
rect 5728 47692 5730 47740
rect 5798 47740 5854 47748
rect 5798 47692 5800 47740
rect 5800 47692 5852 47740
rect 5852 47692 5854 47740
rect 5922 47740 5978 47748
rect 5922 47692 5924 47740
rect 5924 47692 5976 47740
rect 5976 47692 5978 47740
rect 6046 47740 6102 47748
rect 6046 47692 6048 47740
rect 6048 47692 6100 47740
rect 6100 47692 6102 47740
rect 6170 47740 6226 47748
rect 6170 47692 6172 47740
rect 6172 47692 6224 47740
rect 6224 47692 6226 47740
rect 6294 47740 6350 47748
rect 6294 47692 6296 47740
rect 6296 47692 6348 47740
rect 6348 47692 6350 47740
rect 6418 47740 6474 47748
rect 6418 47692 6420 47740
rect 6420 47692 6472 47740
rect 6472 47692 6474 47740
rect 6542 47740 6598 47748
rect 6542 47692 6544 47740
rect 6544 47692 6596 47740
rect 6596 47692 6598 47740
rect 6666 47740 6722 47748
rect 6666 47692 6668 47740
rect 6668 47692 6720 47740
rect 6720 47692 6722 47740
rect 6790 47740 6846 47748
rect 6790 47692 6792 47740
rect 6792 47692 6844 47740
rect 6844 47692 6846 47740
rect 6914 47740 6970 47748
rect 6914 47692 6916 47740
rect 6916 47692 6968 47740
rect 6968 47692 6970 47740
rect 7038 47740 7094 47748
rect 7038 47692 7040 47740
rect 7040 47692 7092 47740
rect 7092 47692 7094 47740
rect 5178 47568 5234 47624
rect 5302 47568 5358 47624
rect 5426 47568 5482 47624
rect 5550 47568 5606 47624
rect 5674 47568 5730 47624
rect 5798 47568 5854 47624
rect 5922 47568 5978 47624
rect 6046 47568 6102 47624
rect 6170 47568 6226 47624
rect 6294 47568 6350 47624
rect 6418 47568 6474 47624
rect 6542 47568 6598 47624
rect 6666 47568 6722 47624
rect 6790 47568 6846 47624
rect 6914 47568 6970 47624
rect 7038 47568 7094 47624
rect 5178 47444 5234 47500
rect 5302 47444 5358 47500
rect 5426 47444 5482 47500
rect 5550 47444 5606 47500
rect 5674 47444 5730 47500
rect 5798 47444 5854 47500
rect 5922 47444 5978 47500
rect 6046 47444 6102 47500
rect 6170 47444 6226 47500
rect 6294 47444 6350 47500
rect 6418 47444 6474 47500
rect 6542 47444 6598 47500
rect 6666 47444 6722 47500
rect 6790 47444 6846 47500
rect 6914 47444 6970 47500
rect 7038 47444 7094 47500
rect 5178 47320 5234 47376
rect 5302 47320 5358 47376
rect 5426 47320 5482 47376
rect 5550 47320 5606 47376
rect 5674 47320 5730 47376
rect 5798 47320 5854 47376
rect 5922 47320 5978 47376
rect 6046 47320 6102 47376
rect 6170 47320 6226 47376
rect 6294 47320 6350 47376
rect 6418 47320 6474 47376
rect 6542 47320 6598 47376
rect 6666 47320 6722 47376
rect 6790 47320 6846 47376
rect 6914 47320 6970 47376
rect 7038 47320 7094 47376
rect 7275 57169 7331 57225
rect 7399 57169 7455 57225
rect 7523 57169 7579 57225
rect 7647 57169 7703 57225
rect 7275 57056 7299 57101
rect 7299 57056 7331 57101
rect 7399 57056 7407 57101
rect 7407 57056 7455 57101
rect 7523 57056 7571 57101
rect 7571 57056 7579 57101
rect 7647 57056 7679 57101
rect 7679 57056 7703 57101
rect 7275 57045 7331 57056
rect 7399 57045 7455 57056
rect 7523 57045 7579 57056
rect 7647 57045 7703 57056
rect 7275 56921 7331 56977
rect 7399 56921 7455 56977
rect 7523 56921 7579 56977
rect 7647 56921 7703 56977
rect 7275 56797 7331 56853
rect 7399 56797 7455 56853
rect 7523 56797 7579 56853
rect 7647 56797 7703 56853
rect 7275 56673 7331 56729
rect 7399 56673 7455 56729
rect 7523 56673 7579 56729
rect 7647 56673 7703 56729
rect 7275 56549 7331 56605
rect 7399 56549 7455 56605
rect 7523 56549 7579 56605
rect 7647 56549 7703 56605
rect 7275 56425 7331 56481
rect 7399 56425 7455 56481
rect 7523 56425 7579 56481
rect 7647 56425 7703 56481
rect 7275 56301 7331 56357
rect 7399 56301 7455 56357
rect 7523 56301 7579 56357
rect 7647 56301 7703 56357
rect 7275 56177 7331 56233
rect 7399 56177 7455 56233
rect 7523 56177 7579 56233
rect 7647 56177 7703 56233
rect 7275 56053 7331 56109
rect 7399 56053 7455 56109
rect 7523 56053 7579 56109
rect 7647 56053 7703 56109
rect 7275 54092 7331 54148
rect 7399 54092 7455 54148
rect 7523 54092 7579 54148
rect 7647 54092 7703 54148
rect 7275 53968 7331 54024
rect 7399 53968 7455 54024
rect 7523 53968 7579 54024
rect 7647 53968 7703 54024
rect 7275 53844 7331 53900
rect 7399 53844 7455 53900
rect 7523 53844 7579 53900
rect 7647 53844 7703 53900
rect 7275 53720 7331 53776
rect 7399 53720 7455 53776
rect 7523 53720 7579 53776
rect 7647 53720 7703 53776
rect 7275 53596 7331 53652
rect 7399 53596 7455 53652
rect 7523 53596 7579 53652
rect 7647 53596 7703 53652
rect 7275 53484 7331 53528
rect 7399 53484 7455 53528
rect 7523 53484 7579 53528
rect 7647 53484 7703 53528
rect 7275 53472 7299 53484
rect 7299 53472 7331 53484
rect 7399 53472 7407 53484
rect 7407 53472 7455 53484
rect 7523 53472 7571 53484
rect 7571 53472 7579 53484
rect 7647 53472 7679 53484
rect 7679 53472 7703 53484
rect 7275 53376 7331 53404
rect 7399 53376 7455 53404
rect 7523 53376 7579 53404
rect 7647 53376 7703 53404
rect 7275 53348 7299 53376
rect 7299 53348 7331 53376
rect 7399 53348 7407 53376
rect 7407 53348 7455 53376
rect 7523 53348 7571 53376
rect 7571 53348 7579 53376
rect 7647 53348 7679 53376
rect 7679 53348 7703 53376
rect 7275 53268 7331 53280
rect 7399 53268 7455 53280
rect 7523 53268 7579 53280
rect 7647 53268 7703 53280
rect 7275 53224 7299 53268
rect 7299 53224 7331 53268
rect 7399 53224 7407 53268
rect 7407 53224 7455 53268
rect 7523 53224 7571 53268
rect 7571 53224 7579 53268
rect 7647 53224 7679 53268
rect 7679 53224 7703 53268
rect 7275 53100 7331 53156
rect 7399 53100 7455 53156
rect 7523 53100 7579 53156
rect 7647 53100 7703 53156
rect 7275 52976 7331 53032
rect 7399 52976 7455 53032
rect 7523 52976 7579 53032
rect 7647 52976 7703 53032
rect 7275 52852 7331 52908
rect 7399 52852 7455 52908
rect 7523 52852 7579 52908
rect 7647 52852 7703 52908
rect 7275 49302 7277 49348
rect 7277 49302 7329 49348
rect 7329 49302 7331 49348
rect 7275 49292 7331 49302
rect 7399 49302 7401 49348
rect 7401 49302 7453 49348
rect 7453 49302 7455 49348
rect 7399 49292 7455 49302
rect 7523 49302 7525 49348
rect 7525 49302 7577 49348
rect 7577 49302 7579 49348
rect 7523 49292 7579 49302
rect 7647 49302 7649 49348
rect 7649 49302 7701 49348
rect 7701 49302 7703 49348
rect 7647 49292 7703 49302
rect 7275 49178 7277 49224
rect 7277 49178 7329 49224
rect 7329 49178 7331 49224
rect 7275 49168 7331 49178
rect 7399 49178 7401 49224
rect 7401 49178 7453 49224
rect 7453 49178 7455 49224
rect 7399 49168 7455 49178
rect 7523 49178 7525 49224
rect 7525 49178 7577 49224
rect 7577 49178 7579 49224
rect 7523 49168 7579 49178
rect 7647 49178 7649 49224
rect 7649 49178 7701 49224
rect 7701 49178 7703 49224
rect 7647 49168 7703 49178
rect 7275 49054 7277 49100
rect 7277 49054 7329 49100
rect 7329 49054 7331 49100
rect 7275 49044 7331 49054
rect 7399 49054 7401 49100
rect 7401 49054 7453 49100
rect 7453 49054 7455 49100
rect 7399 49044 7455 49054
rect 7523 49054 7525 49100
rect 7525 49054 7577 49100
rect 7577 49054 7579 49100
rect 7523 49044 7579 49054
rect 7647 49054 7649 49100
rect 7649 49054 7701 49100
rect 7701 49054 7703 49100
rect 7647 49044 7703 49054
rect 7275 48920 7331 48976
rect 7399 48920 7455 48976
rect 7523 48920 7579 48976
rect 7647 48920 7703 48976
rect 7275 48796 7331 48852
rect 7399 48796 7455 48852
rect 7523 48796 7579 48852
rect 7647 48796 7703 48852
rect 7275 48672 7331 48728
rect 7399 48672 7455 48728
rect 7523 48672 7579 48728
rect 7647 48672 7703 48728
rect 7275 48548 7331 48604
rect 7399 48548 7455 48604
rect 7523 48548 7579 48604
rect 7647 48548 7703 48604
rect 7275 48435 7331 48480
rect 7275 48424 7277 48435
rect 7277 48424 7329 48435
rect 7329 48424 7331 48435
rect 7399 48435 7455 48480
rect 7399 48424 7401 48435
rect 7401 48424 7453 48435
rect 7453 48424 7455 48435
rect 7523 48435 7579 48480
rect 7523 48424 7525 48435
rect 7525 48424 7577 48435
rect 7577 48424 7579 48435
rect 7647 48435 7703 48480
rect 7647 48424 7649 48435
rect 7649 48424 7701 48435
rect 7701 48424 7703 48435
rect 7275 48311 7331 48356
rect 7275 48300 7277 48311
rect 7277 48300 7329 48311
rect 7329 48300 7331 48311
rect 7399 48311 7455 48356
rect 7399 48300 7401 48311
rect 7401 48300 7453 48311
rect 7453 48300 7455 48311
rect 7523 48311 7579 48356
rect 7523 48300 7525 48311
rect 7525 48300 7577 48311
rect 7577 48300 7579 48311
rect 7647 48311 7703 48356
rect 7647 48300 7649 48311
rect 7649 48300 7701 48311
rect 7701 48300 7703 48311
rect 7275 48176 7331 48232
rect 7399 48176 7455 48232
rect 7523 48176 7579 48232
rect 7647 48176 7703 48232
rect 7275 48052 7331 48108
rect 7399 48052 7455 48108
rect 7523 48052 7579 48108
rect 7647 48052 7703 48108
rect 7884 55692 7940 55748
rect 8008 55692 8064 55748
rect 8132 55692 8188 55748
rect 8256 55692 8312 55748
rect 8380 55692 8436 55748
rect 8504 55692 8560 55748
rect 8628 55692 8684 55748
rect 8752 55692 8808 55748
rect 8876 55692 8932 55748
rect 9000 55692 9056 55748
rect 9124 55692 9180 55748
rect 9248 55692 9304 55748
rect 9372 55692 9428 55748
rect 9496 55692 9552 55748
rect 9620 55692 9676 55748
rect 9744 55692 9800 55748
rect 7884 55568 7940 55624
rect 8008 55568 8064 55624
rect 8132 55568 8188 55624
rect 8256 55568 8312 55624
rect 8380 55568 8436 55624
rect 8504 55568 8560 55624
rect 8628 55568 8684 55624
rect 8752 55568 8808 55624
rect 8876 55568 8932 55624
rect 9000 55568 9056 55624
rect 9124 55568 9180 55624
rect 9248 55568 9304 55624
rect 9372 55568 9428 55624
rect 9496 55568 9552 55624
rect 9620 55568 9676 55624
rect 9744 55568 9800 55624
rect 7884 55444 7940 55500
rect 8008 55444 8064 55500
rect 8132 55444 8188 55500
rect 8256 55444 8312 55500
rect 8380 55444 8436 55500
rect 8504 55444 8560 55500
rect 8628 55444 8684 55500
rect 8752 55444 8808 55500
rect 8876 55444 8932 55500
rect 9000 55444 9056 55500
rect 9124 55444 9180 55500
rect 9248 55444 9304 55500
rect 9372 55444 9428 55500
rect 9496 55444 9552 55500
rect 9620 55444 9676 55500
rect 9744 55444 9800 55500
rect 7884 55320 7940 55376
rect 8008 55320 8064 55376
rect 8132 55320 8188 55376
rect 8256 55320 8312 55376
rect 8380 55320 8436 55376
rect 8504 55320 8560 55376
rect 8628 55320 8684 55376
rect 8752 55320 8808 55376
rect 8876 55320 8932 55376
rect 9000 55320 9056 55376
rect 9124 55320 9180 55376
rect 9248 55320 9304 55376
rect 9372 55320 9428 55376
rect 9496 55320 9552 55376
rect 9620 55320 9676 55376
rect 9744 55320 9800 55376
rect 7884 55196 7940 55252
rect 8008 55196 8064 55252
rect 8132 55196 8188 55252
rect 8256 55196 8312 55252
rect 8380 55196 8436 55252
rect 8504 55196 8560 55252
rect 8628 55196 8684 55252
rect 8752 55196 8808 55252
rect 8876 55196 8932 55252
rect 9000 55196 9056 55252
rect 9124 55196 9180 55252
rect 9248 55196 9304 55252
rect 9372 55196 9428 55252
rect 9496 55196 9552 55252
rect 9620 55196 9676 55252
rect 9744 55196 9800 55252
rect 7884 55072 7940 55128
rect 8008 55072 8064 55128
rect 8132 55072 8188 55128
rect 8256 55072 8312 55128
rect 8380 55072 8436 55128
rect 8504 55072 8560 55128
rect 8628 55072 8684 55128
rect 8752 55072 8808 55128
rect 8876 55072 8932 55128
rect 9000 55072 9056 55128
rect 9124 55072 9180 55128
rect 9248 55072 9304 55128
rect 9372 55072 9428 55128
rect 9496 55072 9552 55128
rect 9620 55072 9676 55128
rect 9744 55072 9800 55128
rect 7884 54948 7940 55004
rect 8008 54948 8064 55004
rect 8132 54948 8188 55004
rect 8256 54948 8312 55004
rect 8380 54948 8436 55004
rect 8504 54948 8560 55004
rect 8628 54948 8684 55004
rect 8752 54948 8808 55004
rect 8876 54948 8932 55004
rect 9000 54948 9056 55004
rect 9124 54948 9180 55004
rect 9248 54948 9304 55004
rect 9372 54948 9428 55004
rect 9496 54948 9552 55004
rect 9620 54948 9676 55004
rect 9744 54948 9800 55004
rect 7884 54824 7940 54880
rect 8008 54824 8064 54880
rect 8132 54824 8188 54880
rect 8256 54824 8312 54880
rect 8380 54824 8436 54880
rect 8504 54824 8560 54880
rect 8628 54824 8684 54880
rect 8752 54824 8808 54880
rect 8876 54824 8932 54880
rect 9000 54824 9056 54880
rect 9124 54824 9180 54880
rect 9248 54824 9304 54880
rect 9372 54824 9428 54880
rect 9496 54824 9552 54880
rect 9620 54824 9676 54880
rect 9744 54824 9800 54880
rect 7884 54700 7940 54756
rect 8008 54700 8064 54756
rect 8132 54700 8188 54756
rect 8256 54700 8312 54756
rect 8380 54700 8436 54756
rect 8504 54700 8560 54756
rect 8628 54700 8684 54756
rect 8752 54700 8808 54756
rect 8876 54700 8932 54756
rect 9000 54700 9056 54756
rect 9124 54700 9180 54756
rect 9248 54700 9304 54756
rect 9372 54700 9428 54756
rect 9496 54700 9552 54756
rect 9620 54700 9676 54756
rect 9744 54700 9800 54756
rect 7884 54576 7940 54632
rect 8008 54576 8064 54632
rect 8132 54576 8188 54632
rect 8256 54576 8312 54632
rect 8380 54576 8436 54632
rect 8504 54576 8560 54632
rect 8628 54576 8684 54632
rect 8752 54576 8808 54632
rect 8876 54576 8932 54632
rect 9000 54576 9056 54632
rect 9124 54576 9180 54632
rect 9248 54576 9304 54632
rect 9372 54576 9428 54632
rect 9496 54576 9552 54632
rect 9620 54576 9676 54632
rect 9744 54576 9800 54632
rect 7884 54452 7940 54508
rect 8008 54452 8064 54508
rect 8132 54452 8188 54508
rect 8256 54452 8312 54508
rect 8380 54452 8436 54508
rect 8504 54452 8560 54508
rect 8628 54452 8684 54508
rect 8752 54452 8808 54508
rect 8876 54452 8932 54508
rect 9000 54452 9056 54508
rect 9124 54452 9180 54508
rect 9248 54452 9304 54508
rect 9372 54452 9428 54508
rect 9496 54452 9552 54508
rect 9620 54452 9676 54508
rect 9744 54452 9800 54508
rect 7884 50892 7940 50948
rect 8008 50892 8064 50948
rect 8132 50892 8188 50948
rect 8256 50892 8312 50948
rect 8380 50892 8436 50948
rect 8504 50892 8560 50948
rect 8628 50892 8684 50948
rect 8752 50892 8808 50948
rect 8876 50892 8932 50948
rect 9000 50892 9056 50948
rect 9124 50892 9180 50948
rect 9248 50892 9304 50948
rect 9372 50892 9428 50948
rect 9496 50892 9552 50948
rect 9620 50892 9676 50948
rect 9744 50892 9800 50948
rect 7884 50768 7940 50824
rect 8008 50768 8064 50824
rect 8132 50768 8188 50824
rect 8256 50768 8312 50824
rect 8380 50768 8436 50824
rect 8504 50768 8560 50824
rect 8628 50768 8684 50824
rect 8752 50768 8808 50824
rect 8876 50768 8932 50824
rect 9000 50768 9056 50824
rect 9124 50768 9180 50824
rect 9248 50768 9304 50824
rect 9372 50768 9428 50824
rect 9496 50768 9552 50824
rect 9620 50768 9676 50824
rect 9744 50768 9800 50824
rect 7884 50693 7940 50700
rect 7884 50644 7886 50693
rect 7886 50644 7938 50693
rect 7938 50644 7940 50693
rect 8008 50693 8064 50700
rect 8008 50644 8010 50693
rect 8010 50644 8062 50693
rect 8062 50644 8064 50693
rect 8132 50693 8188 50700
rect 8132 50644 8134 50693
rect 8134 50644 8186 50693
rect 8186 50644 8188 50693
rect 8256 50693 8312 50700
rect 8256 50644 8258 50693
rect 8258 50644 8310 50693
rect 8310 50644 8312 50693
rect 8380 50693 8436 50700
rect 8380 50644 8382 50693
rect 8382 50644 8434 50693
rect 8434 50644 8436 50693
rect 8504 50693 8560 50700
rect 8504 50644 8506 50693
rect 8506 50644 8558 50693
rect 8558 50644 8560 50693
rect 8628 50693 8684 50700
rect 8628 50644 8630 50693
rect 8630 50644 8682 50693
rect 8682 50644 8684 50693
rect 8752 50693 8808 50700
rect 8752 50644 8754 50693
rect 8754 50644 8806 50693
rect 8806 50644 8808 50693
rect 8876 50693 8932 50700
rect 8876 50644 8878 50693
rect 8878 50644 8930 50693
rect 8930 50644 8932 50693
rect 9000 50693 9056 50700
rect 9000 50644 9002 50693
rect 9002 50644 9054 50693
rect 9054 50644 9056 50693
rect 9124 50693 9180 50700
rect 9124 50644 9126 50693
rect 9126 50644 9178 50693
rect 9178 50644 9180 50693
rect 9248 50693 9304 50700
rect 9248 50644 9250 50693
rect 9250 50644 9302 50693
rect 9302 50644 9304 50693
rect 9372 50693 9428 50700
rect 9372 50644 9374 50693
rect 9374 50644 9426 50693
rect 9426 50644 9428 50693
rect 9496 50693 9552 50700
rect 9496 50644 9498 50693
rect 9498 50644 9550 50693
rect 9550 50644 9552 50693
rect 9620 50693 9676 50700
rect 9620 50644 9622 50693
rect 9622 50644 9674 50693
rect 9674 50644 9676 50693
rect 9744 50693 9800 50700
rect 9744 50644 9746 50693
rect 9746 50644 9798 50693
rect 9798 50644 9800 50693
rect 7884 50569 7940 50576
rect 7884 50520 7886 50569
rect 7886 50520 7938 50569
rect 7938 50520 7940 50569
rect 8008 50569 8064 50576
rect 8008 50520 8010 50569
rect 8010 50520 8062 50569
rect 8062 50520 8064 50569
rect 8132 50569 8188 50576
rect 8132 50520 8134 50569
rect 8134 50520 8186 50569
rect 8186 50520 8188 50569
rect 8256 50569 8312 50576
rect 8256 50520 8258 50569
rect 8258 50520 8310 50569
rect 8310 50520 8312 50569
rect 8380 50569 8436 50576
rect 8380 50520 8382 50569
rect 8382 50520 8434 50569
rect 8434 50520 8436 50569
rect 8504 50569 8560 50576
rect 8504 50520 8506 50569
rect 8506 50520 8558 50569
rect 8558 50520 8560 50569
rect 8628 50569 8684 50576
rect 8628 50520 8630 50569
rect 8630 50520 8682 50569
rect 8682 50520 8684 50569
rect 8752 50569 8808 50576
rect 8752 50520 8754 50569
rect 8754 50520 8806 50569
rect 8806 50520 8808 50569
rect 8876 50569 8932 50576
rect 8876 50520 8878 50569
rect 8878 50520 8930 50569
rect 8930 50520 8932 50569
rect 9000 50569 9056 50576
rect 9000 50520 9002 50569
rect 9002 50520 9054 50569
rect 9054 50520 9056 50569
rect 9124 50569 9180 50576
rect 9124 50520 9126 50569
rect 9126 50520 9178 50569
rect 9178 50520 9180 50569
rect 9248 50569 9304 50576
rect 9248 50520 9250 50569
rect 9250 50520 9302 50569
rect 9302 50520 9304 50569
rect 9372 50569 9428 50576
rect 9372 50520 9374 50569
rect 9374 50520 9426 50569
rect 9426 50520 9428 50569
rect 9496 50569 9552 50576
rect 9496 50520 9498 50569
rect 9498 50520 9550 50569
rect 9550 50520 9552 50569
rect 9620 50569 9676 50576
rect 9620 50520 9622 50569
rect 9622 50520 9674 50569
rect 9674 50520 9676 50569
rect 9744 50569 9800 50576
rect 9744 50520 9746 50569
rect 9746 50520 9798 50569
rect 9798 50520 9800 50569
rect 7884 50396 7940 50452
rect 8008 50396 8064 50452
rect 8132 50396 8188 50452
rect 8256 50396 8312 50452
rect 8380 50396 8436 50452
rect 8504 50396 8560 50452
rect 8628 50396 8684 50452
rect 8752 50396 8808 50452
rect 8876 50396 8932 50452
rect 9000 50396 9056 50452
rect 9124 50396 9180 50452
rect 9248 50396 9304 50452
rect 9372 50396 9428 50452
rect 9496 50396 9552 50452
rect 9620 50396 9676 50452
rect 9744 50396 9800 50452
rect 7884 50272 7940 50328
rect 8008 50272 8064 50328
rect 8132 50272 8188 50328
rect 8256 50272 8312 50328
rect 8380 50272 8436 50328
rect 8504 50272 8560 50328
rect 8628 50272 8684 50328
rect 8752 50272 8808 50328
rect 8876 50272 8932 50328
rect 9000 50272 9056 50328
rect 9124 50272 9180 50328
rect 9248 50272 9304 50328
rect 9372 50272 9428 50328
rect 9496 50272 9552 50328
rect 9620 50272 9676 50328
rect 9744 50272 9800 50328
rect 7884 50148 7940 50204
rect 8008 50148 8064 50204
rect 8132 50148 8188 50204
rect 8256 50148 8312 50204
rect 8380 50148 8436 50204
rect 8504 50148 8560 50204
rect 8628 50148 8684 50204
rect 8752 50148 8808 50204
rect 8876 50148 8932 50204
rect 9000 50148 9056 50204
rect 9124 50148 9180 50204
rect 9248 50148 9304 50204
rect 9372 50148 9428 50204
rect 9496 50148 9552 50204
rect 9620 50148 9676 50204
rect 9744 50148 9800 50204
rect 7884 50024 7940 50080
rect 8008 50024 8064 50080
rect 8132 50024 8188 50080
rect 8256 50024 8312 50080
rect 8380 50024 8436 50080
rect 8504 50024 8560 50080
rect 8628 50024 8684 50080
rect 8752 50024 8808 50080
rect 8876 50024 8932 50080
rect 9000 50024 9056 50080
rect 9124 50024 9180 50080
rect 9248 50024 9304 50080
rect 9372 50024 9428 50080
rect 9496 50024 9552 50080
rect 9620 50024 9676 50080
rect 9744 50024 9800 50080
rect 7884 49900 7940 49956
rect 8008 49900 8064 49956
rect 8132 49900 8188 49956
rect 8256 49900 8312 49956
rect 8380 49900 8436 49956
rect 8504 49900 8560 49956
rect 8628 49900 8684 49956
rect 8752 49900 8808 49956
rect 8876 49900 8932 49956
rect 9000 49900 9056 49956
rect 9124 49900 9180 49956
rect 9248 49900 9304 49956
rect 9372 49900 9428 49956
rect 9496 49900 9552 49956
rect 9620 49900 9676 49956
rect 9744 49900 9800 49956
rect 7884 49776 7940 49832
rect 8008 49776 8064 49832
rect 8132 49776 8188 49832
rect 8256 49776 8312 49832
rect 8380 49776 8436 49832
rect 8504 49776 8560 49832
rect 8628 49776 8684 49832
rect 8752 49776 8808 49832
rect 8876 49776 8932 49832
rect 9000 49776 9056 49832
rect 9124 49776 9180 49832
rect 9248 49776 9304 49832
rect 9372 49776 9428 49832
rect 9496 49776 9552 49832
rect 9620 49776 9676 49832
rect 9744 49776 9800 49832
rect 7884 49707 7886 49708
rect 7886 49707 7938 49708
rect 7938 49707 7940 49708
rect 7884 49652 7940 49707
rect 8008 49707 8010 49708
rect 8010 49707 8062 49708
rect 8062 49707 8064 49708
rect 8008 49652 8064 49707
rect 8132 49707 8134 49708
rect 8134 49707 8186 49708
rect 8186 49707 8188 49708
rect 8132 49652 8188 49707
rect 8256 49707 8258 49708
rect 8258 49707 8310 49708
rect 8310 49707 8312 49708
rect 8256 49652 8312 49707
rect 8380 49707 8382 49708
rect 8382 49707 8434 49708
rect 8434 49707 8436 49708
rect 8380 49652 8436 49707
rect 8504 49707 8506 49708
rect 8506 49707 8558 49708
rect 8558 49707 8560 49708
rect 8504 49652 8560 49707
rect 8628 49707 8630 49708
rect 8630 49707 8682 49708
rect 8682 49707 8684 49708
rect 8628 49652 8684 49707
rect 8752 49707 8754 49708
rect 8754 49707 8806 49708
rect 8806 49707 8808 49708
rect 8752 49652 8808 49707
rect 8876 49707 8878 49708
rect 8878 49707 8930 49708
rect 8930 49707 8932 49708
rect 8876 49652 8932 49707
rect 9000 49707 9002 49708
rect 9002 49707 9054 49708
rect 9054 49707 9056 49708
rect 9000 49652 9056 49707
rect 9124 49707 9126 49708
rect 9126 49707 9178 49708
rect 9178 49707 9180 49708
rect 9124 49652 9180 49707
rect 9248 49707 9250 49708
rect 9250 49707 9302 49708
rect 9302 49707 9304 49708
rect 9248 49652 9304 49707
rect 9372 49707 9374 49708
rect 9374 49707 9426 49708
rect 9426 49707 9428 49708
rect 9372 49652 9428 49707
rect 9496 49707 9498 49708
rect 9498 49707 9550 49708
rect 9550 49707 9552 49708
rect 9496 49652 9552 49707
rect 9620 49707 9622 49708
rect 9622 49707 9674 49708
rect 9674 49707 9676 49708
rect 9620 49652 9676 49707
rect 9744 49707 9746 49708
rect 9746 49707 9798 49708
rect 9798 49707 9800 49708
rect 9744 49652 9800 49707
rect 7884 47740 7940 47748
rect 7884 47692 7886 47740
rect 7886 47692 7938 47740
rect 7938 47692 7940 47740
rect 8008 47740 8064 47748
rect 8008 47692 8010 47740
rect 8010 47692 8062 47740
rect 8062 47692 8064 47740
rect 8132 47740 8188 47748
rect 8132 47692 8134 47740
rect 8134 47692 8186 47740
rect 8186 47692 8188 47740
rect 8256 47740 8312 47748
rect 8256 47692 8258 47740
rect 8258 47692 8310 47740
rect 8310 47692 8312 47740
rect 8380 47740 8436 47748
rect 8380 47692 8382 47740
rect 8382 47692 8434 47740
rect 8434 47692 8436 47740
rect 8504 47740 8560 47748
rect 8504 47692 8506 47740
rect 8506 47692 8558 47740
rect 8558 47692 8560 47740
rect 8628 47740 8684 47748
rect 8628 47692 8630 47740
rect 8630 47692 8682 47740
rect 8682 47692 8684 47740
rect 8752 47740 8808 47748
rect 8752 47692 8754 47740
rect 8754 47692 8806 47740
rect 8806 47692 8808 47740
rect 8876 47740 8932 47748
rect 8876 47692 8878 47740
rect 8878 47692 8930 47740
rect 8930 47692 8932 47740
rect 9000 47740 9056 47748
rect 9000 47692 9002 47740
rect 9002 47692 9054 47740
rect 9054 47692 9056 47740
rect 9124 47740 9180 47748
rect 9124 47692 9126 47740
rect 9126 47692 9178 47740
rect 9178 47692 9180 47740
rect 9248 47740 9304 47748
rect 9248 47692 9250 47740
rect 9250 47692 9302 47740
rect 9302 47692 9304 47740
rect 9372 47740 9428 47748
rect 9372 47692 9374 47740
rect 9374 47692 9426 47740
rect 9426 47692 9428 47740
rect 9496 47740 9552 47748
rect 9496 47692 9498 47740
rect 9498 47692 9550 47740
rect 9550 47692 9552 47740
rect 9620 47740 9676 47748
rect 9620 47692 9622 47740
rect 9622 47692 9674 47740
rect 9674 47692 9676 47740
rect 9744 47740 9800 47748
rect 9744 47692 9746 47740
rect 9746 47692 9798 47740
rect 9798 47692 9800 47740
rect 7884 47568 7940 47624
rect 8008 47568 8064 47624
rect 8132 47568 8188 47624
rect 8256 47568 8312 47624
rect 8380 47568 8436 47624
rect 8504 47568 8560 47624
rect 8628 47568 8684 47624
rect 8752 47568 8808 47624
rect 8876 47568 8932 47624
rect 9000 47568 9056 47624
rect 9124 47568 9180 47624
rect 9248 47568 9304 47624
rect 9372 47568 9428 47624
rect 9496 47568 9552 47624
rect 9620 47568 9676 47624
rect 9744 47568 9800 47624
rect 7884 47444 7940 47500
rect 8008 47444 8064 47500
rect 8132 47444 8188 47500
rect 8256 47444 8312 47500
rect 8380 47444 8436 47500
rect 8504 47444 8560 47500
rect 8628 47444 8684 47500
rect 8752 47444 8808 47500
rect 8876 47444 8932 47500
rect 9000 47444 9056 47500
rect 9124 47444 9180 47500
rect 9248 47444 9304 47500
rect 9372 47444 9428 47500
rect 9496 47444 9552 47500
rect 9620 47444 9676 47500
rect 9744 47444 9800 47500
rect 7884 47320 7940 47376
rect 8008 47320 8064 47376
rect 8132 47320 8188 47376
rect 8256 47320 8312 47376
rect 8380 47320 8436 47376
rect 8504 47320 8560 47376
rect 8628 47320 8684 47376
rect 8752 47320 8808 47376
rect 8876 47320 8932 47376
rect 9000 47320 9056 47376
rect 9124 47320 9180 47376
rect 9248 47320 9304 47376
rect 9372 47320 9428 47376
rect 9496 47320 9552 47376
rect 9620 47320 9676 47376
rect 9744 47320 9800 47376
rect 9937 57169 9993 57225
rect 10061 57169 10117 57225
rect 9937 57056 9947 57101
rect 9947 57056 9993 57101
rect 10061 57056 10107 57101
rect 10107 57056 10117 57101
rect 9937 57045 9993 57056
rect 10061 57045 10117 57056
rect 9937 56921 9993 56977
rect 10061 56921 10117 56977
rect 9937 56797 9993 56853
rect 10061 56797 10117 56853
rect 9937 56673 9993 56729
rect 10061 56673 10117 56729
rect 9937 56549 9993 56605
rect 10061 56549 10117 56605
rect 9937 56425 9993 56481
rect 10061 56425 10117 56481
rect 9937 56301 9993 56357
rect 10061 56301 10117 56357
rect 9937 56177 9993 56233
rect 10061 56177 10117 56233
rect 9937 56053 9993 56109
rect 10061 56053 10117 56109
rect 9937 54092 9993 54148
rect 10061 54092 10117 54148
rect 9937 53968 9993 54024
rect 10061 53968 10117 54024
rect 9937 53844 9993 53900
rect 10061 53844 10117 53900
rect 9937 53720 9993 53776
rect 10061 53720 10117 53776
rect 9937 53596 9993 53652
rect 10061 53596 10117 53652
rect 9937 53484 9993 53528
rect 10061 53484 10117 53528
rect 9937 53472 9947 53484
rect 9947 53472 9993 53484
rect 10061 53472 10107 53484
rect 10107 53472 10117 53484
rect 9937 53376 9993 53404
rect 10061 53376 10117 53404
rect 9937 53348 9947 53376
rect 9947 53348 9993 53376
rect 10061 53348 10107 53376
rect 10107 53348 10117 53376
rect 9937 53268 9993 53280
rect 10061 53268 10117 53280
rect 9937 53224 9947 53268
rect 9947 53224 9993 53268
rect 10061 53224 10107 53268
rect 10107 53224 10117 53268
rect 9937 53100 9993 53156
rect 10061 53100 10117 53156
rect 9937 52976 9993 53032
rect 10061 52976 10117 53032
rect 9937 52852 9993 52908
rect 10061 52852 10117 52908
rect 9937 49302 9939 49348
rect 9939 49302 9991 49348
rect 9991 49302 9993 49348
rect 9937 49292 9993 49302
rect 10061 49302 10063 49348
rect 10063 49302 10115 49348
rect 10115 49302 10117 49348
rect 10061 49292 10117 49302
rect 9937 49178 9939 49224
rect 9939 49178 9991 49224
rect 9991 49178 9993 49224
rect 9937 49168 9993 49178
rect 10061 49178 10063 49224
rect 10063 49178 10115 49224
rect 10115 49178 10117 49224
rect 10061 49168 10117 49178
rect 9937 49054 9939 49100
rect 9939 49054 9991 49100
rect 9991 49054 9993 49100
rect 9937 49044 9993 49054
rect 10061 49054 10063 49100
rect 10063 49054 10115 49100
rect 10115 49054 10117 49100
rect 10061 49044 10117 49054
rect 9937 48920 9993 48976
rect 10061 48920 10117 48976
rect 9937 48796 9993 48852
rect 10061 48796 10117 48852
rect 9937 48672 9993 48728
rect 10061 48672 10117 48728
rect 9937 48548 9993 48604
rect 10061 48548 10117 48604
rect 9937 48435 9993 48480
rect 9937 48424 9939 48435
rect 9939 48424 9991 48435
rect 9991 48424 9993 48435
rect 10061 48435 10117 48480
rect 10061 48424 10063 48435
rect 10063 48424 10115 48435
rect 10115 48424 10117 48435
rect 9937 48311 9993 48356
rect 9937 48300 9939 48311
rect 9939 48300 9991 48311
rect 9991 48300 9993 48311
rect 10061 48311 10117 48356
rect 10061 48300 10063 48311
rect 10063 48300 10115 48311
rect 10115 48300 10117 48311
rect 9937 48176 9993 48232
rect 10061 48176 10117 48232
rect 9937 48052 9993 48108
rect 10061 48052 10117 48108
rect 10254 55692 10310 55748
rect 10378 55692 10434 55748
rect 10502 55692 10558 55748
rect 10626 55692 10682 55748
rect 10750 55692 10806 55748
rect 10874 55692 10930 55748
rect 10998 55692 11054 55748
rect 11122 55692 11178 55748
rect 11246 55692 11302 55748
rect 11370 55692 11426 55748
rect 11494 55692 11550 55748
rect 11618 55692 11674 55748
rect 11742 55692 11798 55748
rect 11866 55692 11922 55748
rect 11990 55692 12046 55748
rect 12114 55692 12170 55748
rect 10254 55568 10310 55624
rect 10378 55568 10434 55624
rect 10502 55568 10558 55624
rect 10626 55568 10682 55624
rect 10750 55568 10806 55624
rect 10874 55568 10930 55624
rect 10998 55568 11054 55624
rect 11122 55568 11178 55624
rect 11246 55568 11302 55624
rect 11370 55568 11426 55624
rect 11494 55568 11550 55624
rect 11618 55568 11674 55624
rect 11742 55568 11798 55624
rect 11866 55568 11922 55624
rect 11990 55568 12046 55624
rect 12114 55568 12170 55624
rect 10254 55444 10310 55500
rect 10378 55444 10434 55500
rect 10502 55444 10558 55500
rect 10626 55444 10682 55500
rect 10750 55444 10806 55500
rect 10874 55444 10930 55500
rect 10998 55444 11054 55500
rect 11122 55444 11178 55500
rect 11246 55444 11302 55500
rect 11370 55444 11426 55500
rect 11494 55444 11550 55500
rect 11618 55444 11674 55500
rect 11742 55444 11798 55500
rect 11866 55444 11922 55500
rect 11990 55444 12046 55500
rect 12114 55444 12170 55500
rect 10254 55320 10310 55376
rect 10378 55320 10434 55376
rect 10502 55320 10558 55376
rect 10626 55320 10682 55376
rect 10750 55320 10806 55376
rect 10874 55320 10930 55376
rect 10998 55320 11054 55376
rect 11122 55320 11178 55376
rect 11246 55320 11302 55376
rect 11370 55320 11426 55376
rect 11494 55320 11550 55376
rect 11618 55320 11674 55376
rect 11742 55320 11798 55376
rect 11866 55320 11922 55376
rect 11990 55320 12046 55376
rect 12114 55320 12170 55376
rect 10254 55196 10310 55252
rect 10378 55196 10434 55252
rect 10502 55196 10558 55252
rect 10626 55196 10682 55252
rect 10750 55196 10806 55252
rect 10874 55196 10930 55252
rect 10998 55196 11054 55252
rect 11122 55196 11178 55252
rect 11246 55196 11302 55252
rect 11370 55196 11426 55252
rect 11494 55196 11550 55252
rect 11618 55196 11674 55252
rect 11742 55196 11798 55252
rect 11866 55196 11922 55252
rect 11990 55196 12046 55252
rect 12114 55196 12170 55252
rect 10254 55072 10310 55128
rect 10378 55072 10434 55128
rect 10502 55072 10558 55128
rect 10626 55072 10682 55128
rect 10750 55072 10806 55128
rect 10874 55072 10930 55128
rect 10998 55072 11054 55128
rect 11122 55072 11178 55128
rect 11246 55072 11302 55128
rect 11370 55072 11426 55128
rect 11494 55072 11550 55128
rect 11618 55072 11674 55128
rect 11742 55072 11798 55128
rect 11866 55072 11922 55128
rect 11990 55072 12046 55128
rect 12114 55072 12170 55128
rect 10254 54948 10310 55004
rect 10378 54948 10434 55004
rect 10502 54948 10558 55004
rect 10626 54948 10682 55004
rect 10750 54948 10806 55004
rect 10874 54948 10930 55004
rect 10998 54948 11054 55004
rect 11122 54948 11178 55004
rect 11246 54948 11302 55004
rect 11370 54948 11426 55004
rect 11494 54948 11550 55004
rect 11618 54948 11674 55004
rect 11742 54948 11798 55004
rect 11866 54948 11922 55004
rect 11990 54948 12046 55004
rect 12114 54948 12170 55004
rect 10254 54824 10310 54880
rect 10378 54824 10434 54880
rect 10502 54824 10558 54880
rect 10626 54824 10682 54880
rect 10750 54824 10806 54880
rect 10874 54824 10930 54880
rect 10998 54824 11054 54880
rect 11122 54824 11178 54880
rect 11246 54824 11302 54880
rect 11370 54824 11426 54880
rect 11494 54824 11550 54880
rect 11618 54824 11674 54880
rect 11742 54824 11798 54880
rect 11866 54824 11922 54880
rect 11990 54824 12046 54880
rect 12114 54824 12170 54880
rect 10254 54700 10310 54756
rect 10378 54700 10434 54756
rect 10502 54700 10558 54756
rect 10626 54700 10682 54756
rect 10750 54700 10806 54756
rect 10874 54700 10930 54756
rect 10998 54700 11054 54756
rect 11122 54700 11178 54756
rect 11246 54700 11302 54756
rect 11370 54700 11426 54756
rect 11494 54700 11550 54756
rect 11618 54700 11674 54756
rect 11742 54700 11798 54756
rect 11866 54700 11922 54756
rect 11990 54700 12046 54756
rect 12114 54700 12170 54756
rect 10254 54576 10310 54632
rect 10378 54576 10434 54632
rect 10502 54576 10558 54632
rect 10626 54576 10682 54632
rect 10750 54576 10806 54632
rect 10874 54576 10930 54632
rect 10998 54576 11054 54632
rect 11122 54576 11178 54632
rect 11246 54576 11302 54632
rect 11370 54576 11426 54632
rect 11494 54576 11550 54632
rect 11618 54576 11674 54632
rect 11742 54576 11798 54632
rect 11866 54576 11922 54632
rect 11990 54576 12046 54632
rect 12114 54576 12170 54632
rect 10254 54452 10310 54508
rect 10378 54452 10434 54508
rect 10502 54452 10558 54508
rect 10626 54452 10682 54508
rect 10750 54452 10806 54508
rect 10874 54452 10930 54508
rect 10998 54452 11054 54508
rect 11122 54452 11178 54508
rect 11246 54452 11302 54508
rect 11370 54452 11426 54508
rect 11494 54452 11550 54508
rect 11618 54452 11674 54508
rect 11742 54452 11798 54508
rect 11866 54452 11922 54508
rect 11990 54452 12046 54508
rect 12114 54452 12170 54508
rect 10254 50892 10310 50948
rect 10378 50892 10434 50948
rect 10502 50892 10558 50948
rect 10626 50892 10682 50948
rect 10750 50892 10806 50948
rect 10874 50892 10930 50948
rect 10998 50892 11054 50948
rect 11122 50892 11178 50948
rect 11246 50892 11302 50948
rect 11370 50892 11426 50948
rect 11494 50892 11550 50948
rect 11618 50892 11674 50948
rect 11742 50892 11798 50948
rect 11866 50892 11922 50948
rect 11990 50892 12046 50948
rect 12114 50892 12170 50948
rect 10254 50768 10310 50824
rect 10378 50768 10434 50824
rect 10502 50768 10558 50824
rect 10626 50768 10682 50824
rect 10750 50768 10806 50824
rect 10874 50768 10930 50824
rect 10998 50768 11054 50824
rect 11122 50768 11178 50824
rect 11246 50768 11302 50824
rect 11370 50768 11426 50824
rect 11494 50768 11550 50824
rect 11618 50768 11674 50824
rect 11742 50768 11798 50824
rect 11866 50768 11922 50824
rect 11990 50768 12046 50824
rect 12114 50768 12170 50824
rect 10254 50693 10310 50700
rect 10378 50693 10434 50700
rect 10502 50693 10558 50700
rect 10626 50693 10682 50700
rect 10750 50693 10806 50700
rect 10874 50693 10930 50700
rect 10998 50693 11054 50700
rect 11122 50693 11178 50700
rect 11246 50693 11302 50700
rect 11370 50693 11426 50700
rect 10254 50644 10303 50693
rect 10303 50644 10310 50693
rect 10378 50644 10427 50693
rect 10427 50644 10434 50693
rect 10502 50644 10551 50693
rect 10551 50644 10558 50693
rect 10626 50644 10675 50693
rect 10675 50644 10682 50693
rect 10750 50644 10799 50693
rect 10799 50644 10806 50693
rect 10874 50644 10923 50693
rect 10923 50644 10930 50693
rect 10998 50644 11047 50693
rect 11047 50644 11054 50693
rect 11122 50644 11171 50693
rect 11171 50644 11178 50693
rect 11246 50644 11295 50693
rect 11295 50644 11302 50693
rect 11370 50644 11419 50693
rect 11419 50644 11426 50693
rect 11494 50644 11550 50700
rect 11618 50644 11674 50700
rect 11742 50644 11798 50700
rect 11866 50644 11922 50700
rect 11990 50644 12046 50700
rect 12114 50644 12170 50700
rect 10254 50569 10310 50576
rect 10378 50569 10434 50576
rect 10502 50569 10558 50576
rect 10626 50569 10682 50576
rect 10750 50569 10806 50576
rect 10874 50569 10930 50576
rect 10998 50569 11054 50576
rect 11122 50569 11178 50576
rect 11246 50569 11302 50576
rect 11370 50569 11426 50576
rect 10254 50520 10303 50569
rect 10303 50520 10310 50569
rect 10378 50520 10427 50569
rect 10427 50520 10434 50569
rect 10502 50520 10551 50569
rect 10551 50520 10558 50569
rect 10626 50520 10675 50569
rect 10675 50520 10682 50569
rect 10750 50520 10799 50569
rect 10799 50520 10806 50569
rect 10874 50520 10923 50569
rect 10923 50520 10930 50569
rect 10998 50520 11047 50569
rect 11047 50520 11054 50569
rect 11122 50520 11171 50569
rect 11171 50520 11178 50569
rect 11246 50520 11295 50569
rect 11295 50520 11302 50569
rect 11370 50520 11419 50569
rect 11419 50520 11426 50569
rect 11494 50520 11550 50576
rect 11618 50520 11674 50576
rect 11742 50520 11798 50576
rect 11866 50520 11922 50576
rect 11990 50520 12046 50576
rect 12114 50520 12170 50576
rect 10254 50396 10310 50452
rect 10378 50396 10434 50452
rect 10502 50396 10558 50452
rect 10626 50396 10682 50452
rect 10750 50396 10806 50452
rect 10874 50396 10930 50452
rect 10998 50396 11054 50452
rect 11122 50396 11178 50452
rect 11246 50396 11302 50452
rect 11370 50396 11426 50452
rect 11494 50396 11550 50452
rect 11618 50396 11674 50452
rect 11742 50396 11798 50452
rect 11866 50396 11922 50452
rect 11990 50396 12046 50452
rect 12114 50396 12170 50452
rect 10254 50272 10310 50328
rect 10378 50272 10434 50328
rect 10502 50272 10558 50328
rect 10626 50272 10682 50328
rect 10750 50272 10806 50328
rect 10874 50272 10930 50328
rect 10998 50272 11054 50328
rect 11122 50272 11178 50328
rect 11246 50272 11302 50328
rect 11370 50272 11426 50328
rect 11494 50272 11550 50328
rect 11618 50272 11674 50328
rect 11742 50272 11798 50328
rect 11866 50272 11922 50328
rect 11990 50272 12046 50328
rect 12114 50272 12170 50328
rect 10254 50148 10310 50204
rect 10378 50148 10434 50204
rect 10502 50148 10558 50204
rect 10626 50148 10682 50204
rect 10750 50148 10806 50204
rect 10874 50148 10930 50204
rect 10998 50148 11054 50204
rect 11122 50148 11178 50204
rect 11246 50148 11302 50204
rect 11370 50148 11426 50204
rect 11494 50148 11550 50204
rect 11618 50148 11674 50204
rect 11742 50148 11798 50204
rect 11866 50148 11922 50204
rect 11990 50148 12046 50204
rect 12114 50148 12170 50204
rect 10254 50024 10310 50080
rect 10378 50024 10434 50080
rect 10502 50024 10558 50080
rect 10626 50024 10682 50080
rect 10750 50024 10806 50080
rect 10874 50024 10930 50080
rect 10998 50024 11054 50080
rect 11122 50024 11178 50080
rect 11246 50024 11302 50080
rect 11370 50024 11426 50080
rect 11494 50024 11550 50080
rect 11618 50024 11674 50080
rect 11742 50024 11798 50080
rect 11866 50024 11922 50080
rect 11990 50024 12046 50080
rect 12114 50024 12170 50080
rect 10254 49900 10310 49956
rect 10378 49900 10434 49956
rect 10502 49900 10558 49956
rect 10626 49900 10682 49956
rect 10750 49900 10806 49956
rect 10874 49900 10930 49956
rect 10998 49900 11054 49956
rect 11122 49900 11178 49956
rect 11246 49900 11302 49956
rect 11370 49900 11426 49956
rect 11494 49900 11550 49956
rect 11618 49900 11674 49956
rect 11742 49900 11798 49956
rect 11866 49900 11922 49956
rect 11990 49900 12046 49956
rect 12114 49900 12170 49956
rect 10254 49776 10310 49832
rect 10378 49776 10434 49832
rect 10502 49776 10558 49832
rect 10626 49776 10682 49832
rect 10750 49776 10806 49832
rect 10874 49776 10930 49832
rect 10998 49776 11054 49832
rect 11122 49776 11178 49832
rect 11246 49776 11302 49832
rect 11370 49776 11426 49832
rect 11494 49776 11550 49832
rect 11618 49776 11674 49832
rect 11742 49776 11798 49832
rect 11866 49776 11922 49832
rect 11990 49776 12046 49832
rect 12114 49776 12170 49832
rect 10254 49707 10303 49708
rect 10303 49707 10310 49708
rect 10378 49707 10427 49708
rect 10427 49707 10434 49708
rect 10502 49707 10551 49708
rect 10551 49707 10558 49708
rect 10626 49707 10675 49708
rect 10675 49707 10682 49708
rect 10750 49707 10799 49708
rect 10799 49707 10806 49708
rect 10874 49707 10923 49708
rect 10923 49707 10930 49708
rect 10998 49707 11047 49708
rect 11047 49707 11054 49708
rect 11122 49707 11171 49708
rect 11171 49707 11178 49708
rect 11246 49707 11295 49708
rect 11295 49707 11302 49708
rect 11370 49707 11419 49708
rect 11419 49707 11426 49708
rect 10254 49652 10310 49707
rect 10378 49652 10434 49707
rect 10502 49652 10558 49707
rect 10626 49652 10682 49707
rect 10750 49652 10806 49707
rect 10874 49652 10930 49707
rect 10998 49652 11054 49707
rect 11122 49652 11178 49707
rect 11246 49652 11302 49707
rect 11370 49652 11426 49707
rect 11494 49652 11550 49708
rect 11618 49652 11674 49708
rect 11742 49652 11798 49708
rect 11866 49652 11922 49708
rect 11990 49652 12046 49708
rect 12114 49652 12170 49708
rect 10254 47740 10310 47748
rect 10254 47692 10256 47740
rect 10256 47692 10308 47740
rect 10308 47692 10310 47740
rect 10378 47740 10434 47748
rect 10378 47692 10380 47740
rect 10380 47692 10432 47740
rect 10432 47692 10434 47740
rect 10502 47740 10558 47748
rect 10502 47692 10504 47740
rect 10504 47692 10556 47740
rect 10556 47692 10558 47740
rect 10626 47740 10682 47748
rect 10626 47692 10628 47740
rect 10628 47692 10680 47740
rect 10680 47692 10682 47740
rect 10750 47740 10806 47748
rect 10750 47692 10752 47740
rect 10752 47692 10804 47740
rect 10804 47692 10806 47740
rect 10874 47740 10930 47748
rect 10874 47692 10876 47740
rect 10876 47692 10928 47740
rect 10928 47692 10930 47740
rect 10998 47740 11054 47748
rect 10998 47692 11000 47740
rect 11000 47692 11052 47740
rect 11052 47692 11054 47740
rect 11122 47740 11178 47748
rect 11122 47692 11124 47740
rect 11124 47692 11176 47740
rect 11176 47692 11178 47740
rect 11246 47740 11302 47748
rect 11246 47692 11248 47740
rect 11248 47692 11300 47740
rect 11300 47692 11302 47740
rect 11370 47740 11426 47748
rect 11370 47692 11372 47740
rect 11372 47692 11424 47740
rect 11424 47692 11426 47740
rect 11494 47740 11550 47748
rect 11494 47692 11496 47740
rect 11496 47692 11548 47740
rect 11548 47692 11550 47740
rect 11618 47740 11674 47748
rect 11618 47692 11620 47740
rect 11620 47692 11672 47740
rect 11672 47692 11674 47740
rect 11742 47740 11798 47748
rect 11742 47692 11744 47740
rect 11744 47692 11796 47740
rect 11796 47692 11798 47740
rect 11866 47740 11922 47748
rect 11866 47692 11868 47740
rect 11868 47692 11920 47740
rect 11920 47692 11922 47740
rect 11990 47740 12046 47748
rect 11990 47692 11992 47740
rect 11992 47692 12044 47740
rect 12044 47692 12046 47740
rect 12114 47740 12170 47748
rect 12114 47692 12116 47740
rect 12116 47692 12168 47740
rect 12168 47692 12170 47740
rect 10254 47568 10310 47624
rect 10378 47568 10434 47624
rect 10502 47568 10558 47624
rect 10626 47568 10682 47624
rect 10750 47568 10806 47624
rect 10874 47568 10930 47624
rect 10998 47568 11054 47624
rect 11122 47568 11178 47624
rect 11246 47568 11302 47624
rect 11370 47568 11426 47624
rect 11494 47568 11550 47624
rect 11618 47568 11674 47624
rect 11742 47568 11798 47624
rect 11866 47568 11922 47624
rect 11990 47568 12046 47624
rect 12114 47568 12170 47624
rect 10254 47444 10310 47500
rect 10378 47444 10434 47500
rect 10502 47444 10558 47500
rect 10626 47444 10682 47500
rect 10750 47444 10806 47500
rect 10874 47444 10930 47500
rect 10998 47444 11054 47500
rect 11122 47444 11178 47500
rect 11246 47444 11302 47500
rect 11370 47444 11426 47500
rect 11494 47444 11550 47500
rect 11618 47444 11674 47500
rect 11742 47444 11798 47500
rect 11866 47444 11922 47500
rect 11990 47444 12046 47500
rect 12114 47444 12170 47500
rect 10254 47320 10310 47376
rect 10378 47320 10434 47376
rect 10502 47320 10558 47376
rect 10626 47320 10682 47376
rect 10750 47320 10806 47376
rect 10874 47320 10930 47376
rect 10998 47320 11054 47376
rect 11122 47320 11178 47376
rect 11246 47320 11302 47376
rect 11370 47320 11426 47376
rect 11494 47320 11550 47376
rect 11618 47320 11674 47376
rect 11742 47320 11798 47376
rect 11866 47320 11922 47376
rect 11990 47320 12046 47376
rect 12114 47320 12170 47376
rect 12307 57169 12363 57225
rect 12431 57169 12487 57225
rect 12307 57056 12317 57101
rect 12317 57056 12363 57101
rect 12431 57056 12477 57101
rect 12477 57056 12487 57101
rect 12307 57045 12363 57056
rect 12431 57045 12487 57056
rect 12307 56921 12363 56977
rect 12431 56921 12487 56977
rect 12307 56797 12363 56853
rect 12431 56797 12487 56853
rect 12307 56673 12363 56729
rect 12431 56673 12487 56729
rect 12307 56549 12363 56605
rect 12431 56549 12487 56605
rect 12307 56425 12363 56481
rect 12431 56425 12487 56481
rect 12307 56301 12363 56357
rect 12431 56301 12487 56357
rect 12307 56177 12363 56233
rect 12431 56177 12487 56233
rect 12307 56053 12363 56109
rect 12431 56053 12487 56109
rect 12307 54092 12363 54148
rect 12431 54092 12487 54148
rect 12307 53968 12363 54024
rect 12431 53968 12487 54024
rect 12307 53844 12363 53900
rect 12431 53844 12487 53900
rect 12307 53720 12363 53776
rect 12431 53720 12487 53776
rect 12307 53596 12363 53652
rect 12431 53596 12487 53652
rect 12307 53484 12363 53528
rect 12431 53484 12487 53528
rect 12307 53472 12317 53484
rect 12317 53472 12363 53484
rect 12431 53472 12477 53484
rect 12477 53472 12487 53484
rect 12307 53376 12363 53404
rect 12431 53376 12487 53404
rect 12307 53348 12317 53376
rect 12317 53348 12363 53376
rect 12431 53348 12477 53376
rect 12477 53348 12487 53376
rect 12307 53268 12363 53280
rect 12431 53268 12487 53280
rect 12307 53224 12317 53268
rect 12317 53224 12363 53268
rect 12431 53224 12477 53268
rect 12477 53224 12487 53268
rect 12307 53100 12363 53156
rect 12431 53100 12487 53156
rect 12307 52976 12363 53032
rect 12431 52976 12487 53032
rect 12307 52852 12363 52908
rect 12431 52852 12487 52908
rect 12307 49292 12363 49348
rect 12431 49292 12487 49348
rect 12307 49168 12363 49224
rect 12431 49168 12487 49224
rect 12307 49044 12363 49100
rect 12431 49044 12487 49100
rect 12307 48920 12363 48976
rect 12431 48920 12487 48976
rect 12307 48796 12363 48852
rect 12431 48796 12487 48852
rect 12307 48672 12363 48728
rect 12431 48672 12487 48728
rect 12307 48548 12363 48604
rect 12431 48548 12487 48604
rect 12307 48424 12363 48480
rect 12431 48424 12487 48480
rect 12307 48300 12363 48356
rect 12431 48300 12487 48356
rect 12307 48176 12363 48232
rect 12431 48176 12487 48232
rect 12307 48052 12363 48108
rect 12431 48052 12487 48108
rect 12871 55692 12927 55748
rect 12995 55692 13051 55748
rect 13119 55692 13175 55748
rect 13243 55692 13299 55748
rect 13367 55692 13423 55748
rect 13491 55692 13547 55748
rect 13615 55692 13671 55748
rect 13739 55692 13795 55748
rect 13863 55692 13919 55748
rect 13987 55692 14043 55748
rect 14111 55692 14167 55748
rect 14235 55692 14291 55748
rect 14359 55692 14415 55748
rect 14483 55692 14539 55748
rect 14607 55692 14663 55748
rect 12871 55568 12927 55624
rect 12995 55568 13051 55624
rect 13119 55568 13175 55624
rect 13243 55568 13299 55624
rect 13367 55568 13423 55624
rect 13491 55568 13547 55624
rect 13615 55568 13671 55624
rect 13739 55568 13795 55624
rect 13863 55568 13919 55624
rect 13987 55568 14043 55624
rect 14111 55568 14167 55624
rect 14235 55568 14291 55624
rect 14359 55568 14415 55624
rect 14483 55568 14539 55624
rect 14607 55568 14663 55624
rect 12871 55444 12927 55500
rect 12995 55444 13051 55500
rect 13119 55444 13175 55500
rect 13243 55444 13299 55500
rect 13367 55444 13423 55500
rect 13491 55444 13547 55500
rect 13615 55444 13671 55500
rect 13739 55444 13795 55500
rect 13863 55444 13919 55500
rect 13987 55444 14043 55500
rect 14111 55444 14167 55500
rect 14235 55444 14291 55500
rect 14359 55444 14415 55500
rect 14483 55444 14539 55500
rect 14607 55444 14663 55500
rect 12871 55320 12927 55376
rect 12995 55320 13051 55376
rect 13119 55320 13175 55376
rect 13243 55320 13299 55376
rect 13367 55320 13423 55376
rect 13491 55320 13547 55376
rect 13615 55320 13671 55376
rect 13739 55320 13795 55376
rect 13863 55320 13919 55376
rect 13987 55320 14043 55376
rect 14111 55320 14167 55376
rect 14235 55320 14291 55376
rect 14359 55320 14415 55376
rect 14483 55320 14539 55376
rect 14607 55320 14663 55376
rect 12871 55196 12927 55252
rect 12995 55196 13051 55252
rect 13119 55196 13175 55252
rect 13243 55196 13299 55252
rect 13367 55196 13423 55252
rect 13491 55196 13547 55252
rect 13615 55196 13671 55252
rect 13739 55196 13795 55252
rect 13863 55196 13919 55252
rect 13987 55196 14043 55252
rect 14111 55196 14167 55252
rect 14235 55196 14291 55252
rect 14359 55196 14415 55252
rect 14483 55196 14539 55252
rect 14607 55196 14663 55252
rect 12871 55072 12927 55128
rect 12995 55072 13051 55128
rect 13119 55072 13175 55128
rect 13243 55072 13299 55128
rect 13367 55072 13423 55128
rect 13491 55072 13547 55128
rect 13615 55072 13671 55128
rect 13739 55072 13795 55128
rect 13863 55072 13919 55128
rect 13987 55072 14043 55128
rect 14111 55072 14167 55128
rect 14235 55072 14291 55128
rect 14359 55072 14415 55128
rect 14483 55072 14539 55128
rect 14607 55072 14663 55128
rect 12871 54948 12927 55004
rect 12995 54948 13051 55004
rect 13119 54948 13175 55004
rect 13243 54948 13299 55004
rect 13367 54948 13423 55004
rect 13491 54948 13547 55004
rect 13615 54948 13671 55004
rect 13739 54948 13795 55004
rect 13863 54948 13919 55004
rect 13987 54948 14043 55004
rect 14111 54948 14167 55004
rect 14235 54948 14291 55004
rect 14359 54948 14415 55004
rect 14483 54948 14539 55004
rect 14607 54948 14663 55004
rect 12871 54824 12927 54880
rect 12995 54824 13051 54880
rect 13119 54824 13175 54880
rect 13243 54824 13299 54880
rect 13367 54824 13423 54880
rect 13491 54824 13547 54880
rect 13615 54824 13671 54880
rect 13739 54824 13795 54880
rect 13863 54824 13919 54880
rect 13987 54824 14043 54880
rect 14111 54824 14167 54880
rect 14235 54824 14291 54880
rect 14359 54824 14415 54880
rect 14483 54824 14539 54880
rect 14607 54824 14663 54880
rect 12871 54700 12927 54756
rect 12995 54700 13051 54756
rect 13119 54700 13175 54756
rect 13243 54700 13299 54756
rect 13367 54700 13423 54756
rect 13491 54700 13547 54756
rect 13615 54700 13671 54756
rect 13739 54700 13795 54756
rect 13863 54700 13919 54756
rect 13987 54700 14043 54756
rect 14111 54700 14167 54756
rect 14235 54700 14291 54756
rect 14359 54700 14415 54756
rect 14483 54700 14539 54756
rect 14607 54700 14663 54756
rect 12871 54576 12927 54632
rect 12995 54576 13051 54632
rect 13119 54576 13175 54632
rect 13243 54576 13299 54632
rect 13367 54576 13423 54632
rect 13491 54576 13547 54632
rect 13615 54576 13671 54632
rect 13739 54576 13795 54632
rect 13863 54576 13919 54632
rect 13987 54576 14043 54632
rect 14111 54576 14167 54632
rect 14235 54576 14291 54632
rect 14359 54576 14415 54632
rect 14483 54576 14539 54632
rect 14607 54576 14663 54632
rect 12871 54452 12927 54508
rect 12995 54452 13051 54508
rect 13119 54452 13175 54508
rect 13243 54452 13299 54508
rect 13367 54452 13423 54508
rect 13491 54452 13547 54508
rect 13615 54452 13671 54508
rect 13739 54452 13795 54508
rect 13863 54452 13919 54508
rect 13987 54452 14043 54508
rect 14111 54452 14167 54508
rect 14235 54452 14291 54508
rect 14359 54452 14415 54508
rect 14483 54452 14539 54508
rect 14607 54452 14663 54508
rect 14902 52574 14958 52576
rect 14902 52522 14904 52574
rect 14904 52522 14956 52574
rect 14956 52522 14958 52574
rect 14902 52466 14958 52522
rect 14902 52414 14904 52466
rect 14904 52414 14956 52466
rect 14956 52414 14958 52466
rect 14902 52358 14958 52414
rect 14902 52306 14904 52358
rect 14904 52306 14956 52358
rect 14956 52306 14958 52358
rect 14902 52250 14958 52306
rect 14902 52198 14904 52250
rect 14904 52198 14956 52250
rect 14956 52198 14958 52250
rect 14902 52142 14958 52198
rect 14902 52090 14904 52142
rect 14904 52090 14956 52142
rect 14956 52090 14958 52142
rect 14902 52034 14958 52090
rect 14902 51982 14904 52034
rect 14904 51982 14956 52034
rect 14956 51982 14958 52034
rect 14902 51926 14958 51982
rect 14902 51874 14904 51926
rect 14904 51874 14956 51926
rect 14956 51874 14958 51926
rect 14902 51818 14958 51874
rect 14902 51766 14904 51818
rect 14904 51766 14956 51818
rect 14956 51766 14958 51818
rect 14902 51710 14958 51766
rect 14902 51658 14904 51710
rect 14904 51658 14956 51710
rect 14956 51658 14958 51710
rect 14902 51602 14958 51658
rect 14902 51550 14904 51602
rect 14904 51550 14956 51602
rect 14956 51550 14958 51602
rect 14902 51494 14958 51550
rect 14902 51442 14904 51494
rect 14904 51442 14956 51494
rect 14956 51442 14958 51494
rect 14902 51386 14958 51442
rect 14902 51334 14904 51386
rect 14904 51334 14956 51386
rect 14956 51334 14958 51386
rect 14902 51278 14958 51334
rect 14902 51226 14904 51278
rect 14904 51226 14956 51278
rect 14956 51226 14958 51278
rect 14902 51224 14958 51226
rect 12871 50892 12927 50948
rect 12995 50892 13051 50948
rect 13119 50892 13175 50948
rect 13243 50892 13299 50948
rect 13367 50892 13423 50948
rect 13491 50892 13547 50948
rect 13615 50892 13671 50948
rect 13739 50892 13795 50948
rect 13863 50892 13919 50948
rect 13987 50892 14043 50948
rect 14111 50892 14167 50948
rect 14235 50892 14291 50948
rect 14359 50892 14415 50948
rect 14483 50892 14539 50948
rect 14607 50892 14663 50948
rect 12871 50768 12927 50824
rect 12995 50768 13051 50824
rect 13119 50768 13175 50824
rect 13243 50768 13299 50824
rect 13367 50768 13423 50824
rect 13491 50768 13547 50824
rect 13615 50768 13671 50824
rect 13739 50768 13795 50824
rect 13863 50768 13919 50824
rect 13987 50768 14043 50824
rect 14111 50768 14167 50824
rect 14235 50768 14291 50824
rect 14359 50768 14415 50824
rect 14483 50768 14539 50824
rect 14607 50768 14663 50824
rect 12871 50644 12927 50700
rect 12995 50644 13051 50700
rect 13119 50644 13175 50700
rect 13243 50644 13299 50700
rect 13367 50644 13423 50700
rect 13491 50644 13547 50700
rect 13615 50644 13671 50700
rect 13739 50644 13795 50700
rect 13863 50644 13919 50700
rect 13987 50644 14043 50700
rect 14111 50644 14167 50700
rect 14235 50644 14291 50700
rect 14359 50644 14415 50700
rect 14483 50644 14539 50700
rect 14607 50644 14663 50700
rect 12871 50520 12927 50576
rect 12995 50520 13051 50576
rect 13119 50520 13175 50576
rect 13243 50520 13299 50576
rect 13367 50520 13423 50576
rect 13491 50520 13547 50576
rect 13615 50520 13671 50576
rect 13739 50520 13795 50576
rect 13863 50520 13919 50576
rect 13987 50520 14043 50576
rect 14111 50520 14167 50576
rect 14235 50520 14291 50576
rect 14359 50520 14415 50576
rect 14483 50520 14539 50576
rect 14607 50520 14663 50576
rect 12871 50396 12927 50452
rect 12995 50396 13051 50452
rect 13119 50396 13175 50452
rect 13243 50396 13299 50452
rect 13367 50396 13423 50452
rect 13491 50396 13547 50452
rect 13615 50396 13671 50452
rect 13739 50396 13795 50452
rect 13863 50396 13919 50452
rect 13987 50396 14043 50452
rect 14111 50396 14167 50452
rect 14235 50396 14291 50452
rect 14359 50396 14415 50452
rect 14483 50396 14539 50452
rect 14607 50396 14663 50452
rect 12871 50272 12927 50328
rect 12995 50272 13051 50328
rect 13119 50272 13175 50328
rect 13243 50272 13299 50328
rect 13367 50272 13423 50328
rect 13491 50272 13547 50328
rect 13615 50272 13671 50328
rect 13739 50272 13795 50328
rect 13863 50272 13919 50328
rect 13987 50272 14043 50328
rect 14111 50272 14167 50328
rect 14235 50272 14291 50328
rect 14359 50272 14415 50328
rect 14483 50272 14539 50328
rect 14607 50272 14663 50328
rect 12871 50148 12927 50204
rect 12995 50148 13051 50204
rect 13119 50148 13175 50204
rect 13243 50148 13299 50204
rect 13367 50148 13423 50204
rect 13491 50148 13547 50204
rect 13615 50148 13671 50204
rect 13739 50148 13795 50204
rect 13863 50148 13919 50204
rect 13987 50148 14043 50204
rect 14111 50148 14167 50204
rect 14235 50148 14291 50204
rect 14359 50148 14415 50204
rect 14483 50148 14539 50204
rect 14607 50148 14663 50204
rect 12871 50024 12927 50080
rect 12995 50024 13051 50080
rect 13119 50024 13175 50080
rect 13243 50024 13299 50080
rect 13367 50024 13423 50080
rect 13491 50024 13547 50080
rect 13615 50024 13671 50080
rect 13739 50024 13795 50080
rect 13863 50024 13919 50080
rect 13987 50024 14043 50080
rect 14111 50024 14167 50080
rect 14235 50024 14291 50080
rect 14359 50024 14415 50080
rect 14483 50024 14539 50080
rect 14607 50024 14663 50080
rect 12871 49900 12927 49956
rect 12995 49900 13051 49956
rect 13119 49900 13175 49956
rect 13243 49900 13299 49956
rect 13367 49900 13423 49956
rect 13491 49900 13547 49956
rect 13615 49900 13671 49956
rect 13739 49900 13795 49956
rect 13863 49900 13919 49956
rect 13987 49900 14043 49956
rect 14111 49900 14167 49956
rect 14235 49900 14291 49956
rect 14359 49900 14415 49956
rect 14483 49900 14539 49956
rect 14607 49900 14663 49956
rect 12871 49776 12927 49832
rect 12995 49776 13051 49832
rect 13119 49776 13175 49832
rect 13243 49776 13299 49832
rect 13367 49776 13423 49832
rect 13491 49776 13547 49832
rect 13615 49776 13671 49832
rect 13739 49776 13795 49832
rect 13863 49776 13919 49832
rect 13987 49776 14043 49832
rect 14111 49776 14167 49832
rect 14235 49776 14291 49832
rect 14359 49776 14415 49832
rect 14483 49776 14539 49832
rect 14607 49776 14663 49832
rect 12871 49652 12927 49708
rect 12995 49652 13051 49708
rect 13119 49652 13175 49708
rect 13243 49652 13299 49708
rect 13367 49652 13423 49708
rect 13491 49652 13547 49708
rect 13615 49652 13671 49708
rect 13739 49652 13795 49708
rect 13863 49652 13919 49708
rect 13987 49652 14043 49708
rect 14111 49652 14167 49708
rect 14235 49652 14291 49708
rect 14359 49652 14415 49708
rect 14483 49652 14539 49708
rect 14607 49652 14663 49708
rect 12871 47692 12927 47748
rect 12995 47692 13051 47748
rect 13119 47692 13175 47748
rect 13243 47692 13299 47748
rect 13367 47692 13423 47748
rect 13491 47692 13547 47748
rect 13615 47692 13671 47748
rect 13739 47692 13795 47748
rect 13863 47692 13919 47748
rect 13987 47692 14043 47748
rect 14111 47692 14167 47748
rect 14235 47692 14291 47748
rect 14359 47692 14415 47748
rect 14483 47692 14539 47748
rect 14607 47692 14663 47748
rect 12871 47568 12927 47624
rect 12995 47568 13051 47624
rect 13119 47568 13175 47624
rect 13243 47568 13299 47624
rect 13367 47568 13423 47624
rect 13491 47568 13547 47624
rect 13615 47568 13671 47624
rect 13739 47568 13795 47624
rect 13863 47568 13919 47624
rect 13987 47568 14043 47624
rect 14111 47568 14167 47624
rect 14235 47568 14291 47624
rect 14359 47568 14415 47624
rect 14483 47568 14539 47624
rect 14607 47568 14663 47624
rect 12871 47444 12927 47500
rect 12995 47444 13051 47500
rect 13119 47444 13175 47500
rect 13243 47444 13299 47500
rect 13367 47444 13423 47500
rect 13491 47444 13547 47500
rect 13615 47444 13671 47500
rect 13739 47444 13795 47500
rect 13863 47444 13919 47500
rect 13987 47444 14043 47500
rect 14111 47444 14167 47500
rect 14235 47444 14291 47500
rect 14359 47444 14415 47500
rect 14483 47444 14539 47500
rect 14607 47444 14663 47500
rect 12871 47320 12927 47376
rect 12995 47320 13051 47376
rect 13119 47320 13175 47376
rect 13243 47320 13299 47376
rect 13367 47320 13423 47376
rect 13491 47320 13547 47376
rect 13615 47320 13671 47376
rect 13739 47320 13795 47376
rect 13863 47320 13919 47376
rect 13987 47320 14043 47376
rect 14111 47320 14167 47376
rect 14235 47320 14291 47376
rect 14359 47320 14415 47376
rect 14483 47320 14539 47376
rect 14607 47320 14663 47376
rect 2808 47196 2864 47252
rect 2932 47196 2988 47252
rect 3056 47196 3112 47252
rect 3180 47196 3236 47252
rect 3304 47196 3360 47252
rect 3428 47196 3484 47252
rect 3552 47196 3608 47252
rect 3676 47196 3732 47252
rect 3800 47196 3856 47252
rect 3924 47196 3980 47252
rect 4048 47196 4104 47252
rect 4172 47196 4228 47252
rect 4296 47196 4352 47252
rect 4420 47196 4476 47252
rect 4544 47196 4600 47252
rect 4668 47196 4724 47252
rect 2808 47072 2864 47128
rect 2932 47072 2988 47128
rect 3056 47072 3112 47128
rect 3180 47072 3236 47128
rect 3304 47072 3360 47128
rect 3428 47072 3484 47128
rect 3552 47072 3608 47128
rect 3676 47072 3732 47128
rect 3800 47072 3856 47128
rect 3924 47072 3980 47128
rect 4048 47072 4104 47128
rect 4172 47072 4228 47128
rect 4296 47072 4352 47128
rect 4420 47072 4476 47128
rect 4544 47072 4600 47128
rect 4668 47072 4724 47128
rect 2808 46948 2864 47004
rect 2932 46948 2988 47004
rect 3056 46948 3112 47004
rect 3180 46948 3236 47004
rect 3304 46948 3360 47004
rect 3428 46948 3484 47004
rect 3552 46948 3608 47004
rect 3676 46948 3732 47004
rect 3800 46948 3856 47004
rect 3924 46948 3980 47004
rect 4048 46948 4104 47004
rect 4172 46948 4228 47004
rect 4296 46948 4352 47004
rect 4420 46948 4476 47004
rect 4544 46948 4600 47004
rect 4668 46948 4724 47004
rect 2808 46824 2864 46880
rect 2932 46824 2988 46880
rect 3056 46824 3112 46880
rect 3180 46824 3236 46880
rect 3304 46824 3360 46880
rect 3428 46824 3484 46880
rect 3552 46824 3608 46880
rect 3676 46824 3732 46880
rect 3800 46824 3856 46880
rect 3924 46824 3980 46880
rect 4048 46824 4104 46880
rect 4172 46824 4228 46880
rect 4296 46824 4352 46880
rect 4420 46824 4476 46880
rect 4544 46824 4600 46880
rect 4668 46824 4724 46880
rect 2808 46700 2864 46756
rect 2932 46700 2988 46756
rect 3056 46700 3112 46756
rect 3180 46700 3236 46756
rect 3304 46700 3360 46756
rect 3428 46700 3484 46756
rect 3552 46700 3608 46756
rect 3676 46700 3732 46756
rect 3800 46700 3856 46756
rect 3924 46700 3980 46756
rect 4048 46700 4104 46756
rect 4172 46700 4228 46756
rect 4296 46700 4352 46756
rect 4420 46700 4476 46756
rect 4544 46700 4600 46756
rect 4668 46700 4724 46756
rect 2808 46576 2864 46632
rect 2932 46576 2988 46632
rect 3056 46576 3112 46632
rect 3180 46576 3236 46632
rect 3304 46576 3360 46632
rect 3428 46576 3484 46632
rect 3552 46576 3608 46632
rect 3676 46576 3732 46632
rect 3800 46576 3856 46632
rect 3924 46576 3980 46632
rect 4048 46576 4104 46632
rect 4172 46576 4228 46632
rect 4296 46576 4352 46632
rect 4420 46576 4476 46632
rect 4544 46576 4600 46632
rect 4668 46576 4724 46632
rect 2808 46452 2864 46508
rect 2932 46452 2988 46508
rect 3056 46452 3112 46508
rect 3180 46452 3236 46508
rect 3304 46452 3360 46508
rect 3428 46452 3484 46508
rect 3552 46452 3608 46508
rect 3676 46452 3732 46508
rect 3800 46452 3856 46508
rect 3924 46452 3980 46508
rect 4048 46452 4104 46508
rect 4172 46452 4228 46508
rect 4296 46452 4352 46508
rect 4420 46452 4476 46508
rect 4544 46452 4600 46508
rect 4668 46452 4724 46508
rect 5178 47196 5234 47252
rect 5302 47196 5358 47252
rect 5426 47196 5482 47252
rect 5550 47196 5606 47252
rect 5674 47196 5730 47252
rect 5798 47196 5854 47252
rect 5922 47196 5978 47252
rect 6046 47196 6102 47252
rect 6170 47196 6226 47252
rect 6294 47196 6350 47252
rect 6418 47196 6474 47252
rect 6542 47196 6598 47252
rect 6666 47196 6722 47252
rect 6790 47196 6846 47252
rect 6914 47196 6970 47252
rect 7038 47196 7094 47252
rect 5178 47072 5234 47128
rect 5302 47072 5358 47128
rect 5426 47072 5482 47128
rect 5550 47072 5606 47128
rect 5674 47072 5730 47128
rect 5798 47072 5854 47128
rect 5922 47072 5978 47128
rect 6046 47072 6102 47128
rect 6170 47072 6226 47128
rect 6294 47072 6350 47128
rect 6418 47072 6474 47128
rect 6542 47072 6598 47128
rect 6666 47072 6722 47128
rect 6790 47072 6846 47128
rect 6914 47072 6970 47128
rect 7038 47072 7094 47128
rect 5178 46948 5234 47004
rect 5302 46948 5358 47004
rect 5426 46948 5482 47004
rect 5550 46948 5606 47004
rect 5674 46948 5730 47004
rect 5798 46948 5854 47004
rect 5922 46948 5978 47004
rect 6046 46948 6102 47004
rect 6170 46948 6226 47004
rect 6294 46948 6350 47004
rect 6418 46948 6474 47004
rect 6542 46948 6598 47004
rect 6666 46948 6722 47004
rect 6790 46948 6846 47004
rect 6914 46948 6970 47004
rect 7038 46948 7094 47004
rect 5178 46824 5234 46880
rect 5302 46824 5358 46880
rect 5426 46824 5482 46880
rect 5550 46824 5606 46880
rect 5674 46824 5730 46880
rect 5798 46824 5854 46880
rect 5922 46824 5978 46880
rect 6046 46824 6102 46880
rect 6170 46824 6226 46880
rect 6294 46824 6350 46880
rect 6418 46824 6474 46880
rect 6542 46824 6598 46880
rect 6666 46824 6722 46880
rect 6790 46824 6846 46880
rect 6914 46824 6970 46880
rect 7038 46824 7094 46880
rect 5178 46700 5234 46756
rect 5302 46700 5358 46756
rect 5426 46700 5482 46756
rect 5550 46700 5606 46756
rect 5674 46700 5730 46756
rect 5798 46700 5854 46756
rect 5922 46700 5978 46756
rect 6046 46700 6102 46756
rect 6170 46700 6226 46756
rect 6294 46700 6350 46756
rect 6418 46700 6474 46756
rect 6542 46700 6598 46756
rect 6666 46700 6722 46756
rect 6790 46700 6846 46756
rect 6914 46700 6970 46756
rect 7038 46700 7094 46756
rect 5178 46576 5234 46632
rect 5302 46576 5358 46632
rect 5426 46576 5482 46632
rect 5550 46576 5606 46632
rect 5674 46576 5730 46632
rect 5798 46576 5854 46632
rect 5922 46576 5978 46632
rect 6046 46576 6102 46632
rect 6170 46576 6226 46632
rect 6294 46576 6350 46632
rect 6418 46576 6474 46632
rect 6542 46576 6598 46632
rect 6666 46576 6722 46632
rect 6790 46576 6846 46632
rect 6914 46576 6970 46632
rect 7038 46576 7094 46632
rect 5178 46452 5234 46508
rect 5302 46452 5358 46508
rect 5426 46452 5482 46508
rect 5550 46452 5606 46508
rect 5674 46452 5730 46508
rect 5798 46452 5854 46508
rect 5922 46452 5978 46508
rect 6046 46452 6102 46508
rect 6170 46452 6226 46508
rect 6294 46452 6350 46508
rect 6418 46452 6474 46508
rect 6542 46452 6598 46508
rect 6666 46452 6722 46508
rect 6790 46452 6846 46508
rect 6914 46452 6970 46508
rect 7038 46452 7094 46508
rect 7884 47196 7940 47252
rect 8008 47196 8064 47252
rect 8132 47196 8188 47252
rect 8256 47196 8312 47252
rect 8380 47196 8436 47252
rect 8504 47196 8560 47252
rect 8628 47196 8684 47252
rect 8752 47196 8808 47252
rect 8876 47196 8932 47252
rect 9000 47196 9056 47252
rect 9124 47196 9180 47252
rect 9248 47196 9304 47252
rect 9372 47196 9428 47252
rect 9496 47196 9552 47252
rect 9620 47196 9676 47252
rect 9744 47196 9800 47252
rect 7884 47072 7940 47128
rect 8008 47072 8064 47128
rect 8132 47072 8188 47128
rect 8256 47072 8312 47128
rect 8380 47072 8436 47128
rect 8504 47072 8560 47128
rect 8628 47072 8684 47128
rect 8752 47072 8808 47128
rect 8876 47072 8932 47128
rect 9000 47072 9056 47128
rect 9124 47072 9180 47128
rect 9248 47072 9304 47128
rect 9372 47072 9428 47128
rect 9496 47072 9552 47128
rect 9620 47072 9676 47128
rect 9744 47072 9800 47128
rect 7884 46948 7940 47004
rect 8008 46948 8064 47004
rect 8132 46948 8188 47004
rect 8256 46948 8312 47004
rect 8380 46948 8436 47004
rect 8504 46948 8560 47004
rect 8628 46948 8684 47004
rect 8752 46948 8808 47004
rect 8876 46948 8932 47004
rect 9000 46948 9056 47004
rect 9124 46948 9180 47004
rect 9248 46948 9304 47004
rect 9372 46948 9428 47004
rect 9496 46948 9552 47004
rect 9620 46948 9676 47004
rect 9744 46948 9800 47004
rect 7884 46824 7940 46880
rect 8008 46824 8064 46880
rect 8132 46824 8188 46880
rect 8256 46824 8312 46880
rect 8380 46824 8436 46880
rect 8504 46824 8560 46880
rect 8628 46824 8684 46880
rect 8752 46824 8808 46880
rect 8876 46824 8932 46880
rect 9000 46824 9056 46880
rect 9124 46824 9180 46880
rect 9248 46824 9304 46880
rect 9372 46824 9428 46880
rect 9496 46824 9552 46880
rect 9620 46824 9676 46880
rect 9744 46824 9800 46880
rect 7884 46700 7940 46756
rect 8008 46700 8064 46756
rect 8132 46700 8188 46756
rect 8256 46700 8312 46756
rect 8380 46700 8436 46756
rect 8504 46700 8560 46756
rect 8628 46700 8684 46756
rect 8752 46700 8808 46756
rect 8876 46700 8932 46756
rect 9000 46700 9056 46756
rect 9124 46700 9180 46756
rect 9248 46700 9304 46756
rect 9372 46700 9428 46756
rect 9496 46700 9552 46756
rect 9620 46700 9676 46756
rect 9744 46700 9800 46756
rect 7884 46576 7940 46632
rect 8008 46576 8064 46632
rect 8132 46576 8188 46632
rect 8256 46576 8312 46632
rect 8380 46576 8436 46632
rect 8504 46576 8560 46632
rect 8628 46576 8684 46632
rect 8752 46576 8808 46632
rect 8876 46576 8932 46632
rect 9000 46576 9056 46632
rect 9124 46576 9180 46632
rect 9248 46576 9304 46632
rect 9372 46576 9428 46632
rect 9496 46576 9552 46632
rect 9620 46576 9676 46632
rect 9744 46576 9800 46632
rect 7884 46452 7940 46508
rect 8008 46452 8064 46508
rect 8132 46452 8188 46508
rect 8256 46452 8312 46508
rect 8380 46452 8436 46508
rect 8504 46452 8560 46508
rect 8628 46452 8684 46508
rect 8752 46452 8808 46508
rect 8876 46452 8932 46508
rect 9000 46452 9056 46508
rect 9124 46452 9180 46508
rect 9248 46452 9304 46508
rect 9372 46452 9428 46508
rect 9496 46452 9552 46508
rect 9620 46452 9676 46508
rect 9744 46452 9800 46508
rect 10254 47196 10310 47252
rect 10378 47196 10434 47252
rect 10502 47196 10558 47252
rect 10626 47196 10682 47252
rect 10750 47196 10806 47252
rect 10874 47196 10930 47252
rect 10998 47196 11054 47252
rect 11122 47196 11178 47252
rect 11246 47196 11302 47252
rect 11370 47196 11426 47252
rect 11494 47196 11550 47252
rect 11618 47196 11674 47252
rect 11742 47196 11798 47252
rect 11866 47196 11922 47252
rect 11990 47196 12046 47252
rect 12114 47196 12170 47252
rect 10254 47072 10310 47128
rect 10378 47072 10434 47128
rect 10502 47072 10558 47128
rect 10626 47072 10682 47128
rect 10750 47072 10806 47128
rect 10874 47072 10930 47128
rect 10998 47072 11054 47128
rect 11122 47072 11178 47128
rect 11246 47072 11302 47128
rect 11370 47072 11426 47128
rect 11494 47072 11550 47128
rect 11618 47072 11674 47128
rect 11742 47072 11798 47128
rect 11866 47072 11922 47128
rect 11990 47072 12046 47128
rect 12114 47072 12170 47128
rect 10254 46948 10310 47004
rect 10378 46948 10434 47004
rect 10502 46948 10558 47004
rect 10626 46948 10682 47004
rect 10750 46948 10806 47004
rect 10874 46948 10930 47004
rect 10998 46948 11054 47004
rect 11122 46948 11178 47004
rect 11246 46948 11302 47004
rect 11370 46948 11426 47004
rect 11494 46948 11550 47004
rect 11618 46948 11674 47004
rect 11742 46948 11798 47004
rect 11866 46948 11922 47004
rect 11990 46948 12046 47004
rect 12114 46948 12170 47004
rect 10254 46824 10310 46880
rect 10378 46824 10434 46880
rect 10502 46824 10558 46880
rect 10626 46824 10682 46880
rect 10750 46824 10806 46880
rect 10874 46824 10930 46880
rect 10998 46824 11054 46880
rect 11122 46824 11178 46880
rect 11246 46824 11302 46880
rect 11370 46824 11426 46880
rect 11494 46824 11550 46880
rect 11618 46824 11674 46880
rect 11742 46824 11798 46880
rect 11866 46824 11922 46880
rect 11990 46824 12046 46880
rect 12114 46824 12170 46880
rect 10254 46700 10310 46756
rect 10378 46700 10434 46756
rect 10502 46700 10558 46756
rect 10626 46700 10682 46756
rect 10750 46700 10806 46756
rect 10874 46700 10930 46756
rect 10998 46700 11054 46756
rect 11122 46700 11178 46756
rect 11246 46700 11302 46756
rect 11370 46700 11426 46756
rect 11494 46700 11550 46756
rect 11618 46700 11674 46756
rect 11742 46700 11798 46756
rect 11866 46700 11922 46756
rect 11990 46700 12046 46756
rect 12114 46700 12170 46756
rect 10254 46576 10310 46632
rect 10378 46576 10434 46632
rect 10502 46576 10558 46632
rect 10626 46576 10682 46632
rect 10750 46576 10806 46632
rect 10874 46576 10930 46632
rect 10998 46576 11054 46632
rect 11122 46576 11178 46632
rect 11246 46576 11302 46632
rect 11370 46576 11426 46632
rect 11494 46576 11550 46632
rect 11618 46576 11674 46632
rect 11742 46576 11798 46632
rect 11866 46576 11922 46632
rect 11990 46576 12046 46632
rect 12114 46576 12170 46632
rect 10254 46452 10310 46508
rect 10378 46452 10434 46508
rect 10502 46452 10558 46508
rect 10626 46452 10682 46508
rect 10750 46452 10806 46508
rect 10874 46452 10930 46508
rect 10998 46452 11054 46508
rect 11122 46452 11178 46508
rect 11246 46452 11302 46508
rect 11370 46452 11426 46508
rect 11494 46452 11550 46508
rect 11618 46452 11674 46508
rect 11742 46452 11798 46508
rect 11866 46452 11922 46508
rect 11990 46452 12046 46508
rect 12114 46452 12170 46508
rect 12871 47196 12927 47252
rect 12995 47196 13051 47252
rect 13119 47196 13175 47252
rect 13243 47196 13299 47252
rect 13367 47196 13423 47252
rect 13491 47196 13547 47252
rect 13615 47196 13671 47252
rect 13739 47196 13795 47252
rect 13863 47196 13919 47252
rect 13987 47196 14043 47252
rect 14111 47196 14167 47252
rect 14235 47196 14291 47252
rect 14359 47196 14415 47252
rect 14483 47196 14539 47252
rect 14607 47196 14663 47252
rect 12871 47072 12927 47128
rect 12995 47072 13051 47128
rect 13119 47072 13175 47128
rect 13243 47072 13299 47128
rect 13367 47072 13423 47128
rect 13491 47072 13547 47128
rect 13615 47072 13671 47128
rect 13739 47072 13795 47128
rect 13863 47072 13919 47128
rect 13987 47072 14043 47128
rect 14111 47072 14167 47128
rect 14235 47072 14291 47128
rect 14359 47072 14415 47128
rect 14483 47072 14539 47128
rect 14607 47072 14663 47128
rect 12871 46948 12927 47004
rect 12995 46948 13051 47004
rect 13119 46948 13175 47004
rect 13243 46948 13299 47004
rect 13367 46948 13423 47004
rect 13491 46948 13547 47004
rect 13615 46948 13671 47004
rect 13739 46948 13795 47004
rect 13863 46948 13919 47004
rect 13987 46948 14043 47004
rect 14111 46948 14167 47004
rect 14235 46948 14291 47004
rect 14359 46948 14415 47004
rect 14483 46948 14539 47004
rect 14607 46948 14663 47004
rect 12871 46824 12927 46880
rect 12995 46824 13051 46880
rect 13119 46824 13175 46880
rect 13243 46824 13299 46880
rect 13367 46824 13423 46880
rect 13491 46824 13547 46880
rect 13615 46824 13671 46880
rect 13739 46824 13795 46880
rect 13863 46824 13919 46880
rect 13987 46824 14043 46880
rect 14111 46824 14167 46880
rect 14235 46824 14291 46880
rect 14359 46824 14415 46880
rect 14483 46824 14539 46880
rect 14607 46824 14663 46880
rect 12871 46700 12927 46756
rect 12995 46700 13051 46756
rect 13119 46700 13175 46756
rect 13243 46700 13299 46756
rect 13367 46700 13423 46756
rect 13491 46700 13547 46756
rect 13615 46700 13671 46756
rect 13739 46700 13795 46756
rect 13863 46700 13919 46756
rect 13987 46700 14043 46756
rect 14111 46700 14167 46756
rect 14235 46700 14291 46756
rect 14359 46700 14415 46756
rect 14483 46700 14539 46756
rect 14607 46700 14663 46756
rect 12871 46576 12927 46632
rect 12995 46576 13051 46632
rect 13119 46576 13175 46632
rect 13243 46576 13299 46632
rect 13367 46576 13423 46632
rect 13491 46576 13547 46632
rect 13615 46576 13671 46632
rect 13739 46576 13795 46632
rect 13863 46576 13919 46632
rect 13987 46576 14043 46632
rect 14111 46576 14167 46632
rect 14235 46576 14291 46632
rect 14359 46576 14415 46632
rect 14483 46576 14539 46632
rect 14607 46576 14663 46632
rect 12871 46452 12927 46508
rect 12995 46452 13051 46508
rect 13119 46452 13175 46508
rect 13243 46452 13299 46508
rect 13367 46452 13423 46508
rect 13491 46452 13547 46508
rect 13615 46452 13671 46508
rect 13739 46452 13795 46508
rect 13863 46452 13919 46508
rect 13987 46452 14043 46508
rect 14111 46452 14167 46508
rect 14235 46452 14291 46508
rect 14359 46452 14415 46508
rect 14483 46452 14539 46508
rect 14607 46452 14663 46508
rect 2491 46092 2547 46148
rect 2615 46092 2671 46148
rect 2491 45968 2547 46024
rect 2615 45968 2671 46024
rect 2491 45844 2547 45900
rect 2615 45844 2671 45900
rect 2491 45720 2547 45776
rect 2615 45720 2671 45776
rect 2491 45596 2547 45652
rect 2615 45596 2671 45652
rect 2491 45472 2547 45528
rect 2615 45472 2671 45528
rect 2491 45348 2547 45404
rect 2615 45348 2671 45404
rect 2491 45224 2547 45280
rect 2615 45224 2671 45280
rect 2491 45100 2547 45156
rect 2615 45100 2671 45156
rect 2491 44976 2547 45032
rect 2615 44976 2671 45032
rect 2491 44852 2547 44908
rect 2615 44852 2671 44908
rect 4861 46092 4917 46148
rect 4985 46092 5041 46148
rect 4861 45968 4917 46024
rect 4985 45968 5041 46024
rect 4861 45844 4917 45900
rect 4985 45844 5041 45900
rect 4861 45720 4917 45776
rect 4985 45720 5041 45776
rect 4861 45596 4917 45652
rect 4985 45596 5041 45652
rect 4861 45472 4917 45528
rect 4985 45472 5041 45528
rect 4861 45348 4917 45404
rect 4985 45348 5041 45404
rect 4861 45224 4917 45280
rect 4985 45224 5041 45280
rect 4861 45100 4917 45156
rect 4985 45100 5041 45156
rect 4861 44976 4917 45032
rect 4985 44976 5041 45032
rect 4861 44852 4917 44908
rect 4985 44852 5041 44908
rect 7275 46092 7331 46148
rect 7399 46092 7455 46148
rect 7523 46092 7579 46148
rect 7647 46092 7703 46148
rect 7275 45968 7331 46024
rect 7399 45968 7455 46024
rect 7523 45968 7579 46024
rect 7647 45968 7703 46024
rect 7275 45844 7331 45900
rect 7399 45844 7455 45900
rect 7523 45844 7579 45900
rect 7647 45844 7703 45900
rect 7275 45720 7331 45776
rect 7399 45720 7455 45776
rect 7523 45720 7579 45776
rect 7647 45720 7703 45776
rect 7275 45596 7331 45652
rect 7399 45596 7455 45652
rect 7523 45596 7579 45652
rect 7647 45596 7703 45652
rect 7275 45472 7331 45528
rect 7399 45472 7455 45528
rect 7523 45472 7579 45528
rect 7647 45472 7703 45528
rect 7275 45348 7331 45404
rect 7399 45348 7455 45404
rect 7523 45348 7579 45404
rect 7647 45348 7703 45404
rect 7275 45224 7331 45280
rect 7399 45224 7455 45280
rect 7523 45224 7579 45280
rect 7647 45224 7703 45280
rect 7275 45100 7331 45156
rect 7399 45100 7455 45156
rect 7523 45100 7579 45156
rect 7647 45100 7703 45156
rect 7275 44976 7331 45032
rect 7399 44976 7455 45032
rect 7523 44976 7579 45032
rect 7647 44976 7703 45032
rect 7275 44852 7331 44908
rect 7399 44852 7455 44908
rect 7523 44852 7579 44908
rect 7647 44852 7703 44908
rect 9937 46092 9993 46148
rect 10061 46092 10117 46148
rect 9937 45968 9993 46024
rect 10061 45968 10117 46024
rect 9937 45844 9993 45900
rect 10061 45844 10117 45900
rect 9937 45720 9993 45776
rect 10061 45720 10117 45776
rect 9937 45596 9993 45652
rect 10061 45596 10117 45652
rect 9937 45472 9993 45528
rect 10061 45472 10117 45528
rect 9937 45348 9993 45404
rect 10061 45348 10117 45404
rect 9937 45224 9993 45280
rect 10061 45224 10117 45280
rect 9937 45100 9993 45156
rect 10061 45100 10117 45156
rect 9937 44976 9993 45032
rect 10061 44976 10117 45032
rect 9937 44852 9993 44908
rect 10061 44852 10117 44908
rect 12307 46092 12363 46148
rect 12431 46092 12487 46148
rect 12307 45968 12363 46024
rect 12431 45968 12487 46024
rect 12307 45844 12363 45900
rect 12431 45844 12487 45900
rect 12307 45720 12363 45776
rect 12431 45720 12487 45776
rect 12307 45596 12363 45652
rect 12431 45596 12487 45652
rect 12307 45472 12363 45528
rect 12431 45472 12487 45528
rect 12307 45348 12363 45404
rect 12431 45348 12487 45404
rect 12307 45224 12363 45280
rect 12431 45224 12487 45280
rect 12307 45100 12363 45156
rect 12431 45100 12487 45156
rect 12307 44976 12363 45032
rect 12431 44976 12487 45032
rect 12307 44852 12363 44908
rect 12431 44852 12487 44908
rect 2808 44492 2864 44548
rect 2932 44492 2988 44548
rect 3056 44492 3112 44548
rect 3180 44492 3236 44548
rect 3304 44492 3360 44548
rect 3428 44492 3484 44548
rect 3552 44492 3608 44548
rect 3676 44492 3732 44548
rect 3800 44492 3856 44548
rect 3924 44492 3980 44548
rect 4048 44492 4104 44548
rect 4172 44492 4228 44548
rect 4296 44492 4352 44548
rect 4420 44492 4476 44548
rect 4544 44492 4600 44548
rect 4668 44492 4724 44548
rect 2808 44368 2864 44424
rect 2932 44368 2988 44424
rect 3056 44368 3112 44424
rect 3180 44368 3236 44424
rect 3304 44368 3360 44424
rect 3428 44368 3484 44424
rect 3552 44368 3608 44424
rect 3676 44368 3732 44424
rect 3800 44368 3856 44424
rect 3924 44368 3980 44424
rect 4048 44368 4104 44424
rect 4172 44368 4228 44424
rect 4296 44368 4352 44424
rect 4420 44368 4476 44424
rect 4544 44368 4600 44424
rect 4668 44368 4724 44424
rect 2808 44244 2864 44300
rect 2932 44244 2988 44300
rect 3056 44244 3112 44300
rect 3180 44244 3236 44300
rect 3304 44244 3360 44300
rect 3428 44244 3484 44300
rect 3552 44244 3608 44300
rect 3676 44244 3732 44300
rect 3800 44244 3856 44300
rect 3924 44244 3980 44300
rect 4048 44244 4104 44300
rect 4172 44244 4228 44300
rect 4296 44244 4352 44300
rect 4420 44244 4476 44300
rect 4544 44244 4600 44300
rect 4668 44244 4724 44300
rect 2808 44120 2864 44176
rect 2932 44120 2988 44176
rect 3056 44120 3112 44176
rect 3180 44120 3236 44176
rect 3304 44120 3360 44176
rect 3428 44120 3484 44176
rect 3552 44120 3608 44176
rect 3676 44120 3732 44176
rect 3800 44120 3856 44176
rect 3924 44120 3980 44176
rect 4048 44120 4104 44176
rect 4172 44120 4228 44176
rect 4296 44120 4352 44176
rect 4420 44120 4476 44176
rect 4544 44120 4600 44176
rect 4668 44120 4724 44176
rect 2808 43996 2864 44052
rect 2932 43996 2988 44052
rect 3056 43996 3112 44052
rect 3180 43996 3236 44052
rect 3304 43996 3360 44052
rect 3428 43996 3484 44052
rect 3552 43996 3608 44052
rect 3676 43996 3732 44052
rect 3800 43996 3856 44052
rect 3924 43996 3980 44052
rect 4048 43996 4104 44052
rect 4172 43996 4228 44052
rect 4296 43996 4352 44052
rect 4420 43996 4476 44052
rect 4544 43996 4600 44052
rect 4668 43996 4724 44052
rect 2808 43872 2864 43928
rect 2932 43872 2988 43928
rect 3056 43872 3112 43928
rect 3180 43872 3236 43928
rect 3304 43872 3360 43928
rect 3428 43872 3484 43928
rect 3552 43872 3608 43928
rect 3676 43872 3732 43928
rect 3800 43872 3856 43928
rect 3924 43872 3980 43928
rect 4048 43872 4104 43928
rect 4172 43872 4228 43928
rect 4296 43872 4352 43928
rect 4420 43872 4476 43928
rect 4544 43872 4600 43928
rect 4668 43872 4724 43928
rect 2808 43748 2864 43804
rect 2932 43748 2988 43804
rect 3056 43748 3112 43804
rect 3180 43748 3236 43804
rect 3304 43748 3360 43804
rect 3428 43748 3484 43804
rect 3552 43748 3608 43804
rect 3676 43748 3732 43804
rect 3800 43748 3856 43804
rect 3924 43748 3980 43804
rect 4048 43748 4104 43804
rect 4172 43748 4228 43804
rect 4296 43748 4352 43804
rect 4420 43748 4476 43804
rect 4544 43748 4600 43804
rect 4668 43748 4724 43804
rect 2808 43624 2864 43680
rect 2932 43624 2988 43680
rect 3056 43624 3112 43680
rect 3180 43624 3236 43680
rect 3304 43624 3360 43680
rect 3428 43624 3484 43680
rect 3552 43624 3608 43680
rect 3676 43624 3732 43680
rect 3800 43624 3856 43680
rect 3924 43624 3980 43680
rect 4048 43624 4104 43680
rect 4172 43624 4228 43680
rect 4296 43624 4352 43680
rect 4420 43624 4476 43680
rect 4544 43624 4600 43680
rect 4668 43624 4724 43680
rect 2808 43500 2864 43556
rect 2932 43500 2988 43556
rect 3056 43500 3112 43556
rect 3180 43500 3236 43556
rect 3304 43500 3360 43556
rect 3428 43500 3484 43556
rect 3552 43500 3608 43556
rect 3676 43500 3732 43556
rect 3800 43500 3856 43556
rect 3924 43500 3980 43556
rect 4048 43500 4104 43556
rect 4172 43500 4228 43556
rect 4296 43500 4352 43556
rect 4420 43500 4476 43556
rect 4544 43500 4600 43556
rect 4668 43500 4724 43556
rect 2808 43376 2864 43432
rect 2932 43376 2988 43432
rect 3056 43376 3112 43432
rect 3180 43376 3236 43432
rect 3304 43376 3360 43432
rect 3428 43376 3484 43432
rect 3552 43376 3608 43432
rect 3676 43376 3732 43432
rect 3800 43376 3856 43432
rect 3924 43376 3980 43432
rect 4048 43376 4104 43432
rect 4172 43376 4228 43432
rect 4296 43376 4352 43432
rect 4420 43376 4476 43432
rect 4544 43376 4600 43432
rect 4668 43376 4724 43432
rect 2808 43252 2864 43308
rect 2932 43252 2988 43308
rect 3056 43252 3112 43308
rect 3180 43252 3236 43308
rect 3304 43252 3360 43308
rect 3428 43252 3484 43308
rect 3552 43252 3608 43308
rect 3676 43252 3732 43308
rect 3800 43252 3856 43308
rect 3924 43252 3980 43308
rect 4048 43252 4104 43308
rect 4172 43252 4228 43308
rect 4296 43252 4352 43308
rect 4420 43252 4476 43308
rect 4544 43252 4600 43308
rect 4668 43252 4724 43308
rect 5178 44492 5234 44548
rect 5302 44492 5358 44548
rect 5426 44492 5482 44548
rect 5550 44492 5606 44548
rect 5674 44492 5730 44548
rect 5798 44492 5854 44548
rect 5922 44492 5978 44548
rect 6046 44492 6102 44548
rect 6170 44492 6226 44548
rect 6294 44492 6350 44548
rect 6418 44492 6474 44548
rect 6542 44492 6598 44548
rect 6666 44492 6722 44548
rect 6790 44492 6846 44548
rect 6914 44492 6970 44548
rect 7038 44492 7094 44548
rect 5178 44368 5234 44424
rect 5302 44368 5358 44424
rect 5426 44368 5482 44424
rect 5550 44368 5606 44424
rect 5674 44368 5730 44424
rect 5798 44368 5854 44424
rect 5922 44368 5978 44424
rect 6046 44368 6102 44424
rect 6170 44368 6226 44424
rect 6294 44368 6350 44424
rect 6418 44368 6474 44424
rect 6542 44368 6598 44424
rect 6666 44368 6722 44424
rect 6790 44368 6846 44424
rect 6914 44368 6970 44424
rect 7038 44368 7094 44424
rect 5178 44244 5234 44300
rect 5302 44244 5358 44300
rect 5426 44244 5482 44300
rect 5550 44244 5606 44300
rect 5674 44244 5730 44300
rect 5798 44244 5854 44300
rect 5922 44244 5978 44300
rect 6046 44244 6102 44300
rect 6170 44244 6226 44300
rect 6294 44244 6350 44300
rect 6418 44244 6474 44300
rect 6542 44244 6598 44300
rect 6666 44244 6722 44300
rect 6790 44244 6846 44300
rect 6914 44244 6970 44300
rect 7038 44244 7094 44300
rect 5178 44120 5234 44176
rect 5302 44120 5358 44176
rect 5426 44120 5482 44176
rect 5550 44120 5606 44176
rect 5674 44120 5730 44176
rect 5798 44120 5854 44176
rect 5922 44120 5978 44176
rect 6046 44120 6102 44176
rect 6170 44120 6226 44176
rect 6294 44120 6350 44176
rect 6418 44120 6474 44176
rect 6542 44120 6598 44176
rect 6666 44120 6722 44176
rect 6790 44120 6846 44176
rect 6914 44120 6970 44176
rect 7038 44120 7094 44176
rect 5178 43996 5234 44052
rect 5302 43996 5358 44052
rect 5426 43996 5482 44052
rect 5550 43996 5606 44052
rect 5674 43996 5730 44052
rect 5798 43996 5854 44052
rect 5922 43996 5978 44052
rect 6046 43996 6102 44052
rect 6170 43996 6226 44052
rect 6294 43996 6350 44052
rect 6418 43996 6474 44052
rect 6542 43996 6598 44052
rect 6666 43996 6722 44052
rect 6790 43996 6846 44052
rect 6914 43996 6970 44052
rect 7038 43996 7094 44052
rect 5178 43872 5234 43928
rect 5302 43872 5358 43928
rect 5426 43872 5482 43928
rect 5550 43872 5606 43928
rect 5674 43872 5730 43928
rect 5798 43872 5854 43928
rect 5922 43872 5978 43928
rect 6046 43872 6102 43928
rect 6170 43872 6226 43928
rect 6294 43872 6350 43928
rect 6418 43872 6474 43928
rect 6542 43872 6598 43928
rect 6666 43872 6722 43928
rect 6790 43872 6846 43928
rect 6914 43872 6970 43928
rect 7038 43872 7094 43928
rect 5178 43748 5234 43804
rect 5302 43748 5358 43804
rect 5426 43748 5482 43804
rect 5550 43748 5606 43804
rect 5674 43748 5730 43804
rect 5798 43748 5854 43804
rect 5922 43748 5978 43804
rect 6046 43748 6102 43804
rect 6170 43748 6226 43804
rect 6294 43748 6350 43804
rect 6418 43748 6474 43804
rect 6542 43748 6598 43804
rect 6666 43748 6722 43804
rect 6790 43748 6846 43804
rect 6914 43748 6970 43804
rect 7038 43748 7094 43804
rect 5178 43624 5234 43680
rect 5302 43624 5358 43680
rect 5426 43624 5482 43680
rect 5550 43624 5606 43680
rect 5674 43624 5730 43680
rect 5798 43624 5854 43680
rect 5922 43624 5978 43680
rect 6046 43624 6102 43680
rect 6170 43624 6226 43680
rect 6294 43624 6350 43680
rect 6418 43624 6474 43680
rect 6542 43624 6598 43680
rect 6666 43624 6722 43680
rect 6790 43624 6846 43680
rect 6914 43624 6970 43680
rect 7038 43624 7094 43680
rect 5178 43500 5234 43556
rect 5302 43500 5358 43556
rect 5426 43500 5482 43556
rect 5550 43500 5606 43556
rect 5674 43500 5730 43556
rect 5798 43500 5854 43556
rect 5922 43500 5978 43556
rect 6046 43500 6102 43556
rect 6170 43500 6226 43556
rect 6294 43500 6350 43556
rect 6418 43500 6474 43556
rect 6542 43500 6598 43556
rect 6666 43500 6722 43556
rect 6790 43500 6846 43556
rect 6914 43500 6970 43556
rect 7038 43500 7094 43556
rect 5178 43376 5234 43432
rect 5302 43376 5358 43432
rect 5426 43376 5482 43432
rect 5550 43376 5606 43432
rect 5674 43376 5730 43432
rect 5798 43376 5854 43432
rect 5922 43376 5978 43432
rect 6046 43376 6102 43432
rect 6170 43376 6226 43432
rect 6294 43376 6350 43432
rect 6418 43376 6474 43432
rect 6542 43376 6598 43432
rect 6666 43376 6722 43432
rect 6790 43376 6846 43432
rect 6914 43376 6970 43432
rect 7038 43376 7094 43432
rect 5178 43252 5234 43308
rect 5302 43252 5358 43308
rect 5426 43252 5482 43308
rect 5550 43252 5606 43308
rect 5674 43252 5730 43308
rect 5798 43252 5854 43308
rect 5922 43252 5978 43308
rect 6046 43252 6102 43308
rect 6170 43252 6226 43308
rect 6294 43252 6350 43308
rect 6418 43252 6474 43308
rect 6542 43252 6598 43308
rect 6666 43252 6722 43308
rect 6790 43252 6846 43308
rect 6914 43252 6970 43308
rect 7038 43252 7094 43308
rect 7884 44492 7940 44548
rect 8008 44492 8064 44548
rect 8132 44492 8188 44548
rect 8256 44492 8312 44548
rect 8380 44492 8436 44548
rect 8504 44492 8560 44548
rect 8628 44492 8684 44548
rect 8752 44492 8808 44548
rect 8876 44492 8932 44548
rect 9000 44492 9056 44548
rect 9124 44492 9180 44548
rect 9248 44492 9304 44548
rect 9372 44492 9428 44548
rect 9496 44492 9552 44548
rect 9620 44492 9676 44548
rect 9744 44492 9800 44548
rect 7884 44368 7940 44424
rect 8008 44368 8064 44424
rect 8132 44368 8188 44424
rect 8256 44368 8312 44424
rect 8380 44368 8436 44424
rect 8504 44368 8560 44424
rect 8628 44368 8684 44424
rect 8752 44368 8808 44424
rect 8876 44368 8932 44424
rect 9000 44368 9056 44424
rect 9124 44368 9180 44424
rect 9248 44368 9304 44424
rect 9372 44368 9428 44424
rect 9496 44368 9552 44424
rect 9620 44368 9676 44424
rect 9744 44368 9800 44424
rect 7884 44244 7940 44300
rect 8008 44244 8064 44300
rect 8132 44244 8188 44300
rect 8256 44244 8312 44300
rect 8380 44244 8436 44300
rect 8504 44244 8560 44300
rect 8628 44244 8684 44300
rect 8752 44244 8808 44300
rect 8876 44244 8932 44300
rect 9000 44244 9056 44300
rect 9124 44244 9180 44300
rect 9248 44244 9304 44300
rect 9372 44244 9428 44300
rect 9496 44244 9552 44300
rect 9620 44244 9676 44300
rect 9744 44244 9800 44300
rect 7884 44120 7940 44176
rect 8008 44120 8064 44176
rect 8132 44120 8188 44176
rect 8256 44120 8312 44176
rect 8380 44120 8436 44176
rect 8504 44120 8560 44176
rect 8628 44120 8684 44176
rect 8752 44120 8808 44176
rect 8876 44120 8932 44176
rect 9000 44120 9056 44176
rect 9124 44120 9180 44176
rect 9248 44120 9304 44176
rect 9372 44120 9428 44176
rect 9496 44120 9552 44176
rect 9620 44120 9676 44176
rect 9744 44120 9800 44176
rect 7884 43996 7940 44052
rect 8008 43996 8064 44052
rect 8132 43996 8188 44052
rect 8256 43996 8312 44052
rect 8380 43996 8436 44052
rect 8504 43996 8560 44052
rect 8628 43996 8684 44052
rect 8752 43996 8808 44052
rect 8876 43996 8932 44052
rect 9000 43996 9056 44052
rect 9124 43996 9180 44052
rect 9248 43996 9304 44052
rect 9372 43996 9428 44052
rect 9496 43996 9552 44052
rect 9620 43996 9676 44052
rect 9744 43996 9800 44052
rect 7884 43872 7940 43928
rect 8008 43872 8064 43928
rect 8132 43872 8188 43928
rect 8256 43872 8312 43928
rect 8380 43872 8436 43928
rect 8504 43872 8560 43928
rect 8628 43872 8684 43928
rect 8752 43872 8808 43928
rect 8876 43872 8932 43928
rect 9000 43872 9056 43928
rect 9124 43872 9180 43928
rect 9248 43872 9304 43928
rect 9372 43872 9428 43928
rect 9496 43872 9552 43928
rect 9620 43872 9676 43928
rect 9744 43872 9800 43928
rect 7884 43748 7940 43804
rect 8008 43748 8064 43804
rect 8132 43748 8188 43804
rect 8256 43748 8312 43804
rect 8380 43748 8436 43804
rect 8504 43748 8560 43804
rect 8628 43748 8684 43804
rect 8752 43748 8808 43804
rect 8876 43748 8932 43804
rect 9000 43748 9056 43804
rect 9124 43748 9180 43804
rect 9248 43748 9304 43804
rect 9372 43748 9428 43804
rect 9496 43748 9552 43804
rect 9620 43748 9676 43804
rect 9744 43748 9800 43804
rect 7884 43624 7940 43680
rect 8008 43624 8064 43680
rect 8132 43624 8188 43680
rect 8256 43624 8312 43680
rect 8380 43624 8436 43680
rect 8504 43624 8560 43680
rect 8628 43624 8684 43680
rect 8752 43624 8808 43680
rect 8876 43624 8932 43680
rect 9000 43624 9056 43680
rect 9124 43624 9180 43680
rect 9248 43624 9304 43680
rect 9372 43624 9428 43680
rect 9496 43624 9552 43680
rect 9620 43624 9676 43680
rect 9744 43624 9800 43680
rect 7884 43500 7940 43556
rect 8008 43500 8064 43556
rect 8132 43500 8188 43556
rect 8256 43500 8312 43556
rect 8380 43500 8436 43556
rect 8504 43500 8560 43556
rect 8628 43500 8684 43556
rect 8752 43500 8808 43556
rect 8876 43500 8932 43556
rect 9000 43500 9056 43556
rect 9124 43500 9180 43556
rect 9248 43500 9304 43556
rect 9372 43500 9428 43556
rect 9496 43500 9552 43556
rect 9620 43500 9676 43556
rect 9744 43500 9800 43556
rect 7884 43376 7940 43432
rect 8008 43376 8064 43432
rect 8132 43376 8188 43432
rect 8256 43376 8312 43432
rect 8380 43376 8436 43432
rect 8504 43376 8560 43432
rect 8628 43376 8684 43432
rect 8752 43376 8808 43432
rect 8876 43376 8932 43432
rect 9000 43376 9056 43432
rect 9124 43376 9180 43432
rect 9248 43376 9304 43432
rect 9372 43376 9428 43432
rect 9496 43376 9552 43432
rect 9620 43376 9676 43432
rect 9744 43376 9800 43432
rect 7884 43252 7940 43308
rect 8008 43252 8064 43308
rect 8132 43252 8188 43308
rect 8256 43252 8312 43308
rect 8380 43252 8436 43308
rect 8504 43252 8560 43308
rect 8628 43252 8684 43308
rect 8752 43252 8808 43308
rect 8876 43252 8932 43308
rect 9000 43252 9056 43308
rect 9124 43252 9180 43308
rect 9248 43252 9304 43308
rect 9372 43252 9428 43308
rect 9496 43252 9552 43308
rect 9620 43252 9676 43308
rect 9744 43252 9800 43308
rect 10254 44492 10310 44548
rect 10378 44492 10434 44548
rect 10502 44492 10558 44548
rect 10626 44492 10682 44548
rect 10750 44492 10806 44548
rect 10874 44492 10930 44548
rect 10998 44492 11054 44548
rect 11122 44492 11178 44548
rect 11246 44492 11302 44548
rect 11370 44492 11426 44548
rect 11494 44492 11550 44548
rect 11618 44492 11674 44548
rect 11742 44492 11798 44548
rect 11866 44492 11922 44548
rect 11990 44492 12046 44548
rect 12114 44492 12170 44548
rect 10254 44368 10310 44424
rect 10378 44368 10434 44424
rect 10502 44368 10558 44424
rect 10626 44368 10682 44424
rect 10750 44368 10806 44424
rect 10874 44368 10930 44424
rect 10998 44368 11054 44424
rect 11122 44368 11178 44424
rect 11246 44368 11302 44424
rect 11370 44368 11426 44424
rect 11494 44368 11550 44424
rect 11618 44368 11674 44424
rect 11742 44368 11798 44424
rect 11866 44368 11922 44424
rect 11990 44368 12046 44424
rect 12114 44368 12170 44424
rect 10254 44244 10310 44300
rect 10378 44244 10434 44300
rect 10502 44244 10558 44300
rect 10626 44244 10682 44300
rect 10750 44244 10806 44300
rect 10874 44244 10930 44300
rect 10998 44244 11054 44300
rect 11122 44244 11178 44300
rect 11246 44244 11302 44300
rect 11370 44244 11426 44300
rect 11494 44244 11550 44300
rect 11618 44244 11674 44300
rect 11742 44244 11798 44300
rect 11866 44244 11922 44300
rect 11990 44244 12046 44300
rect 12114 44244 12170 44300
rect 10254 44120 10310 44176
rect 10378 44120 10434 44176
rect 10502 44120 10558 44176
rect 10626 44120 10682 44176
rect 10750 44120 10806 44176
rect 10874 44120 10930 44176
rect 10998 44120 11054 44176
rect 11122 44120 11178 44176
rect 11246 44120 11302 44176
rect 11370 44120 11426 44176
rect 11494 44120 11550 44176
rect 11618 44120 11674 44176
rect 11742 44120 11798 44176
rect 11866 44120 11922 44176
rect 11990 44120 12046 44176
rect 12114 44120 12170 44176
rect 10254 43996 10310 44052
rect 10378 43996 10434 44052
rect 10502 43996 10558 44052
rect 10626 43996 10682 44052
rect 10750 43996 10806 44052
rect 10874 43996 10930 44052
rect 10998 43996 11054 44052
rect 11122 43996 11178 44052
rect 11246 43996 11302 44052
rect 11370 43996 11426 44052
rect 11494 43996 11550 44052
rect 11618 43996 11674 44052
rect 11742 43996 11798 44052
rect 11866 43996 11922 44052
rect 11990 43996 12046 44052
rect 12114 43996 12170 44052
rect 10254 43872 10310 43928
rect 10378 43872 10434 43928
rect 10502 43872 10558 43928
rect 10626 43872 10682 43928
rect 10750 43872 10806 43928
rect 10874 43872 10930 43928
rect 10998 43872 11054 43928
rect 11122 43872 11178 43928
rect 11246 43872 11302 43928
rect 11370 43872 11426 43928
rect 11494 43872 11550 43928
rect 11618 43872 11674 43928
rect 11742 43872 11798 43928
rect 11866 43872 11922 43928
rect 11990 43872 12046 43928
rect 12114 43872 12170 43928
rect 10254 43748 10310 43804
rect 10378 43748 10434 43804
rect 10502 43748 10558 43804
rect 10626 43748 10682 43804
rect 10750 43748 10806 43804
rect 10874 43748 10930 43804
rect 10998 43748 11054 43804
rect 11122 43748 11178 43804
rect 11246 43748 11302 43804
rect 11370 43748 11426 43804
rect 11494 43748 11550 43804
rect 11618 43748 11674 43804
rect 11742 43748 11798 43804
rect 11866 43748 11922 43804
rect 11990 43748 12046 43804
rect 12114 43748 12170 43804
rect 10254 43624 10310 43680
rect 10378 43624 10434 43680
rect 10502 43624 10558 43680
rect 10626 43624 10682 43680
rect 10750 43624 10806 43680
rect 10874 43624 10930 43680
rect 10998 43624 11054 43680
rect 11122 43624 11178 43680
rect 11246 43624 11302 43680
rect 11370 43624 11426 43680
rect 11494 43624 11550 43680
rect 11618 43624 11674 43680
rect 11742 43624 11798 43680
rect 11866 43624 11922 43680
rect 11990 43624 12046 43680
rect 12114 43624 12170 43680
rect 10254 43500 10310 43556
rect 10378 43500 10434 43556
rect 10502 43500 10558 43556
rect 10626 43500 10682 43556
rect 10750 43500 10806 43556
rect 10874 43500 10930 43556
rect 10998 43500 11054 43556
rect 11122 43500 11178 43556
rect 11246 43500 11302 43556
rect 11370 43500 11426 43556
rect 11494 43500 11550 43556
rect 11618 43500 11674 43556
rect 11742 43500 11798 43556
rect 11866 43500 11922 43556
rect 11990 43500 12046 43556
rect 12114 43500 12170 43556
rect 10254 43376 10310 43432
rect 10378 43376 10434 43432
rect 10502 43376 10558 43432
rect 10626 43376 10682 43432
rect 10750 43376 10806 43432
rect 10874 43376 10930 43432
rect 10998 43376 11054 43432
rect 11122 43376 11178 43432
rect 11246 43376 11302 43432
rect 11370 43376 11426 43432
rect 11494 43376 11550 43432
rect 11618 43376 11674 43432
rect 11742 43376 11798 43432
rect 11866 43376 11922 43432
rect 11990 43376 12046 43432
rect 12114 43376 12170 43432
rect 10254 43252 10310 43308
rect 10378 43252 10434 43308
rect 10502 43252 10558 43308
rect 10626 43252 10682 43308
rect 10750 43252 10806 43308
rect 10874 43252 10930 43308
rect 10998 43252 11054 43308
rect 11122 43252 11178 43308
rect 11246 43252 11302 43308
rect 11370 43252 11426 43308
rect 11494 43252 11550 43308
rect 11618 43252 11674 43308
rect 11742 43252 11798 43308
rect 11866 43252 11922 43308
rect 11990 43252 12046 43308
rect 12114 43252 12170 43308
rect 12871 44492 12927 44548
rect 12995 44492 13051 44548
rect 13119 44492 13175 44548
rect 13243 44492 13299 44548
rect 13367 44492 13423 44548
rect 13491 44492 13547 44548
rect 13615 44492 13671 44548
rect 13739 44492 13795 44548
rect 13863 44492 13919 44548
rect 13987 44492 14043 44548
rect 14111 44492 14167 44548
rect 14235 44492 14291 44548
rect 14359 44492 14415 44548
rect 14483 44492 14539 44548
rect 14607 44492 14663 44548
rect 12871 44368 12927 44424
rect 12995 44368 13051 44424
rect 13119 44368 13175 44424
rect 13243 44368 13299 44424
rect 13367 44368 13423 44424
rect 13491 44368 13547 44424
rect 13615 44368 13671 44424
rect 13739 44368 13795 44424
rect 13863 44368 13919 44424
rect 13987 44368 14043 44424
rect 14111 44368 14167 44424
rect 14235 44368 14291 44424
rect 14359 44368 14415 44424
rect 14483 44368 14539 44424
rect 14607 44368 14663 44424
rect 12871 44244 12927 44300
rect 12995 44244 13051 44300
rect 13119 44244 13175 44300
rect 13243 44244 13299 44300
rect 13367 44244 13423 44300
rect 13491 44244 13547 44300
rect 13615 44244 13671 44300
rect 13739 44244 13795 44300
rect 13863 44244 13919 44300
rect 13987 44244 14043 44300
rect 14111 44244 14167 44300
rect 14235 44244 14291 44300
rect 14359 44244 14415 44300
rect 14483 44244 14539 44300
rect 14607 44244 14663 44300
rect 12871 44120 12927 44176
rect 12995 44120 13051 44176
rect 13119 44120 13175 44176
rect 13243 44120 13299 44176
rect 13367 44120 13423 44176
rect 13491 44120 13547 44176
rect 13615 44120 13671 44176
rect 13739 44120 13795 44176
rect 13863 44120 13919 44176
rect 13987 44120 14043 44176
rect 14111 44120 14167 44176
rect 14235 44120 14291 44176
rect 14359 44120 14415 44176
rect 14483 44120 14539 44176
rect 14607 44120 14663 44176
rect 12871 43996 12927 44052
rect 12995 43996 13051 44052
rect 13119 43996 13175 44052
rect 13243 43996 13299 44052
rect 13367 43996 13423 44052
rect 13491 43996 13547 44052
rect 13615 43996 13671 44052
rect 13739 43996 13795 44052
rect 13863 43996 13919 44052
rect 13987 43996 14043 44052
rect 14111 43996 14167 44052
rect 14235 43996 14291 44052
rect 14359 43996 14415 44052
rect 14483 43996 14539 44052
rect 14607 43996 14663 44052
rect 12871 43872 12927 43928
rect 12995 43872 13051 43928
rect 13119 43872 13175 43928
rect 13243 43872 13299 43928
rect 13367 43872 13423 43928
rect 13491 43872 13547 43928
rect 13615 43872 13671 43928
rect 13739 43872 13795 43928
rect 13863 43872 13919 43928
rect 13987 43872 14043 43928
rect 14111 43872 14167 43928
rect 14235 43872 14291 43928
rect 14359 43872 14415 43928
rect 14483 43872 14539 43928
rect 14607 43872 14663 43928
rect 12871 43748 12927 43804
rect 12995 43748 13051 43804
rect 13119 43748 13175 43804
rect 13243 43748 13299 43804
rect 13367 43748 13423 43804
rect 13491 43748 13547 43804
rect 13615 43748 13671 43804
rect 13739 43748 13795 43804
rect 13863 43748 13919 43804
rect 13987 43748 14043 43804
rect 14111 43748 14167 43804
rect 14235 43748 14291 43804
rect 14359 43748 14415 43804
rect 14483 43748 14539 43804
rect 14607 43748 14663 43804
rect 12871 43624 12927 43680
rect 12995 43624 13051 43680
rect 13119 43624 13175 43680
rect 13243 43624 13299 43680
rect 13367 43624 13423 43680
rect 13491 43624 13547 43680
rect 13615 43624 13671 43680
rect 13739 43624 13795 43680
rect 13863 43624 13919 43680
rect 13987 43624 14043 43680
rect 14111 43624 14167 43680
rect 14235 43624 14291 43680
rect 14359 43624 14415 43680
rect 14483 43624 14539 43680
rect 14607 43624 14663 43680
rect 12871 43500 12927 43556
rect 12995 43500 13051 43556
rect 13119 43500 13175 43556
rect 13243 43500 13299 43556
rect 13367 43500 13423 43556
rect 13491 43500 13547 43556
rect 13615 43500 13671 43556
rect 13739 43500 13795 43556
rect 13863 43500 13919 43556
rect 13987 43500 14043 43556
rect 14111 43500 14167 43556
rect 14235 43500 14291 43556
rect 14359 43500 14415 43556
rect 14483 43500 14539 43556
rect 14607 43500 14663 43556
rect 12871 43376 12927 43432
rect 12995 43376 13051 43432
rect 13119 43376 13175 43432
rect 13243 43376 13299 43432
rect 13367 43376 13423 43432
rect 13491 43376 13547 43432
rect 13615 43376 13671 43432
rect 13739 43376 13795 43432
rect 13863 43376 13919 43432
rect 13987 43376 14043 43432
rect 14111 43376 14167 43432
rect 14235 43376 14291 43432
rect 14359 43376 14415 43432
rect 14483 43376 14539 43432
rect 14607 43376 14663 43432
rect 12871 43252 12927 43308
rect 12995 43252 13051 43308
rect 13119 43252 13175 43308
rect 13243 43252 13299 43308
rect 13367 43252 13423 43308
rect 13491 43252 13547 43308
rect 13615 43252 13671 43308
rect 13739 43252 13795 43308
rect 13863 43252 13919 43308
rect 13987 43252 14043 43308
rect 14111 43252 14167 43308
rect 14235 43252 14291 43308
rect 14359 43252 14415 43308
rect 14483 43252 14539 43308
rect 14607 43252 14663 43308
rect 2808 42892 2864 42948
rect 2932 42892 2988 42948
rect 3056 42892 3112 42948
rect 3180 42892 3236 42948
rect 3304 42892 3360 42948
rect 3428 42892 3484 42948
rect 3552 42892 3608 42948
rect 3676 42892 3732 42948
rect 3800 42892 3856 42948
rect 3924 42892 3980 42948
rect 4048 42892 4104 42948
rect 4172 42892 4228 42948
rect 4296 42892 4352 42948
rect 4420 42892 4476 42948
rect 4544 42892 4600 42948
rect 4668 42892 4724 42948
rect 2808 42768 2864 42824
rect 2932 42768 2988 42824
rect 3056 42768 3112 42824
rect 3180 42768 3236 42824
rect 3304 42768 3360 42824
rect 3428 42768 3484 42824
rect 3552 42768 3608 42824
rect 3676 42768 3732 42824
rect 3800 42768 3856 42824
rect 3924 42768 3980 42824
rect 4048 42768 4104 42824
rect 4172 42768 4228 42824
rect 4296 42768 4352 42824
rect 4420 42768 4476 42824
rect 4544 42768 4600 42824
rect 4668 42768 4724 42824
rect 2808 42644 2864 42700
rect 2932 42644 2988 42700
rect 3056 42644 3112 42700
rect 3180 42644 3236 42700
rect 3304 42644 3360 42700
rect 3428 42644 3484 42700
rect 3552 42644 3608 42700
rect 3676 42644 3732 42700
rect 3800 42644 3856 42700
rect 3924 42644 3980 42700
rect 4048 42644 4104 42700
rect 4172 42644 4228 42700
rect 4296 42644 4352 42700
rect 4420 42644 4476 42700
rect 4544 42644 4600 42700
rect 4668 42644 4724 42700
rect 2808 42520 2864 42576
rect 2932 42520 2988 42576
rect 3056 42520 3112 42576
rect 3180 42520 3236 42576
rect 3304 42520 3360 42576
rect 3428 42520 3484 42576
rect 3552 42520 3608 42576
rect 3676 42520 3732 42576
rect 3800 42520 3856 42576
rect 3924 42520 3980 42576
rect 4048 42520 4104 42576
rect 4172 42520 4228 42576
rect 4296 42520 4352 42576
rect 4420 42520 4476 42576
rect 4544 42520 4600 42576
rect 4668 42520 4724 42576
rect 2808 42396 2864 42452
rect 2932 42396 2988 42452
rect 3056 42396 3112 42452
rect 3180 42396 3236 42452
rect 3304 42396 3360 42452
rect 3428 42396 3484 42452
rect 3552 42396 3608 42452
rect 3676 42396 3732 42452
rect 3800 42396 3856 42452
rect 3924 42396 3980 42452
rect 4048 42396 4104 42452
rect 4172 42396 4228 42452
rect 4296 42396 4352 42452
rect 4420 42396 4476 42452
rect 4544 42396 4600 42452
rect 4668 42396 4724 42452
rect 2808 42272 2864 42328
rect 2932 42272 2988 42328
rect 3056 42272 3112 42328
rect 3180 42272 3236 42328
rect 3304 42272 3360 42328
rect 3428 42272 3484 42328
rect 3552 42272 3608 42328
rect 3676 42272 3732 42328
rect 3800 42272 3856 42328
rect 3924 42272 3980 42328
rect 4048 42272 4104 42328
rect 4172 42272 4228 42328
rect 4296 42272 4352 42328
rect 4420 42272 4476 42328
rect 4544 42272 4600 42328
rect 4668 42272 4724 42328
rect 2808 42148 2864 42204
rect 2932 42148 2988 42204
rect 3056 42148 3112 42204
rect 3180 42148 3236 42204
rect 3304 42148 3360 42204
rect 3428 42148 3484 42204
rect 3552 42148 3608 42204
rect 3676 42148 3732 42204
rect 3800 42148 3856 42204
rect 3924 42148 3980 42204
rect 4048 42148 4104 42204
rect 4172 42148 4228 42204
rect 4296 42148 4352 42204
rect 4420 42148 4476 42204
rect 4544 42148 4600 42204
rect 4668 42148 4724 42204
rect 2808 42024 2864 42080
rect 2932 42024 2988 42080
rect 3056 42024 3112 42080
rect 3180 42024 3236 42080
rect 3304 42024 3360 42080
rect 3428 42024 3484 42080
rect 3552 42024 3608 42080
rect 3676 42024 3732 42080
rect 3800 42024 3856 42080
rect 3924 42024 3980 42080
rect 4048 42024 4104 42080
rect 4172 42024 4228 42080
rect 4296 42024 4352 42080
rect 4420 42024 4476 42080
rect 4544 42024 4600 42080
rect 4668 42024 4724 42080
rect 2808 41900 2864 41956
rect 2932 41900 2988 41956
rect 3056 41900 3112 41956
rect 3180 41900 3236 41956
rect 3304 41900 3360 41956
rect 3428 41900 3484 41956
rect 3552 41900 3608 41956
rect 3676 41900 3732 41956
rect 3800 41900 3856 41956
rect 3924 41900 3980 41956
rect 4048 41900 4104 41956
rect 4172 41900 4228 41956
rect 4296 41900 4352 41956
rect 4420 41900 4476 41956
rect 4544 41900 4600 41956
rect 4668 41900 4724 41956
rect 2808 41776 2864 41832
rect 2932 41776 2988 41832
rect 3056 41776 3112 41832
rect 3180 41776 3236 41832
rect 3304 41776 3360 41832
rect 3428 41776 3484 41832
rect 3552 41776 3608 41832
rect 3676 41776 3732 41832
rect 3800 41776 3856 41832
rect 3924 41776 3980 41832
rect 4048 41776 4104 41832
rect 4172 41776 4228 41832
rect 4296 41776 4352 41832
rect 4420 41776 4476 41832
rect 4544 41776 4600 41832
rect 4668 41776 4724 41832
rect 2808 41652 2864 41708
rect 2932 41652 2988 41708
rect 3056 41652 3112 41708
rect 3180 41652 3236 41708
rect 3304 41652 3360 41708
rect 3428 41652 3484 41708
rect 3552 41652 3608 41708
rect 3676 41652 3732 41708
rect 3800 41652 3856 41708
rect 3924 41652 3980 41708
rect 4048 41652 4104 41708
rect 4172 41652 4228 41708
rect 4296 41652 4352 41708
rect 4420 41652 4476 41708
rect 4544 41652 4600 41708
rect 4668 41652 4724 41708
rect 5178 42892 5234 42948
rect 5302 42892 5358 42948
rect 5426 42892 5482 42948
rect 5550 42892 5606 42948
rect 5674 42892 5730 42948
rect 5798 42892 5854 42948
rect 5922 42892 5978 42948
rect 6046 42892 6102 42948
rect 6170 42892 6226 42948
rect 6294 42892 6350 42948
rect 6418 42892 6474 42948
rect 6542 42892 6598 42948
rect 6666 42892 6722 42948
rect 6790 42892 6846 42948
rect 6914 42892 6970 42948
rect 7038 42892 7094 42948
rect 5178 42768 5234 42824
rect 5302 42768 5358 42824
rect 5426 42768 5482 42824
rect 5550 42768 5606 42824
rect 5674 42768 5730 42824
rect 5798 42768 5854 42824
rect 5922 42768 5978 42824
rect 6046 42768 6102 42824
rect 6170 42768 6226 42824
rect 6294 42768 6350 42824
rect 6418 42768 6474 42824
rect 6542 42768 6598 42824
rect 6666 42768 6722 42824
rect 6790 42768 6846 42824
rect 6914 42768 6970 42824
rect 7038 42768 7094 42824
rect 5178 42644 5234 42700
rect 5302 42644 5358 42700
rect 5426 42644 5482 42700
rect 5550 42644 5606 42700
rect 5674 42644 5730 42700
rect 5798 42644 5854 42700
rect 5922 42644 5978 42700
rect 6046 42644 6102 42700
rect 6170 42644 6226 42700
rect 6294 42644 6350 42700
rect 6418 42644 6474 42700
rect 6542 42644 6598 42700
rect 6666 42644 6722 42700
rect 6790 42644 6846 42700
rect 6914 42644 6970 42700
rect 7038 42644 7094 42700
rect 5178 42520 5234 42576
rect 5302 42520 5358 42576
rect 5426 42520 5482 42576
rect 5550 42520 5606 42576
rect 5674 42520 5730 42576
rect 5798 42520 5854 42576
rect 5922 42520 5978 42576
rect 6046 42520 6102 42576
rect 6170 42520 6226 42576
rect 6294 42520 6350 42576
rect 6418 42520 6474 42576
rect 6542 42520 6598 42576
rect 6666 42520 6722 42576
rect 6790 42520 6846 42576
rect 6914 42520 6970 42576
rect 7038 42520 7094 42576
rect 5178 42396 5234 42452
rect 5302 42396 5358 42452
rect 5426 42396 5482 42452
rect 5550 42396 5606 42452
rect 5674 42396 5730 42452
rect 5798 42396 5854 42452
rect 5922 42396 5978 42452
rect 6046 42396 6102 42452
rect 6170 42396 6226 42452
rect 6294 42396 6350 42452
rect 6418 42396 6474 42452
rect 6542 42396 6598 42452
rect 6666 42396 6722 42452
rect 6790 42396 6846 42452
rect 6914 42396 6970 42452
rect 7038 42396 7094 42452
rect 5178 42272 5234 42328
rect 5302 42272 5358 42328
rect 5426 42272 5482 42328
rect 5550 42272 5606 42328
rect 5674 42272 5730 42328
rect 5798 42272 5854 42328
rect 5922 42272 5978 42328
rect 6046 42272 6102 42328
rect 6170 42272 6226 42328
rect 6294 42272 6350 42328
rect 6418 42272 6474 42328
rect 6542 42272 6598 42328
rect 6666 42272 6722 42328
rect 6790 42272 6846 42328
rect 6914 42272 6970 42328
rect 7038 42272 7094 42328
rect 5178 42148 5234 42204
rect 5302 42148 5358 42204
rect 5426 42148 5482 42204
rect 5550 42148 5606 42204
rect 5674 42148 5730 42204
rect 5798 42148 5854 42204
rect 5922 42148 5978 42204
rect 6046 42148 6102 42204
rect 6170 42148 6226 42204
rect 6294 42148 6350 42204
rect 6418 42148 6474 42204
rect 6542 42148 6598 42204
rect 6666 42148 6722 42204
rect 6790 42148 6846 42204
rect 6914 42148 6970 42204
rect 7038 42148 7094 42204
rect 5178 42024 5234 42080
rect 5302 42024 5358 42080
rect 5426 42024 5482 42080
rect 5550 42024 5606 42080
rect 5674 42024 5730 42080
rect 5798 42024 5854 42080
rect 5922 42024 5978 42080
rect 6046 42024 6102 42080
rect 6170 42024 6226 42080
rect 6294 42024 6350 42080
rect 6418 42024 6474 42080
rect 6542 42024 6598 42080
rect 6666 42024 6722 42080
rect 6790 42024 6846 42080
rect 6914 42024 6970 42080
rect 7038 42024 7094 42080
rect 5178 41900 5234 41956
rect 5302 41900 5358 41956
rect 5426 41900 5482 41956
rect 5550 41900 5606 41956
rect 5674 41900 5730 41956
rect 5798 41900 5854 41956
rect 5922 41900 5978 41956
rect 6046 41900 6102 41956
rect 6170 41900 6226 41956
rect 6294 41900 6350 41956
rect 6418 41900 6474 41956
rect 6542 41900 6598 41956
rect 6666 41900 6722 41956
rect 6790 41900 6846 41956
rect 6914 41900 6970 41956
rect 7038 41900 7094 41956
rect 5178 41776 5234 41832
rect 5302 41776 5358 41832
rect 5426 41776 5482 41832
rect 5550 41776 5606 41832
rect 5674 41776 5730 41832
rect 5798 41776 5854 41832
rect 5922 41776 5978 41832
rect 6046 41776 6102 41832
rect 6170 41776 6226 41832
rect 6294 41776 6350 41832
rect 6418 41776 6474 41832
rect 6542 41776 6598 41832
rect 6666 41776 6722 41832
rect 6790 41776 6846 41832
rect 6914 41776 6970 41832
rect 7038 41776 7094 41832
rect 5178 41652 5234 41708
rect 5302 41652 5358 41708
rect 5426 41652 5482 41708
rect 5550 41652 5606 41708
rect 5674 41652 5730 41708
rect 5798 41652 5854 41708
rect 5922 41652 5978 41708
rect 6046 41652 6102 41708
rect 6170 41652 6226 41708
rect 6294 41652 6350 41708
rect 6418 41652 6474 41708
rect 6542 41652 6598 41708
rect 6666 41652 6722 41708
rect 6790 41652 6846 41708
rect 6914 41652 6970 41708
rect 7038 41652 7094 41708
rect 7884 42892 7940 42948
rect 8008 42892 8064 42948
rect 8132 42892 8188 42948
rect 8256 42892 8312 42948
rect 8380 42892 8436 42948
rect 8504 42892 8560 42948
rect 8628 42892 8684 42948
rect 8752 42892 8808 42948
rect 8876 42892 8932 42948
rect 9000 42892 9056 42948
rect 9124 42892 9180 42948
rect 9248 42892 9304 42948
rect 9372 42892 9428 42948
rect 9496 42892 9552 42948
rect 9620 42892 9676 42948
rect 9744 42892 9800 42948
rect 7884 42768 7940 42824
rect 8008 42768 8064 42824
rect 8132 42768 8188 42824
rect 8256 42768 8312 42824
rect 8380 42768 8436 42824
rect 8504 42768 8560 42824
rect 8628 42768 8684 42824
rect 8752 42768 8808 42824
rect 8876 42768 8932 42824
rect 9000 42768 9056 42824
rect 9124 42768 9180 42824
rect 9248 42768 9304 42824
rect 9372 42768 9428 42824
rect 9496 42768 9552 42824
rect 9620 42768 9676 42824
rect 9744 42768 9800 42824
rect 7884 42644 7940 42700
rect 8008 42644 8064 42700
rect 8132 42644 8188 42700
rect 8256 42644 8312 42700
rect 8380 42644 8436 42700
rect 8504 42644 8560 42700
rect 8628 42644 8684 42700
rect 8752 42644 8808 42700
rect 8876 42644 8932 42700
rect 9000 42644 9056 42700
rect 9124 42644 9180 42700
rect 9248 42644 9304 42700
rect 9372 42644 9428 42700
rect 9496 42644 9552 42700
rect 9620 42644 9676 42700
rect 9744 42644 9800 42700
rect 7884 42520 7940 42576
rect 8008 42520 8064 42576
rect 8132 42520 8188 42576
rect 8256 42520 8312 42576
rect 8380 42520 8436 42576
rect 8504 42520 8560 42576
rect 8628 42520 8684 42576
rect 8752 42520 8808 42576
rect 8876 42520 8932 42576
rect 9000 42520 9056 42576
rect 9124 42520 9180 42576
rect 9248 42520 9304 42576
rect 9372 42520 9428 42576
rect 9496 42520 9552 42576
rect 9620 42520 9676 42576
rect 9744 42520 9800 42576
rect 7884 42396 7940 42452
rect 8008 42396 8064 42452
rect 8132 42396 8188 42452
rect 8256 42396 8312 42452
rect 8380 42396 8436 42452
rect 8504 42396 8560 42452
rect 8628 42396 8684 42452
rect 8752 42396 8808 42452
rect 8876 42396 8932 42452
rect 9000 42396 9056 42452
rect 9124 42396 9180 42452
rect 9248 42396 9304 42452
rect 9372 42396 9428 42452
rect 9496 42396 9552 42452
rect 9620 42396 9676 42452
rect 9744 42396 9800 42452
rect 7884 42272 7940 42328
rect 8008 42272 8064 42328
rect 8132 42272 8188 42328
rect 8256 42272 8312 42328
rect 8380 42272 8436 42328
rect 8504 42272 8560 42328
rect 8628 42272 8684 42328
rect 8752 42272 8808 42328
rect 8876 42272 8932 42328
rect 9000 42272 9056 42328
rect 9124 42272 9180 42328
rect 9248 42272 9304 42328
rect 9372 42272 9428 42328
rect 9496 42272 9552 42328
rect 9620 42272 9676 42328
rect 9744 42272 9800 42328
rect 7884 42148 7940 42204
rect 8008 42148 8064 42204
rect 8132 42148 8188 42204
rect 8256 42148 8312 42204
rect 8380 42148 8436 42204
rect 8504 42148 8560 42204
rect 8628 42148 8684 42204
rect 8752 42148 8808 42204
rect 8876 42148 8932 42204
rect 9000 42148 9056 42204
rect 9124 42148 9180 42204
rect 9248 42148 9304 42204
rect 9372 42148 9428 42204
rect 9496 42148 9552 42204
rect 9620 42148 9676 42204
rect 9744 42148 9800 42204
rect 7884 42024 7940 42080
rect 8008 42024 8064 42080
rect 8132 42024 8188 42080
rect 8256 42024 8312 42080
rect 8380 42024 8436 42080
rect 8504 42024 8560 42080
rect 8628 42024 8684 42080
rect 8752 42024 8808 42080
rect 8876 42024 8932 42080
rect 9000 42024 9056 42080
rect 9124 42024 9180 42080
rect 9248 42024 9304 42080
rect 9372 42024 9428 42080
rect 9496 42024 9552 42080
rect 9620 42024 9676 42080
rect 9744 42024 9800 42080
rect 7884 41900 7940 41956
rect 8008 41900 8064 41956
rect 8132 41900 8188 41956
rect 8256 41900 8312 41956
rect 8380 41900 8436 41956
rect 8504 41900 8560 41956
rect 8628 41900 8684 41956
rect 8752 41900 8808 41956
rect 8876 41900 8932 41956
rect 9000 41900 9056 41956
rect 9124 41900 9180 41956
rect 9248 41900 9304 41956
rect 9372 41900 9428 41956
rect 9496 41900 9552 41956
rect 9620 41900 9676 41956
rect 9744 41900 9800 41956
rect 7884 41776 7940 41832
rect 8008 41776 8064 41832
rect 8132 41776 8188 41832
rect 8256 41776 8312 41832
rect 8380 41776 8436 41832
rect 8504 41776 8560 41832
rect 8628 41776 8684 41832
rect 8752 41776 8808 41832
rect 8876 41776 8932 41832
rect 9000 41776 9056 41832
rect 9124 41776 9180 41832
rect 9248 41776 9304 41832
rect 9372 41776 9428 41832
rect 9496 41776 9552 41832
rect 9620 41776 9676 41832
rect 9744 41776 9800 41832
rect 7884 41652 7940 41708
rect 8008 41652 8064 41708
rect 8132 41652 8188 41708
rect 8256 41652 8312 41708
rect 8380 41652 8436 41708
rect 8504 41652 8560 41708
rect 8628 41652 8684 41708
rect 8752 41652 8808 41708
rect 8876 41652 8932 41708
rect 9000 41652 9056 41708
rect 9124 41652 9180 41708
rect 9248 41652 9304 41708
rect 9372 41652 9428 41708
rect 9496 41652 9552 41708
rect 9620 41652 9676 41708
rect 9744 41652 9800 41708
rect 10254 42892 10310 42948
rect 10378 42892 10434 42948
rect 10502 42892 10558 42948
rect 10626 42892 10682 42948
rect 10750 42892 10806 42948
rect 10874 42892 10930 42948
rect 10998 42892 11054 42948
rect 11122 42892 11178 42948
rect 11246 42892 11302 42948
rect 11370 42892 11426 42948
rect 11494 42892 11550 42948
rect 11618 42892 11674 42948
rect 11742 42892 11798 42948
rect 11866 42892 11922 42948
rect 11990 42892 12046 42948
rect 12114 42892 12170 42948
rect 10254 42768 10310 42824
rect 10378 42768 10434 42824
rect 10502 42768 10558 42824
rect 10626 42768 10682 42824
rect 10750 42768 10806 42824
rect 10874 42768 10930 42824
rect 10998 42768 11054 42824
rect 11122 42768 11178 42824
rect 11246 42768 11302 42824
rect 11370 42768 11426 42824
rect 11494 42768 11550 42824
rect 11618 42768 11674 42824
rect 11742 42768 11798 42824
rect 11866 42768 11922 42824
rect 11990 42768 12046 42824
rect 12114 42768 12170 42824
rect 10254 42644 10310 42700
rect 10378 42644 10434 42700
rect 10502 42644 10558 42700
rect 10626 42644 10682 42700
rect 10750 42644 10806 42700
rect 10874 42644 10930 42700
rect 10998 42644 11054 42700
rect 11122 42644 11178 42700
rect 11246 42644 11302 42700
rect 11370 42644 11426 42700
rect 11494 42644 11550 42700
rect 11618 42644 11674 42700
rect 11742 42644 11798 42700
rect 11866 42644 11922 42700
rect 11990 42644 12046 42700
rect 12114 42644 12170 42700
rect 10254 42520 10310 42576
rect 10378 42520 10434 42576
rect 10502 42520 10558 42576
rect 10626 42520 10682 42576
rect 10750 42520 10806 42576
rect 10874 42520 10930 42576
rect 10998 42520 11054 42576
rect 11122 42520 11178 42576
rect 11246 42520 11302 42576
rect 11370 42520 11426 42576
rect 11494 42520 11550 42576
rect 11618 42520 11674 42576
rect 11742 42520 11798 42576
rect 11866 42520 11922 42576
rect 11990 42520 12046 42576
rect 12114 42520 12170 42576
rect 10254 42396 10310 42452
rect 10378 42396 10434 42452
rect 10502 42396 10558 42452
rect 10626 42396 10682 42452
rect 10750 42396 10806 42452
rect 10874 42396 10930 42452
rect 10998 42396 11054 42452
rect 11122 42396 11178 42452
rect 11246 42396 11302 42452
rect 11370 42396 11426 42452
rect 11494 42396 11550 42452
rect 11618 42396 11674 42452
rect 11742 42396 11798 42452
rect 11866 42396 11922 42452
rect 11990 42396 12046 42452
rect 12114 42396 12170 42452
rect 10254 42272 10310 42328
rect 10378 42272 10434 42328
rect 10502 42272 10558 42328
rect 10626 42272 10682 42328
rect 10750 42272 10806 42328
rect 10874 42272 10930 42328
rect 10998 42272 11054 42328
rect 11122 42272 11178 42328
rect 11246 42272 11302 42328
rect 11370 42272 11426 42328
rect 11494 42272 11550 42328
rect 11618 42272 11674 42328
rect 11742 42272 11798 42328
rect 11866 42272 11922 42328
rect 11990 42272 12046 42328
rect 12114 42272 12170 42328
rect 10254 42148 10310 42204
rect 10378 42148 10434 42204
rect 10502 42148 10558 42204
rect 10626 42148 10682 42204
rect 10750 42148 10806 42204
rect 10874 42148 10930 42204
rect 10998 42148 11054 42204
rect 11122 42148 11178 42204
rect 11246 42148 11302 42204
rect 11370 42148 11426 42204
rect 11494 42148 11550 42204
rect 11618 42148 11674 42204
rect 11742 42148 11798 42204
rect 11866 42148 11922 42204
rect 11990 42148 12046 42204
rect 12114 42148 12170 42204
rect 10254 42024 10310 42080
rect 10378 42024 10434 42080
rect 10502 42024 10558 42080
rect 10626 42024 10682 42080
rect 10750 42024 10806 42080
rect 10874 42024 10930 42080
rect 10998 42024 11054 42080
rect 11122 42024 11178 42080
rect 11246 42024 11302 42080
rect 11370 42024 11426 42080
rect 11494 42024 11550 42080
rect 11618 42024 11674 42080
rect 11742 42024 11798 42080
rect 11866 42024 11922 42080
rect 11990 42024 12046 42080
rect 12114 42024 12170 42080
rect 10254 41900 10310 41956
rect 10378 41900 10434 41956
rect 10502 41900 10558 41956
rect 10626 41900 10682 41956
rect 10750 41900 10806 41956
rect 10874 41900 10930 41956
rect 10998 41900 11054 41956
rect 11122 41900 11178 41956
rect 11246 41900 11302 41956
rect 11370 41900 11426 41956
rect 11494 41900 11550 41956
rect 11618 41900 11674 41956
rect 11742 41900 11798 41956
rect 11866 41900 11922 41956
rect 11990 41900 12046 41956
rect 12114 41900 12170 41956
rect 10254 41776 10310 41832
rect 10378 41776 10434 41832
rect 10502 41776 10558 41832
rect 10626 41776 10682 41832
rect 10750 41776 10806 41832
rect 10874 41776 10930 41832
rect 10998 41776 11054 41832
rect 11122 41776 11178 41832
rect 11246 41776 11302 41832
rect 11370 41776 11426 41832
rect 11494 41776 11550 41832
rect 11618 41776 11674 41832
rect 11742 41776 11798 41832
rect 11866 41776 11922 41832
rect 11990 41776 12046 41832
rect 12114 41776 12170 41832
rect 10254 41652 10310 41708
rect 10378 41652 10434 41708
rect 10502 41652 10558 41708
rect 10626 41652 10682 41708
rect 10750 41652 10806 41708
rect 10874 41652 10930 41708
rect 10998 41652 11054 41708
rect 11122 41652 11178 41708
rect 11246 41652 11302 41708
rect 11370 41652 11426 41708
rect 11494 41652 11550 41708
rect 11618 41652 11674 41708
rect 11742 41652 11798 41708
rect 11866 41652 11922 41708
rect 11990 41652 12046 41708
rect 12114 41652 12170 41708
rect 12871 42892 12927 42948
rect 12995 42892 13051 42948
rect 13119 42892 13175 42948
rect 13243 42892 13299 42948
rect 13367 42892 13423 42948
rect 13491 42892 13547 42948
rect 13615 42892 13671 42948
rect 13739 42892 13795 42948
rect 13863 42892 13919 42948
rect 13987 42892 14043 42948
rect 14111 42892 14167 42948
rect 14235 42892 14291 42948
rect 14359 42892 14415 42948
rect 14483 42892 14539 42948
rect 14607 42892 14663 42948
rect 12871 42768 12927 42824
rect 12995 42768 13051 42824
rect 13119 42768 13175 42824
rect 13243 42768 13299 42824
rect 13367 42768 13423 42824
rect 13491 42768 13547 42824
rect 13615 42768 13671 42824
rect 13739 42768 13795 42824
rect 13863 42768 13919 42824
rect 13987 42768 14043 42824
rect 14111 42768 14167 42824
rect 14235 42768 14291 42824
rect 14359 42768 14415 42824
rect 14483 42768 14539 42824
rect 14607 42768 14663 42824
rect 12871 42644 12927 42700
rect 12995 42644 13051 42700
rect 13119 42644 13175 42700
rect 13243 42644 13299 42700
rect 13367 42644 13423 42700
rect 13491 42644 13547 42700
rect 13615 42644 13671 42700
rect 13739 42644 13795 42700
rect 13863 42644 13919 42700
rect 13987 42644 14043 42700
rect 14111 42644 14167 42700
rect 14235 42644 14291 42700
rect 14359 42644 14415 42700
rect 14483 42644 14539 42700
rect 14607 42644 14663 42700
rect 12871 42520 12927 42576
rect 12995 42520 13051 42576
rect 13119 42520 13175 42576
rect 13243 42520 13299 42576
rect 13367 42520 13423 42576
rect 13491 42520 13547 42576
rect 13615 42520 13671 42576
rect 13739 42520 13795 42576
rect 13863 42520 13919 42576
rect 13987 42520 14043 42576
rect 14111 42520 14167 42576
rect 14235 42520 14291 42576
rect 14359 42520 14415 42576
rect 14483 42520 14539 42576
rect 14607 42520 14663 42576
rect 12871 42396 12927 42452
rect 12995 42396 13051 42452
rect 13119 42396 13175 42452
rect 13243 42396 13299 42452
rect 13367 42396 13423 42452
rect 13491 42396 13547 42452
rect 13615 42396 13671 42452
rect 13739 42396 13795 42452
rect 13863 42396 13919 42452
rect 13987 42396 14043 42452
rect 14111 42396 14167 42452
rect 14235 42396 14291 42452
rect 14359 42396 14415 42452
rect 14483 42396 14539 42452
rect 14607 42396 14663 42452
rect 12871 42272 12927 42328
rect 12995 42272 13051 42328
rect 13119 42272 13175 42328
rect 13243 42272 13299 42328
rect 13367 42272 13423 42328
rect 13491 42272 13547 42328
rect 13615 42272 13671 42328
rect 13739 42272 13795 42328
rect 13863 42272 13919 42328
rect 13987 42272 14043 42328
rect 14111 42272 14167 42328
rect 14235 42272 14291 42328
rect 14359 42272 14415 42328
rect 14483 42272 14539 42328
rect 14607 42272 14663 42328
rect 12871 42148 12927 42204
rect 12995 42148 13051 42204
rect 13119 42148 13175 42204
rect 13243 42148 13299 42204
rect 13367 42148 13423 42204
rect 13491 42148 13547 42204
rect 13615 42148 13671 42204
rect 13739 42148 13795 42204
rect 13863 42148 13919 42204
rect 13987 42148 14043 42204
rect 14111 42148 14167 42204
rect 14235 42148 14291 42204
rect 14359 42148 14415 42204
rect 14483 42148 14539 42204
rect 14607 42148 14663 42204
rect 12871 42024 12927 42080
rect 12995 42024 13051 42080
rect 13119 42024 13175 42080
rect 13243 42024 13299 42080
rect 13367 42024 13423 42080
rect 13491 42024 13547 42080
rect 13615 42024 13671 42080
rect 13739 42024 13795 42080
rect 13863 42024 13919 42080
rect 13987 42024 14043 42080
rect 14111 42024 14167 42080
rect 14235 42024 14291 42080
rect 14359 42024 14415 42080
rect 14483 42024 14539 42080
rect 14607 42024 14663 42080
rect 12871 41900 12927 41956
rect 12995 41900 13051 41956
rect 13119 41900 13175 41956
rect 13243 41900 13299 41956
rect 13367 41900 13423 41956
rect 13491 41900 13547 41956
rect 13615 41900 13671 41956
rect 13739 41900 13795 41956
rect 13863 41900 13919 41956
rect 13987 41900 14043 41956
rect 14111 41900 14167 41956
rect 14235 41900 14291 41956
rect 14359 41900 14415 41956
rect 14483 41900 14539 41956
rect 14607 41900 14663 41956
rect 12871 41776 12927 41832
rect 12995 41776 13051 41832
rect 13119 41776 13175 41832
rect 13243 41776 13299 41832
rect 13367 41776 13423 41832
rect 13491 41776 13547 41832
rect 13615 41776 13671 41832
rect 13739 41776 13795 41832
rect 13863 41776 13919 41832
rect 13987 41776 14043 41832
rect 14111 41776 14167 41832
rect 14235 41776 14291 41832
rect 14359 41776 14415 41832
rect 14483 41776 14539 41832
rect 14607 41776 14663 41832
rect 12871 41652 12927 41708
rect 12995 41652 13051 41708
rect 13119 41652 13175 41708
rect 13243 41652 13299 41708
rect 13367 41652 13423 41708
rect 13491 41652 13547 41708
rect 13615 41652 13671 41708
rect 13739 41652 13795 41708
rect 13863 41652 13919 41708
rect 13987 41652 14043 41708
rect 14111 41652 14167 41708
rect 14235 41652 14291 41708
rect 14359 41652 14415 41708
rect 14483 41652 14539 41708
rect 14607 41652 14663 41708
rect 2808 41292 2864 41348
rect 2932 41292 2988 41348
rect 3056 41292 3112 41348
rect 3180 41292 3236 41348
rect 3304 41292 3360 41348
rect 3428 41292 3484 41348
rect 3552 41292 3608 41348
rect 3676 41292 3732 41348
rect 3800 41292 3856 41348
rect 3924 41292 3980 41348
rect 4048 41292 4104 41348
rect 4172 41292 4228 41348
rect 4296 41292 4352 41348
rect 4420 41292 4476 41348
rect 4544 41292 4600 41348
rect 4668 41292 4724 41348
rect 2808 41168 2864 41224
rect 2932 41168 2988 41224
rect 3056 41168 3112 41224
rect 3180 41168 3236 41224
rect 3304 41168 3360 41224
rect 3428 41168 3484 41224
rect 3552 41168 3608 41224
rect 3676 41168 3732 41224
rect 3800 41168 3856 41224
rect 3924 41168 3980 41224
rect 4048 41168 4104 41224
rect 4172 41168 4228 41224
rect 4296 41168 4352 41224
rect 4420 41168 4476 41224
rect 4544 41168 4600 41224
rect 4668 41168 4724 41224
rect 2808 41044 2864 41100
rect 2932 41044 2988 41100
rect 3056 41044 3112 41100
rect 3180 41044 3236 41100
rect 3304 41044 3360 41100
rect 3428 41044 3484 41100
rect 3552 41044 3608 41100
rect 3676 41044 3732 41100
rect 3800 41044 3856 41100
rect 3924 41044 3980 41100
rect 4048 41044 4104 41100
rect 4172 41044 4228 41100
rect 4296 41044 4352 41100
rect 4420 41044 4476 41100
rect 4544 41044 4600 41100
rect 4668 41044 4724 41100
rect 2808 40920 2864 40976
rect 2932 40920 2988 40976
rect 3056 40920 3112 40976
rect 3180 40920 3236 40976
rect 3304 40920 3360 40976
rect 3428 40920 3484 40976
rect 3552 40920 3608 40976
rect 3676 40920 3732 40976
rect 3800 40920 3856 40976
rect 3924 40920 3980 40976
rect 4048 40920 4104 40976
rect 4172 40920 4228 40976
rect 4296 40920 4352 40976
rect 4420 40920 4476 40976
rect 4544 40920 4600 40976
rect 4668 40920 4724 40976
rect 2808 40796 2864 40852
rect 2932 40796 2988 40852
rect 3056 40796 3112 40852
rect 3180 40796 3236 40852
rect 3304 40796 3360 40852
rect 3428 40796 3484 40852
rect 3552 40796 3608 40852
rect 3676 40796 3732 40852
rect 3800 40796 3856 40852
rect 3924 40796 3980 40852
rect 4048 40796 4104 40852
rect 4172 40796 4228 40852
rect 4296 40796 4352 40852
rect 4420 40796 4476 40852
rect 4544 40796 4600 40852
rect 4668 40796 4724 40852
rect 2808 40672 2864 40728
rect 2932 40672 2988 40728
rect 3056 40672 3112 40728
rect 3180 40672 3236 40728
rect 3304 40672 3360 40728
rect 3428 40672 3484 40728
rect 3552 40672 3608 40728
rect 3676 40672 3732 40728
rect 3800 40672 3856 40728
rect 3924 40672 3980 40728
rect 4048 40672 4104 40728
rect 4172 40672 4228 40728
rect 4296 40672 4352 40728
rect 4420 40672 4476 40728
rect 4544 40672 4600 40728
rect 4668 40672 4724 40728
rect 2808 40548 2864 40604
rect 2932 40548 2988 40604
rect 3056 40548 3112 40604
rect 3180 40548 3236 40604
rect 3304 40548 3360 40604
rect 3428 40548 3484 40604
rect 3552 40548 3608 40604
rect 3676 40548 3732 40604
rect 3800 40548 3856 40604
rect 3924 40548 3980 40604
rect 4048 40548 4104 40604
rect 4172 40548 4228 40604
rect 4296 40548 4352 40604
rect 4420 40548 4476 40604
rect 4544 40548 4600 40604
rect 4668 40548 4724 40604
rect 2808 40424 2864 40480
rect 2932 40424 2988 40480
rect 3056 40424 3112 40480
rect 3180 40424 3236 40480
rect 3304 40424 3360 40480
rect 3428 40424 3484 40480
rect 3552 40424 3608 40480
rect 3676 40424 3732 40480
rect 3800 40424 3856 40480
rect 3924 40424 3980 40480
rect 4048 40424 4104 40480
rect 4172 40424 4228 40480
rect 4296 40424 4352 40480
rect 4420 40424 4476 40480
rect 4544 40424 4600 40480
rect 4668 40424 4724 40480
rect 2808 40300 2864 40356
rect 2932 40300 2988 40356
rect 3056 40300 3112 40356
rect 3180 40300 3236 40356
rect 3304 40300 3360 40356
rect 3428 40300 3484 40356
rect 3552 40300 3608 40356
rect 3676 40300 3732 40356
rect 3800 40300 3856 40356
rect 3924 40300 3980 40356
rect 4048 40300 4104 40356
rect 4172 40300 4228 40356
rect 4296 40300 4352 40356
rect 4420 40300 4476 40356
rect 4544 40300 4600 40356
rect 4668 40300 4724 40356
rect 2808 40176 2864 40232
rect 2932 40176 2988 40232
rect 3056 40176 3112 40232
rect 3180 40176 3236 40232
rect 3304 40176 3360 40232
rect 3428 40176 3484 40232
rect 3552 40176 3608 40232
rect 3676 40176 3732 40232
rect 3800 40176 3856 40232
rect 3924 40176 3980 40232
rect 4048 40176 4104 40232
rect 4172 40176 4228 40232
rect 4296 40176 4352 40232
rect 4420 40176 4476 40232
rect 4544 40176 4600 40232
rect 4668 40176 4724 40232
rect 2808 40052 2864 40108
rect 2932 40052 2988 40108
rect 3056 40052 3112 40108
rect 3180 40052 3236 40108
rect 3304 40052 3360 40108
rect 3428 40052 3484 40108
rect 3552 40052 3608 40108
rect 3676 40052 3732 40108
rect 3800 40052 3856 40108
rect 3924 40052 3980 40108
rect 4048 40052 4104 40108
rect 4172 40052 4228 40108
rect 4296 40052 4352 40108
rect 4420 40052 4476 40108
rect 4544 40052 4600 40108
rect 4668 40052 4724 40108
rect 5178 41292 5234 41348
rect 5302 41292 5358 41348
rect 5426 41292 5482 41348
rect 5550 41292 5606 41348
rect 5674 41292 5730 41348
rect 5798 41292 5854 41348
rect 5922 41292 5978 41348
rect 6046 41292 6102 41348
rect 6170 41292 6226 41348
rect 6294 41292 6350 41348
rect 6418 41292 6474 41348
rect 6542 41292 6598 41348
rect 6666 41292 6722 41348
rect 6790 41292 6846 41348
rect 6914 41292 6970 41348
rect 7038 41292 7094 41348
rect 5178 41168 5234 41224
rect 5302 41168 5358 41224
rect 5426 41168 5482 41224
rect 5550 41168 5606 41224
rect 5674 41168 5730 41224
rect 5798 41168 5854 41224
rect 5922 41168 5978 41224
rect 6046 41168 6102 41224
rect 6170 41168 6226 41224
rect 6294 41168 6350 41224
rect 6418 41168 6474 41224
rect 6542 41168 6598 41224
rect 6666 41168 6722 41224
rect 6790 41168 6846 41224
rect 6914 41168 6970 41224
rect 7038 41168 7094 41224
rect 5178 41044 5234 41100
rect 5302 41044 5358 41100
rect 5426 41044 5482 41100
rect 5550 41044 5606 41100
rect 5674 41044 5730 41100
rect 5798 41044 5854 41100
rect 5922 41044 5978 41100
rect 6046 41044 6102 41100
rect 6170 41044 6226 41100
rect 6294 41044 6350 41100
rect 6418 41044 6474 41100
rect 6542 41044 6598 41100
rect 6666 41044 6722 41100
rect 6790 41044 6846 41100
rect 6914 41044 6970 41100
rect 7038 41044 7094 41100
rect 5178 40920 5234 40976
rect 5302 40920 5358 40976
rect 5426 40920 5482 40976
rect 5550 40920 5606 40976
rect 5674 40920 5730 40976
rect 5798 40920 5854 40976
rect 5922 40920 5978 40976
rect 6046 40920 6102 40976
rect 6170 40920 6226 40976
rect 6294 40920 6350 40976
rect 6418 40920 6474 40976
rect 6542 40920 6598 40976
rect 6666 40920 6722 40976
rect 6790 40920 6846 40976
rect 6914 40920 6970 40976
rect 7038 40920 7094 40976
rect 5178 40796 5234 40852
rect 5302 40796 5358 40852
rect 5426 40796 5482 40852
rect 5550 40796 5606 40852
rect 5674 40796 5730 40852
rect 5798 40796 5854 40852
rect 5922 40796 5978 40852
rect 6046 40796 6102 40852
rect 6170 40796 6226 40852
rect 6294 40796 6350 40852
rect 6418 40796 6474 40852
rect 6542 40796 6598 40852
rect 6666 40796 6722 40852
rect 6790 40796 6846 40852
rect 6914 40796 6970 40852
rect 7038 40796 7094 40852
rect 5178 40672 5234 40728
rect 5302 40672 5358 40728
rect 5426 40672 5482 40728
rect 5550 40672 5606 40728
rect 5674 40672 5730 40728
rect 5798 40672 5854 40728
rect 5922 40672 5978 40728
rect 6046 40672 6102 40728
rect 6170 40672 6226 40728
rect 6294 40672 6350 40728
rect 6418 40672 6474 40728
rect 6542 40672 6598 40728
rect 6666 40672 6722 40728
rect 6790 40672 6846 40728
rect 6914 40672 6970 40728
rect 7038 40672 7094 40728
rect 5178 40548 5234 40604
rect 5302 40548 5358 40604
rect 5426 40548 5482 40604
rect 5550 40548 5606 40604
rect 5674 40548 5730 40604
rect 5798 40548 5854 40604
rect 5922 40548 5978 40604
rect 6046 40548 6102 40604
rect 6170 40548 6226 40604
rect 6294 40548 6350 40604
rect 6418 40548 6474 40604
rect 6542 40548 6598 40604
rect 6666 40548 6722 40604
rect 6790 40548 6846 40604
rect 6914 40548 6970 40604
rect 7038 40548 7094 40604
rect 5178 40424 5234 40480
rect 5302 40424 5358 40480
rect 5426 40424 5482 40480
rect 5550 40424 5606 40480
rect 5674 40424 5730 40480
rect 5798 40424 5854 40480
rect 5922 40424 5978 40480
rect 6046 40424 6102 40480
rect 6170 40424 6226 40480
rect 6294 40424 6350 40480
rect 6418 40424 6474 40480
rect 6542 40424 6598 40480
rect 6666 40424 6722 40480
rect 6790 40424 6846 40480
rect 6914 40424 6970 40480
rect 7038 40424 7094 40480
rect 5178 40300 5234 40356
rect 5302 40300 5358 40356
rect 5426 40300 5482 40356
rect 5550 40300 5606 40356
rect 5674 40300 5730 40356
rect 5798 40300 5854 40356
rect 5922 40300 5978 40356
rect 6046 40300 6102 40356
rect 6170 40300 6226 40356
rect 6294 40300 6350 40356
rect 6418 40300 6474 40356
rect 6542 40300 6598 40356
rect 6666 40300 6722 40356
rect 6790 40300 6846 40356
rect 6914 40300 6970 40356
rect 7038 40300 7094 40356
rect 5178 40176 5234 40232
rect 5302 40176 5358 40232
rect 5426 40176 5482 40232
rect 5550 40176 5606 40232
rect 5674 40176 5730 40232
rect 5798 40176 5854 40232
rect 5922 40176 5978 40232
rect 6046 40176 6102 40232
rect 6170 40176 6226 40232
rect 6294 40176 6350 40232
rect 6418 40176 6474 40232
rect 6542 40176 6598 40232
rect 6666 40176 6722 40232
rect 6790 40176 6846 40232
rect 6914 40176 6970 40232
rect 7038 40176 7094 40232
rect 5178 40052 5234 40108
rect 5302 40052 5358 40108
rect 5426 40052 5482 40108
rect 5550 40052 5606 40108
rect 5674 40052 5730 40108
rect 5798 40052 5854 40108
rect 5922 40052 5978 40108
rect 6046 40052 6102 40108
rect 6170 40052 6226 40108
rect 6294 40052 6350 40108
rect 6418 40052 6474 40108
rect 6542 40052 6598 40108
rect 6666 40052 6722 40108
rect 6790 40052 6846 40108
rect 6914 40052 6970 40108
rect 7038 40052 7094 40108
rect 7884 41292 7940 41348
rect 8008 41292 8064 41348
rect 8132 41292 8188 41348
rect 8256 41292 8312 41348
rect 8380 41292 8436 41348
rect 8504 41292 8560 41348
rect 8628 41292 8684 41348
rect 8752 41292 8808 41348
rect 8876 41292 8932 41348
rect 9000 41292 9056 41348
rect 9124 41292 9180 41348
rect 9248 41292 9304 41348
rect 9372 41292 9428 41348
rect 9496 41292 9552 41348
rect 9620 41292 9676 41348
rect 9744 41292 9800 41348
rect 7884 41168 7940 41224
rect 8008 41168 8064 41224
rect 8132 41168 8188 41224
rect 8256 41168 8312 41224
rect 8380 41168 8436 41224
rect 8504 41168 8560 41224
rect 8628 41168 8684 41224
rect 8752 41168 8808 41224
rect 8876 41168 8932 41224
rect 9000 41168 9056 41224
rect 9124 41168 9180 41224
rect 9248 41168 9304 41224
rect 9372 41168 9428 41224
rect 9496 41168 9552 41224
rect 9620 41168 9676 41224
rect 9744 41168 9800 41224
rect 7884 41044 7940 41100
rect 8008 41044 8064 41100
rect 8132 41044 8188 41100
rect 8256 41044 8312 41100
rect 8380 41044 8436 41100
rect 8504 41044 8560 41100
rect 8628 41044 8684 41100
rect 8752 41044 8808 41100
rect 8876 41044 8932 41100
rect 9000 41044 9056 41100
rect 9124 41044 9180 41100
rect 9248 41044 9304 41100
rect 9372 41044 9428 41100
rect 9496 41044 9552 41100
rect 9620 41044 9676 41100
rect 9744 41044 9800 41100
rect 7884 40920 7940 40976
rect 8008 40920 8064 40976
rect 8132 40920 8188 40976
rect 8256 40920 8312 40976
rect 8380 40920 8436 40976
rect 8504 40920 8560 40976
rect 8628 40920 8684 40976
rect 8752 40920 8808 40976
rect 8876 40920 8932 40976
rect 9000 40920 9056 40976
rect 9124 40920 9180 40976
rect 9248 40920 9304 40976
rect 9372 40920 9428 40976
rect 9496 40920 9552 40976
rect 9620 40920 9676 40976
rect 9744 40920 9800 40976
rect 7884 40796 7940 40852
rect 8008 40796 8064 40852
rect 8132 40796 8188 40852
rect 8256 40796 8312 40852
rect 8380 40796 8436 40852
rect 8504 40796 8560 40852
rect 8628 40796 8684 40852
rect 8752 40796 8808 40852
rect 8876 40796 8932 40852
rect 9000 40796 9056 40852
rect 9124 40796 9180 40852
rect 9248 40796 9304 40852
rect 9372 40796 9428 40852
rect 9496 40796 9552 40852
rect 9620 40796 9676 40852
rect 9744 40796 9800 40852
rect 7884 40672 7940 40728
rect 8008 40672 8064 40728
rect 8132 40672 8188 40728
rect 8256 40672 8312 40728
rect 8380 40672 8436 40728
rect 8504 40672 8560 40728
rect 8628 40672 8684 40728
rect 8752 40672 8808 40728
rect 8876 40672 8932 40728
rect 9000 40672 9056 40728
rect 9124 40672 9180 40728
rect 9248 40672 9304 40728
rect 9372 40672 9428 40728
rect 9496 40672 9552 40728
rect 9620 40672 9676 40728
rect 9744 40672 9800 40728
rect 7884 40548 7940 40604
rect 8008 40548 8064 40604
rect 8132 40548 8188 40604
rect 8256 40548 8312 40604
rect 8380 40548 8436 40604
rect 8504 40548 8560 40604
rect 8628 40548 8684 40604
rect 8752 40548 8808 40604
rect 8876 40548 8932 40604
rect 9000 40548 9056 40604
rect 9124 40548 9180 40604
rect 9248 40548 9304 40604
rect 9372 40548 9428 40604
rect 9496 40548 9552 40604
rect 9620 40548 9676 40604
rect 9744 40548 9800 40604
rect 7884 40424 7940 40480
rect 8008 40424 8064 40480
rect 8132 40424 8188 40480
rect 8256 40424 8312 40480
rect 8380 40424 8436 40480
rect 8504 40424 8560 40480
rect 8628 40424 8684 40480
rect 8752 40424 8808 40480
rect 8876 40424 8932 40480
rect 9000 40424 9056 40480
rect 9124 40424 9180 40480
rect 9248 40424 9304 40480
rect 9372 40424 9428 40480
rect 9496 40424 9552 40480
rect 9620 40424 9676 40480
rect 9744 40424 9800 40480
rect 7884 40300 7940 40356
rect 8008 40300 8064 40356
rect 8132 40300 8188 40356
rect 8256 40300 8312 40356
rect 8380 40300 8436 40356
rect 8504 40300 8560 40356
rect 8628 40300 8684 40356
rect 8752 40300 8808 40356
rect 8876 40300 8932 40356
rect 9000 40300 9056 40356
rect 9124 40300 9180 40356
rect 9248 40300 9304 40356
rect 9372 40300 9428 40356
rect 9496 40300 9552 40356
rect 9620 40300 9676 40356
rect 9744 40300 9800 40356
rect 7884 40176 7940 40232
rect 8008 40176 8064 40232
rect 8132 40176 8188 40232
rect 8256 40176 8312 40232
rect 8380 40176 8436 40232
rect 8504 40176 8560 40232
rect 8628 40176 8684 40232
rect 8752 40176 8808 40232
rect 8876 40176 8932 40232
rect 9000 40176 9056 40232
rect 9124 40176 9180 40232
rect 9248 40176 9304 40232
rect 9372 40176 9428 40232
rect 9496 40176 9552 40232
rect 9620 40176 9676 40232
rect 9744 40176 9800 40232
rect 7884 40052 7940 40108
rect 8008 40052 8064 40108
rect 8132 40052 8188 40108
rect 8256 40052 8312 40108
rect 8380 40052 8436 40108
rect 8504 40052 8560 40108
rect 8628 40052 8684 40108
rect 8752 40052 8808 40108
rect 8876 40052 8932 40108
rect 9000 40052 9056 40108
rect 9124 40052 9180 40108
rect 9248 40052 9304 40108
rect 9372 40052 9428 40108
rect 9496 40052 9552 40108
rect 9620 40052 9676 40108
rect 9744 40052 9800 40108
rect 10254 41292 10310 41348
rect 10378 41292 10434 41348
rect 10502 41292 10558 41348
rect 10626 41292 10682 41348
rect 10750 41292 10806 41348
rect 10874 41292 10930 41348
rect 10998 41292 11054 41348
rect 11122 41292 11178 41348
rect 11246 41292 11302 41348
rect 11370 41292 11426 41348
rect 11494 41292 11550 41348
rect 11618 41292 11674 41348
rect 11742 41292 11798 41348
rect 11866 41292 11922 41348
rect 11990 41292 12046 41348
rect 12114 41292 12170 41348
rect 10254 41168 10310 41224
rect 10378 41168 10434 41224
rect 10502 41168 10558 41224
rect 10626 41168 10682 41224
rect 10750 41168 10806 41224
rect 10874 41168 10930 41224
rect 10998 41168 11054 41224
rect 11122 41168 11178 41224
rect 11246 41168 11302 41224
rect 11370 41168 11426 41224
rect 11494 41168 11550 41224
rect 11618 41168 11674 41224
rect 11742 41168 11798 41224
rect 11866 41168 11922 41224
rect 11990 41168 12046 41224
rect 12114 41168 12170 41224
rect 10254 41044 10310 41100
rect 10378 41044 10434 41100
rect 10502 41044 10558 41100
rect 10626 41044 10682 41100
rect 10750 41044 10806 41100
rect 10874 41044 10930 41100
rect 10998 41044 11054 41100
rect 11122 41044 11178 41100
rect 11246 41044 11302 41100
rect 11370 41044 11426 41100
rect 11494 41044 11550 41100
rect 11618 41044 11674 41100
rect 11742 41044 11798 41100
rect 11866 41044 11922 41100
rect 11990 41044 12046 41100
rect 12114 41044 12170 41100
rect 10254 40920 10310 40976
rect 10378 40920 10434 40976
rect 10502 40920 10558 40976
rect 10626 40920 10682 40976
rect 10750 40920 10806 40976
rect 10874 40920 10930 40976
rect 10998 40920 11054 40976
rect 11122 40920 11178 40976
rect 11246 40920 11302 40976
rect 11370 40920 11426 40976
rect 11494 40920 11550 40976
rect 11618 40920 11674 40976
rect 11742 40920 11798 40976
rect 11866 40920 11922 40976
rect 11990 40920 12046 40976
rect 12114 40920 12170 40976
rect 10254 40796 10310 40852
rect 10378 40796 10434 40852
rect 10502 40796 10558 40852
rect 10626 40796 10682 40852
rect 10750 40796 10806 40852
rect 10874 40796 10930 40852
rect 10998 40796 11054 40852
rect 11122 40796 11178 40852
rect 11246 40796 11302 40852
rect 11370 40796 11426 40852
rect 11494 40796 11550 40852
rect 11618 40796 11674 40852
rect 11742 40796 11798 40852
rect 11866 40796 11922 40852
rect 11990 40796 12046 40852
rect 12114 40796 12170 40852
rect 10254 40672 10310 40728
rect 10378 40672 10434 40728
rect 10502 40672 10558 40728
rect 10626 40672 10682 40728
rect 10750 40672 10806 40728
rect 10874 40672 10930 40728
rect 10998 40672 11054 40728
rect 11122 40672 11178 40728
rect 11246 40672 11302 40728
rect 11370 40672 11426 40728
rect 11494 40672 11550 40728
rect 11618 40672 11674 40728
rect 11742 40672 11798 40728
rect 11866 40672 11922 40728
rect 11990 40672 12046 40728
rect 12114 40672 12170 40728
rect 10254 40548 10310 40604
rect 10378 40548 10434 40604
rect 10502 40548 10558 40604
rect 10626 40548 10682 40604
rect 10750 40548 10806 40604
rect 10874 40548 10930 40604
rect 10998 40548 11054 40604
rect 11122 40548 11178 40604
rect 11246 40548 11302 40604
rect 11370 40548 11426 40604
rect 11494 40548 11550 40604
rect 11618 40548 11674 40604
rect 11742 40548 11798 40604
rect 11866 40548 11922 40604
rect 11990 40548 12046 40604
rect 12114 40548 12170 40604
rect 10254 40424 10310 40480
rect 10378 40424 10434 40480
rect 10502 40424 10558 40480
rect 10626 40424 10682 40480
rect 10750 40424 10806 40480
rect 10874 40424 10930 40480
rect 10998 40424 11054 40480
rect 11122 40424 11178 40480
rect 11246 40424 11302 40480
rect 11370 40424 11426 40480
rect 11494 40424 11550 40480
rect 11618 40424 11674 40480
rect 11742 40424 11798 40480
rect 11866 40424 11922 40480
rect 11990 40424 12046 40480
rect 12114 40424 12170 40480
rect 10254 40300 10310 40356
rect 10378 40300 10434 40356
rect 10502 40300 10558 40356
rect 10626 40300 10682 40356
rect 10750 40300 10806 40356
rect 10874 40300 10930 40356
rect 10998 40300 11054 40356
rect 11122 40300 11178 40356
rect 11246 40300 11302 40356
rect 11370 40300 11426 40356
rect 11494 40300 11550 40356
rect 11618 40300 11674 40356
rect 11742 40300 11798 40356
rect 11866 40300 11922 40356
rect 11990 40300 12046 40356
rect 12114 40300 12170 40356
rect 10254 40176 10310 40232
rect 10378 40176 10434 40232
rect 10502 40176 10558 40232
rect 10626 40176 10682 40232
rect 10750 40176 10806 40232
rect 10874 40176 10930 40232
rect 10998 40176 11054 40232
rect 11122 40176 11178 40232
rect 11246 40176 11302 40232
rect 11370 40176 11426 40232
rect 11494 40176 11550 40232
rect 11618 40176 11674 40232
rect 11742 40176 11798 40232
rect 11866 40176 11922 40232
rect 11990 40176 12046 40232
rect 12114 40176 12170 40232
rect 10254 40052 10310 40108
rect 10378 40052 10434 40108
rect 10502 40052 10558 40108
rect 10626 40052 10682 40108
rect 10750 40052 10806 40108
rect 10874 40052 10930 40108
rect 10998 40052 11054 40108
rect 11122 40052 11178 40108
rect 11246 40052 11302 40108
rect 11370 40052 11426 40108
rect 11494 40052 11550 40108
rect 11618 40052 11674 40108
rect 11742 40052 11798 40108
rect 11866 40052 11922 40108
rect 11990 40052 12046 40108
rect 12114 40052 12170 40108
rect 12871 41292 12927 41348
rect 12995 41292 13051 41348
rect 13119 41292 13175 41348
rect 13243 41292 13299 41348
rect 13367 41292 13423 41348
rect 13491 41292 13547 41348
rect 13615 41292 13671 41348
rect 13739 41292 13795 41348
rect 13863 41292 13919 41348
rect 13987 41292 14043 41348
rect 14111 41292 14167 41348
rect 14235 41292 14291 41348
rect 14359 41292 14415 41348
rect 14483 41292 14539 41348
rect 14607 41292 14663 41348
rect 12871 41168 12927 41224
rect 12995 41168 13051 41224
rect 13119 41168 13175 41224
rect 13243 41168 13299 41224
rect 13367 41168 13423 41224
rect 13491 41168 13547 41224
rect 13615 41168 13671 41224
rect 13739 41168 13795 41224
rect 13863 41168 13919 41224
rect 13987 41168 14043 41224
rect 14111 41168 14167 41224
rect 14235 41168 14291 41224
rect 14359 41168 14415 41224
rect 14483 41168 14539 41224
rect 14607 41168 14663 41224
rect 12871 41044 12927 41100
rect 12995 41044 13051 41100
rect 13119 41044 13175 41100
rect 13243 41044 13299 41100
rect 13367 41044 13423 41100
rect 13491 41044 13547 41100
rect 13615 41044 13671 41100
rect 13739 41044 13795 41100
rect 13863 41044 13919 41100
rect 13987 41044 14043 41100
rect 14111 41044 14167 41100
rect 14235 41044 14291 41100
rect 14359 41044 14415 41100
rect 14483 41044 14539 41100
rect 14607 41044 14663 41100
rect 12871 40920 12927 40976
rect 12995 40920 13051 40976
rect 13119 40920 13175 40976
rect 13243 40920 13299 40976
rect 13367 40920 13423 40976
rect 13491 40920 13547 40976
rect 13615 40920 13671 40976
rect 13739 40920 13795 40976
rect 13863 40920 13919 40976
rect 13987 40920 14043 40976
rect 14111 40920 14167 40976
rect 14235 40920 14291 40976
rect 14359 40920 14415 40976
rect 14483 40920 14539 40976
rect 14607 40920 14663 40976
rect 12871 40796 12927 40852
rect 12995 40796 13051 40852
rect 13119 40796 13175 40852
rect 13243 40796 13299 40852
rect 13367 40796 13423 40852
rect 13491 40796 13547 40852
rect 13615 40796 13671 40852
rect 13739 40796 13795 40852
rect 13863 40796 13919 40852
rect 13987 40796 14043 40852
rect 14111 40796 14167 40852
rect 14235 40796 14291 40852
rect 14359 40796 14415 40852
rect 14483 40796 14539 40852
rect 14607 40796 14663 40852
rect 12871 40672 12927 40728
rect 12995 40672 13051 40728
rect 13119 40672 13175 40728
rect 13243 40672 13299 40728
rect 13367 40672 13423 40728
rect 13491 40672 13547 40728
rect 13615 40672 13671 40728
rect 13739 40672 13795 40728
rect 13863 40672 13919 40728
rect 13987 40672 14043 40728
rect 14111 40672 14167 40728
rect 14235 40672 14291 40728
rect 14359 40672 14415 40728
rect 14483 40672 14539 40728
rect 14607 40672 14663 40728
rect 12871 40548 12927 40604
rect 12995 40548 13051 40604
rect 13119 40548 13175 40604
rect 13243 40548 13299 40604
rect 13367 40548 13423 40604
rect 13491 40548 13547 40604
rect 13615 40548 13671 40604
rect 13739 40548 13795 40604
rect 13863 40548 13919 40604
rect 13987 40548 14043 40604
rect 14111 40548 14167 40604
rect 14235 40548 14291 40604
rect 14359 40548 14415 40604
rect 14483 40548 14539 40604
rect 14607 40548 14663 40604
rect 12871 40424 12927 40480
rect 12995 40424 13051 40480
rect 13119 40424 13175 40480
rect 13243 40424 13299 40480
rect 13367 40424 13423 40480
rect 13491 40424 13547 40480
rect 13615 40424 13671 40480
rect 13739 40424 13795 40480
rect 13863 40424 13919 40480
rect 13987 40424 14043 40480
rect 14111 40424 14167 40480
rect 14235 40424 14291 40480
rect 14359 40424 14415 40480
rect 14483 40424 14539 40480
rect 14607 40424 14663 40480
rect 12871 40300 12927 40356
rect 12995 40300 13051 40356
rect 13119 40300 13175 40356
rect 13243 40300 13299 40356
rect 13367 40300 13423 40356
rect 13491 40300 13547 40356
rect 13615 40300 13671 40356
rect 13739 40300 13795 40356
rect 13863 40300 13919 40356
rect 13987 40300 14043 40356
rect 14111 40300 14167 40356
rect 14235 40300 14291 40356
rect 14359 40300 14415 40356
rect 14483 40300 14539 40356
rect 14607 40300 14663 40356
rect 12871 40176 12927 40232
rect 12995 40176 13051 40232
rect 13119 40176 13175 40232
rect 13243 40176 13299 40232
rect 13367 40176 13423 40232
rect 13491 40176 13547 40232
rect 13615 40176 13671 40232
rect 13739 40176 13795 40232
rect 13863 40176 13919 40232
rect 13987 40176 14043 40232
rect 14111 40176 14167 40232
rect 14235 40176 14291 40232
rect 14359 40176 14415 40232
rect 14483 40176 14539 40232
rect 14607 40176 14663 40232
rect 12871 40052 12927 40108
rect 12995 40052 13051 40108
rect 13119 40052 13175 40108
rect 13243 40052 13299 40108
rect 13367 40052 13423 40108
rect 13491 40052 13547 40108
rect 13615 40052 13671 40108
rect 13739 40052 13795 40108
rect 13863 40052 13919 40108
rect 13987 40052 14043 40108
rect 14111 40052 14167 40108
rect 14235 40052 14291 40108
rect 14359 40052 14415 40108
rect 14483 40052 14539 40108
rect 14607 40052 14663 40108
rect 2808 39692 2864 39748
rect 2932 39692 2988 39748
rect 3056 39692 3112 39748
rect 3180 39692 3236 39748
rect 3304 39692 3360 39748
rect 3428 39692 3484 39748
rect 3552 39692 3608 39748
rect 3676 39692 3732 39748
rect 3800 39692 3856 39748
rect 3924 39692 3980 39748
rect 4048 39692 4104 39748
rect 4172 39692 4228 39748
rect 4296 39692 4352 39748
rect 4420 39692 4476 39748
rect 4544 39692 4600 39748
rect 4668 39692 4724 39748
rect 2808 39568 2864 39624
rect 2932 39568 2988 39624
rect 3056 39568 3112 39624
rect 3180 39568 3236 39624
rect 3304 39568 3360 39624
rect 3428 39568 3484 39624
rect 3552 39568 3608 39624
rect 3676 39568 3732 39624
rect 3800 39568 3856 39624
rect 3924 39568 3980 39624
rect 4048 39568 4104 39624
rect 4172 39568 4228 39624
rect 4296 39568 4352 39624
rect 4420 39568 4476 39624
rect 4544 39568 4600 39624
rect 4668 39568 4724 39624
rect 2808 39444 2864 39500
rect 2932 39444 2988 39500
rect 3056 39444 3112 39500
rect 3180 39444 3236 39500
rect 3304 39444 3360 39500
rect 3428 39444 3484 39500
rect 3552 39444 3608 39500
rect 3676 39444 3732 39500
rect 3800 39444 3856 39500
rect 3924 39444 3980 39500
rect 4048 39444 4104 39500
rect 4172 39444 4228 39500
rect 4296 39444 4352 39500
rect 4420 39444 4476 39500
rect 4544 39444 4600 39500
rect 4668 39444 4724 39500
rect 2808 39320 2864 39376
rect 2932 39320 2988 39376
rect 3056 39320 3112 39376
rect 3180 39320 3236 39376
rect 3304 39320 3360 39376
rect 3428 39320 3484 39376
rect 3552 39320 3608 39376
rect 3676 39320 3732 39376
rect 3800 39320 3856 39376
rect 3924 39320 3980 39376
rect 4048 39320 4104 39376
rect 4172 39320 4228 39376
rect 4296 39320 4352 39376
rect 4420 39320 4476 39376
rect 4544 39320 4600 39376
rect 4668 39320 4724 39376
rect 2808 39196 2864 39252
rect 2932 39196 2988 39252
rect 3056 39196 3112 39252
rect 3180 39196 3236 39252
rect 3304 39196 3360 39252
rect 3428 39196 3484 39252
rect 3552 39196 3608 39252
rect 3676 39196 3732 39252
rect 3800 39196 3856 39252
rect 3924 39196 3980 39252
rect 4048 39196 4104 39252
rect 4172 39196 4228 39252
rect 4296 39196 4352 39252
rect 4420 39196 4476 39252
rect 4544 39196 4600 39252
rect 4668 39196 4724 39252
rect 2808 39072 2864 39128
rect 2932 39072 2988 39128
rect 3056 39072 3112 39128
rect 3180 39072 3236 39128
rect 3304 39072 3360 39128
rect 3428 39072 3484 39128
rect 3552 39072 3608 39128
rect 3676 39072 3732 39128
rect 3800 39072 3856 39128
rect 3924 39072 3980 39128
rect 4048 39072 4104 39128
rect 4172 39072 4228 39128
rect 4296 39072 4352 39128
rect 4420 39072 4476 39128
rect 4544 39072 4600 39128
rect 4668 39072 4724 39128
rect 2808 38948 2864 39004
rect 2932 38948 2988 39004
rect 3056 38948 3112 39004
rect 3180 38948 3236 39004
rect 3304 38948 3360 39004
rect 3428 38948 3484 39004
rect 3552 38948 3608 39004
rect 3676 38948 3732 39004
rect 3800 38948 3856 39004
rect 3924 38948 3980 39004
rect 4048 38948 4104 39004
rect 4172 38948 4228 39004
rect 4296 38948 4352 39004
rect 4420 38948 4476 39004
rect 4544 38948 4600 39004
rect 4668 38948 4724 39004
rect 2808 38824 2864 38880
rect 2932 38824 2988 38880
rect 3056 38824 3112 38880
rect 3180 38824 3236 38880
rect 3304 38824 3360 38880
rect 3428 38824 3484 38880
rect 3552 38824 3608 38880
rect 3676 38824 3732 38880
rect 3800 38824 3856 38880
rect 3924 38824 3980 38880
rect 4048 38824 4104 38880
rect 4172 38824 4228 38880
rect 4296 38824 4352 38880
rect 4420 38824 4476 38880
rect 4544 38824 4600 38880
rect 4668 38824 4724 38880
rect 2808 38700 2864 38756
rect 2932 38700 2988 38756
rect 3056 38700 3112 38756
rect 3180 38700 3236 38756
rect 3304 38700 3360 38756
rect 3428 38700 3484 38756
rect 3552 38700 3608 38756
rect 3676 38700 3732 38756
rect 3800 38700 3856 38756
rect 3924 38700 3980 38756
rect 4048 38700 4104 38756
rect 4172 38700 4228 38756
rect 4296 38700 4352 38756
rect 4420 38700 4476 38756
rect 4544 38700 4600 38756
rect 4668 38700 4724 38756
rect 2808 38576 2864 38632
rect 2932 38576 2988 38632
rect 3056 38576 3112 38632
rect 3180 38576 3236 38632
rect 3304 38576 3360 38632
rect 3428 38576 3484 38632
rect 3552 38576 3608 38632
rect 3676 38576 3732 38632
rect 3800 38576 3856 38632
rect 3924 38576 3980 38632
rect 4048 38576 4104 38632
rect 4172 38576 4228 38632
rect 4296 38576 4352 38632
rect 4420 38576 4476 38632
rect 4544 38576 4600 38632
rect 4668 38576 4724 38632
rect 2808 38452 2864 38508
rect 2932 38452 2988 38508
rect 3056 38452 3112 38508
rect 3180 38452 3236 38508
rect 3304 38452 3360 38508
rect 3428 38452 3484 38508
rect 3552 38452 3608 38508
rect 3676 38452 3732 38508
rect 3800 38452 3856 38508
rect 3924 38452 3980 38508
rect 4048 38452 4104 38508
rect 4172 38452 4228 38508
rect 4296 38452 4352 38508
rect 4420 38452 4476 38508
rect 4544 38452 4600 38508
rect 4668 38452 4724 38508
rect 5178 39692 5234 39748
rect 5302 39692 5358 39748
rect 5426 39692 5482 39748
rect 5550 39692 5606 39748
rect 5674 39692 5730 39748
rect 5798 39692 5854 39748
rect 5922 39692 5978 39748
rect 6046 39692 6102 39748
rect 6170 39692 6226 39748
rect 6294 39692 6350 39748
rect 6418 39692 6474 39748
rect 6542 39692 6598 39748
rect 6666 39692 6722 39748
rect 6790 39692 6846 39748
rect 6914 39692 6970 39748
rect 7038 39692 7094 39748
rect 5178 39568 5234 39624
rect 5302 39568 5358 39624
rect 5426 39568 5482 39624
rect 5550 39568 5606 39624
rect 5674 39568 5730 39624
rect 5798 39568 5854 39624
rect 5922 39568 5978 39624
rect 6046 39568 6102 39624
rect 6170 39568 6226 39624
rect 6294 39568 6350 39624
rect 6418 39568 6474 39624
rect 6542 39568 6598 39624
rect 6666 39568 6722 39624
rect 6790 39568 6846 39624
rect 6914 39568 6970 39624
rect 7038 39568 7094 39624
rect 5178 39444 5234 39500
rect 5302 39444 5358 39500
rect 5426 39444 5482 39500
rect 5550 39444 5606 39500
rect 5674 39444 5730 39500
rect 5798 39444 5854 39500
rect 5922 39444 5978 39500
rect 6046 39444 6102 39500
rect 6170 39444 6226 39500
rect 6294 39444 6350 39500
rect 6418 39444 6474 39500
rect 6542 39444 6598 39500
rect 6666 39444 6722 39500
rect 6790 39444 6846 39500
rect 6914 39444 6970 39500
rect 7038 39444 7094 39500
rect 5178 39320 5234 39376
rect 5302 39320 5358 39376
rect 5426 39320 5482 39376
rect 5550 39320 5606 39376
rect 5674 39320 5730 39376
rect 5798 39320 5854 39376
rect 5922 39320 5978 39376
rect 6046 39320 6102 39376
rect 6170 39320 6226 39376
rect 6294 39320 6350 39376
rect 6418 39320 6474 39376
rect 6542 39320 6598 39376
rect 6666 39320 6722 39376
rect 6790 39320 6846 39376
rect 6914 39320 6970 39376
rect 7038 39320 7094 39376
rect 5178 39196 5234 39252
rect 5302 39196 5358 39252
rect 5426 39196 5482 39252
rect 5550 39196 5606 39252
rect 5674 39196 5730 39252
rect 5798 39196 5854 39252
rect 5922 39196 5978 39252
rect 6046 39196 6102 39252
rect 6170 39196 6226 39252
rect 6294 39196 6350 39252
rect 6418 39196 6474 39252
rect 6542 39196 6598 39252
rect 6666 39196 6722 39252
rect 6790 39196 6846 39252
rect 6914 39196 6970 39252
rect 7038 39196 7094 39252
rect 5178 39072 5234 39128
rect 5302 39072 5358 39128
rect 5426 39072 5482 39128
rect 5550 39072 5606 39128
rect 5674 39072 5730 39128
rect 5798 39072 5854 39128
rect 5922 39072 5978 39128
rect 6046 39072 6102 39128
rect 6170 39072 6226 39128
rect 6294 39072 6350 39128
rect 6418 39072 6474 39128
rect 6542 39072 6598 39128
rect 6666 39072 6722 39128
rect 6790 39072 6846 39128
rect 6914 39072 6970 39128
rect 7038 39072 7094 39128
rect 5178 38948 5234 39004
rect 5302 38948 5358 39004
rect 5426 38948 5482 39004
rect 5550 38948 5606 39004
rect 5674 38948 5730 39004
rect 5798 38948 5854 39004
rect 5922 38948 5978 39004
rect 6046 38948 6102 39004
rect 6170 38948 6226 39004
rect 6294 38948 6350 39004
rect 6418 38948 6474 39004
rect 6542 38948 6598 39004
rect 6666 38948 6722 39004
rect 6790 38948 6846 39004
rect 6914 38948 6970 39004
rect 7038 38948 7094 39004
rect 5178 38824 5234 38880
rect 5302 38824 5358 38880
rect 5426 38824 5482 38880
rect 5550 38824 5606 38880
rect 5674 38824 5730 38880
rect 5798 38824 5854 38880
rect 5922 38824 5978 38880
rect 6046 38824 6102 38880
rect 6170 38824 6226 38880
rect 6294 38824 6350 38880
rect 6418 38824 6474 38880
rect 6542 38824 6598 38880
rect 6666 38824 6722 38880
rect 6790 38824 6846 38880
rect 6914 38824 6970 38880
rect 7038 38824 7094 38880
rect 5178 38700 5234 38756
rect 5302 38700 5358 38756
rect 5426 38700 5482 38756
rect 5550 38700 5606 38756
rect 5674 38700 5730 38756
rect 5798 38700 5854 38756
rect 5922 38700 5978 38756
rect 6046 38700 6102 38756
rect 6170 38700 6226 38756
rect 6294 38700 6350 38756
rect 6418 38700 6474 38756
rect 6542 38700 6598 38756
rect 6666 38700 6722 38756
rect 6790 38700 6846 38756
rect 6914 38700 6970 38756
rect 7038 38700 7094 38756
rect 5178 38576 5234 38632
rect 5302 38576 5358 38632
rect 5426 38576 5482 38632
rect 5550 38576 5606 38632
rect 5674 38576 5730 38632
rect 5798 38576 5854 38632
rect 5922 38576 5978 38632
rect 6046 38576 6102 38632
rect 6170 38576 6226 38632
rect 6294 38576 6350 38632
rect 6418 38576 6474 38632
rect 6542 38576 6598 38632
rect 6666 38576 6722 38632
rect 6790 38576 6846 38632
rect 6914 38576 6970 38632
rect 7038 38576 7094 38632
rect 5178 38452 5234 38508
rect 5302 38452 5358 38508
rect 5426 38452 5482 38508
rect 5550 38452 5606 38508
rect 5674 38452 5730 38508
rect 5798 38452 5854 38508
rect 5922 38452 5978 38508
rect 6046 38452 6102 38508
rect 6170 38452 6226 38508
rect 6294 38452 6350 38508
rect 6418 38452 6474 38508
rect 6542 38452 6598 38508
rect 6666 38452 6722 38508
rect 6790 38452 6846 38508
rect 6914 38452 6970 38508
rect 7038 38452 7094 38508
rect 7884 39692 7940 39748
rect 8008 39692 8064 39748
rect 8132 39692 8188 39748
rect 8256 39692 8312 39748
rect 8380 39692 8436 39748
rect 8504 39692 8560 39748
rect 8628 39692 8684 39748
rect 8752 39692 8808 39748
rect 8876 39692 8932 39748
rect 9000 39692 9056 39748
rect 9124 39692 9180 39748
rect 9248 39692 9304 39748
rect 9372 39692 9428 39748
rect 9496 39692 9552 39748
rect 9620 39692 9676 39748
rect 9744 39692 9800 39748
rect 7884 39568 7940 39624
rect 8008 39568 8064 39624
rect 8132 39568 8188 39624
rect 8256 39568 8312 39624
rect 8380 39568 8436 39624
rect 8504 39568 8560 39624
rect 8628 39568 8684 39624
rect 8752 39568 8808 39624
rect 8876 39568 8932 39624
rect 9000 39568 9056 39624
rect 9124 39568 9180 39624
rect 9248 39568 9304 39624
rect 9372 39568 9428 39624
rect 9496 39568 9552 39624
rect 9620 39568 9676 39624
rect 9744 39568 9800 39624
rect 7884 39444 7940 39500
rect 8008 39444 8064 39500
rect 8132 39444 8188 39500
rect 8256 39444 8312 39500
rect 8380 39444 8436 39500
rect 8504 39444 8560 39500
rect 8628 39444 8684 39500
rect 8752 39444 8808 39500
rect 8876 39444 8932 39500
rect 9000 39444 9056 39500
rect 9124 39444 9180 39500
rect 9248 39444 9304 39500
rect 9372 39444 9428 39500
rect 9496 39444 9552 39500
rect 9620 39444 9676 39500
rect 9744 39444 9800 39500
rect 7884 39320 7940 39376
rect 8008 39320 8064 39376
rect 8132 39320 8188 39376
rect 8256 39320 8312 39376
rect 8380 39320 8436 39376
rect 8504 39320 8560 39376
rect 8628 39320 8684 39376
rect 8752 39320 8808 39376
rect 8876 39320 8932 39376
rect 9000 39320 9056 39376
rect 9124 39320 9180 39376
rect 9248 39320 9304 39376
rect 9372 39320 9428 39376
rect 9496 39320 9552 39376
rect 9620 39320 9676 39376
rect 9744 39320 9800 39376
rect 7884 39196 7940 39252
rect 8008 39196 8064 39252
rect 8132 39196 8188 39252
rect 8256 39196 8312 39252
rect 8380 39196 8436 39252
rect 8504 39196 8560 39252
rect 8628 39196 8684 39252
rect 8752 39196 8808 39252
rect 8876 39196 8932 39252
rect 9000 39196 9056 39252
rect 9124 39196 9180 39252
rect 9248 39196 9304 39252
rect 9372 39196 9428 39252
rect 9496 39196 9552 39252
rect 9620 39196 9676 39252
rect 9744 39196 9800 39252
rect 7884 39072 7940 39128
rect 8008 39072 8064 39128
rect 8132 39072 8188 39128
rect 8256 39072 8312 39128
rect 8380 39072 8436 39128
rect 8504 39072 8560 39128
rect 8628 39072 8684 39128
rect 8752 39072 8808 39128
rect 8876 39072 8932 39128
rect 9000 39072 9056 39128
rect 9124 39072 9180 39128
rect 9248 39072 9304 39128
rect 9372 39072 9428 39128
rect 9496 39072 9552 39128
rect 9620 39072 9676 39128
rect 9744 39072 9800 39128
rect 7884 38948 7940 39004
rect 8008 38948 8064 39004
rect 8132 38948 8188 39004
rect 8256 38948 8312 39004
rect 8380 38948 8436 39004
rect 8504 38948 8560 39004
rect 8628 38948 8684 39004
rect 8752 38948 8808 39004
rect 8876 38948 8932 39004
rect 9000 38948 9056 39004
rect 9124 38948 9180 39004
rect 9248 38948 9304 39004
rect 9372 38948 9428 39004
rect 9496 38948 9552 39004
rect 9620 38948 9676 39004
rect 9744 38948 9800 39004
rect 7884 38824 7940 38880
rect 8008 38824 8064 38880
rect 8132 38824 8188 38880
rect 8256 38824 8312 38880
rect 8380 38824 8436 38880
rect 8504 38824 8560 38880
rect 8628 38824 8684 38880
rect 8752 38824 8808 38880
rect 8876 38824 8932 38880
rect 9000 38824 9056 38880
rect 9124 38824 9180 38880
rect 9248 38824 9304 38880
rect 9372 38824 9428 38880
rect 9496 38824 9552 38880
rect 9620 38824 9676 38880
rect 9744 38824 9800 38880
rect 7884 38700 7940 38756
rect 8008 38700 8064 38756
rect 8132 38700 8188 38756
rect 8256 38700 8312 38756
rect 8380 38700 8436 38756
rect 8504 38700 8560 38756
rect 8628 38700 8684 38756
rect 8752 38700 8808 38756
rect 8876 38700 8932 38756
rect 9000 38700 9056 38756
rect 9124 38700 9180 38756
rect 9248 38700 9304 38756
rect 9372 38700 9428 38756
rect 9496 38700 9552 38756
rect 9620 38700 9676 38756
rect 9744 38700 9800 38756
rect 7884 38576 7940 38632
rect 8008 38576 8064 38632
rect 8132 38576 8188 38632
rect 8256 38576 8312 38632
rect 8380 38576 8436 38632
rect 8504 38576 8560 38632
rect 8628 38576 8684 38632
rect 8752 38576 8808 38632
rect 8876 38576 8932 38632
rect 9000 38576 9056 38632
rect 9124 38576 9180 38632
rect 9248 38576 9304 38632
rect 9372 38576 9428 38632
rect 9496 38576 9552 38632
rect 9620 38576 9676 38632
rect 9744 38576 9800 38632
rect 7884 38452 7940 38508
rect 8008 38452 8064 38508
rect 8132 38452 8188 38508
rect 8256 38452 8312 38508
rect 8380 38452 8436 38508
rect 8504 38452 8560 38508
rect 8628 38452 8684 38508
rect 8752 38452 8808 38508
rect 8876 38452 8932 38508
rect 9000 38452 9056 38508
rect 9124 38452 9180 38508
rect 9248 38452 9304 38508
rect 9372 38452 9428 38508
rect 9496 38452 9552 38508
rect 9620 38452 9676 38508
rect 9744 38452 9800 38508
rect 10254 39692 10310 39748
rect 10378 39692 10434 39748
rect 10502 39692 10558 39748
rect 10626 39692 10682 39748
rect 10750 39692 10806 39748
rect 10874 39692 10930 39748
rect 10998 39692 11054 39748
rect 11122 39692 11178 39748
rect 11246 39692 11302 39748
rect 11370 39692 11426 39748
rect 11494 39692 11550 39748
rect 11618 39692 11674 39748
rect 11742 39692 11798 39748
rect 11866 39692 11922 39748
rect 11990 39692 12046 39748
rect 12114 39692 12170 39748
rect 10254 39568 10310 39624
rect 10378 39568 10434 39624
rect 10502 39568 10558 39624
rect 10626 39568 10682 39624
rect 10750 39568 10806 39624
rect 10874 39568 10930 39624
rect 10998 39568 11054 39624
rect 11122 39568 11178 39624
rect 11246 39568 11302 39624
rect 11370 39568 11426 39624
rect 11494 39568 11550 39624
rect 11618 39568 11674 39624
rect 11742 39568 11798 39624
rect 11866 39568 11922 39624
rect 11990 39568 12046 39624
rect 12114 39568 12170 39624
rect 10254 39444 10310 39500
rect 10378 39444 10434 39500
rect 10502 39444 10558 39500
rect 10626 39444 10682 39500
rect 10750 39444 10806 39500
rect 10874 39444 10930 39500
rect 10998 39444 11054 39500
rect 11122 39444 11178 39500
rect 11246 39444 11302 39500
rect 11370 39444 11426 39500
rect 11494 39444 11550 39500
rect 11618 39444 11674 39500
rect 11742 39444 11798 39500
rect 11866 39444 11922 39500
rect 11990 39444 12046 39500
rect 12114 39444 12170 39500
rect 10254 39320 10310 39376
rect 10378 39320 10434 39376
rect 10502 39320 10558 39376
rect 10626 39320 10682 39376
rect 10750 39320 10806 39376
rect 10874 39320 10930 39376
rect 10998 39320 11054 39376
rect 11122 39320 11178 39376
rect 11246 39320 11302 39376
rect 11370 39320 11426 39376
rect 11494 39320 11550 39376
rect 11618 39320 11674 39376
rect 11742 39320 11798 39376
rect 11866 39320 11922 39376
rect 11990 39320 12046 39376
rect 12114 39320 12170 39376
rect 10254 39196 10310 39252
rect 10378 39196 10434 39252
rect 10502 39196 10558 39252
rect 10626 39196 10682 39252
rect 10750 39196 10806 39252
rect 10874 39196 10930 39252
rect 10998 39196 11054 39252
rect 11122 39196 11178 39252
rect 11246 39196 11302 39252
rect 11370 39196 11426 39252
rect 11494 39196 11550 39252
rect 11618 39196 11674 39252
rect 11742 39196 11798 39252
rect 11866 39196 11922 39252
rect 11990 39196 12046 39252
rect 12114 39196 12170 39252
rect 10254 39072 10310 39128
rect 10378 39072 10434 39128
rect 10502 39072 10558 39128
rect 10626 39072 10682 39128
rect 10750 39072 10806 39128
rect 10874 39072 10930 39128
rect 10998 39072 11054 39128
rect 11122 39072 11178 39128
rect 11246 39072 11302 39128
rect 11370 39072 11426 39128
rect 11494 39072 11550 39128
rect 11618 39072 11674 39128
rect 11742 39072 11798 39128
rect 11866 39072 11922 39128
rect 11990 39072 12046 39128
rect 12114 39072 12170 39128
rect 10254 38948 10310 39004
rect 10378 38948 10434 39004
rect 10502 38948 10558 39004
rect 10626 38948 10682 39004
rect 10750 38948 10806 39004
rect 10874 38948 10930 39004
rect 10998 38948 11054 39004
rect 11122 38948 11178 39004
rect 11246 38948 11302 39004
rect 11370 38948 11426 39004
rect 11494 38948 11550 39004
rect 11618 38948 11674 39004
rect 11742 38948 11798 39004
rect 11866 38948 11922 39004
rect 11990 38948 12046 39004
rect 12114 38948 12170 39004
rect 10254 38824 10310 38880
rect 10378 38824 10434 38880
rect 10502 38824 10558 38880
rect 10626 38824 10682 38880
rect 10750 38824 10806 38880
rect 10874 38824 10930 38880
rect 10998 38824 11054 38880
rect 11122 38824 11178 38880
rect 11246 38824 11302 38880
rect 11370 38824 11426 38880
rect 11494 38824 11550 38880
rect 11618 38824 11674 38880
rect 11742 38824 11798 38880
rect 11866 38824 11922 38880
rect 11990 38824 12046 38880
rect 12114 38824 12170 38880
rect 10254 38700 10310 38756
rect 10378 38700 10434 38756
rect 10502 38700 10558 38756
rect 10626 38700 10682 38756
rect 10750 38700 10806 38756
rect 10874 38700 10930 38756
rect 10998 38700 11054 38756
rect 11122 38700 11178 38756
rect 11246 38700 11302 38756
rect 11370 38700 11426 38756
rect 11494 38700 11550 38756
rect 11618 38700 11674 38756
rect 11742 38700 11798 38756
rect 11866 38700 11922 38756
rect 11990 38700 12046 38756
rect 12114 38700 12170 38756
rect 10254 38576 10310 38632
rect 10378 38576 10434 38632
rect 10502 38576 10558 38632
rect 10626 38576 10682 38632
rect 10750 38576 10806 38632
rect 10874 38576 10930 38632
rect 10998 38576 11054 38632
rect 11122 38576 11178 38632
rect 11246 38576 11302 38632
rect 11370 38576 11426 38632
rect 11494 38576 11550 38632
rect 11618 38576 11674 38632
rect 11742 38576 11798 38632
rect 11866 38576 11922 38632
rect 11990 38576 12046 38632
rect 12114 38576 12170 38632
rect 10254 38452 10310 38508
rect 10378 38452 10434 38508
rect 10502 38452 10558 38508
rect 10626 38452 10682 38508
rect 10750 38452 10806 38508
rect 10874 38452 10930 38508
rect 10998 38452 11054 38508
rect 11122 38452 11178 38508
rect 11246 38452 11302 38508
rect 11370 38452 11426 38508
rect 11494 38452 11550 38508
rect 11618 38452 11674 38508
rect 11742 38452 11798 38508
rect 11866 38452 11922 38508
rect 11990 38452 12046 38508
rect 12114 38452 12170 38508
rect 12871 39692 12927 39748
rect 12995 39692 13051 39748
rect 13119 39692 13175 39748
rect 13243 39692 13299 39748
rect 13367 39692 13423 39748
rect 13491 39692 13547 39748
rect 13615 39692 13671 39748
rect 13739 39692 13795 39748
rect 13863 39692 13919 39748
rect 13987 39692 14043 39748
rect 14111 39692 14167 39748
rect 14235 39692 14291 39748
rect 14359 39692 14415 39748
rect 14483 39692 14539 39748
rect 14607 39692 14663 39748
rect 12871 39568 12927 39624
rect 12995 39568 13051 39624
rect 13119 39568 13175 39624
rect 13243 39568 13299 39624
rect 13367 39568 13423 39624
rect 13491 39568 13547 39624
rect 13615 39568 13671 39624
rect 13739 39568 13795 39624
rect 13863 39568 13919 39624
rect 13987 39568 14043 39624
rect 14111 39568 14167 39624
rect 14235 39568 14291 39624
rect 14359 39568 14415 39624
rect 14483 39568 14539 39624
rect 14607 39568 14663 39624
rect 12871 39444 12927 39500
rect 12995 39444 13051 39500
rect 13119 39444 13175 39500
rect 13243 39444 13299 39500
rect 13367 39444 13423 39500
rect 13491 39444 13547 39500
rect 13615 39444 13671 39500
rect 13739 39444 13795 39500
rect 13863 39444 13919 39500
rect 13987 39444 14043 39500
rect 14111 39444 14167 39500
rect 14235 39444 14291 39500
rect 14359 39444 14415 39500
rect 14483 39444 14539 39500
rect 14607 39444 14663 39500
rect 12871 39320 12927 39376
rect 12995 39320 13051 39376
rect 13119 39320 13175 39376
rect 13243 39320 13299 39376
rect 13367 39320 13423 39376
rect 13491 39320 13547 39376
rect 13615 39320 13671 39376
rect 13739 39320 13795 39376
rect 13863 39320 13919 39376
rect 13987 39320 14043 39376
rect 14111 39320 14167 39376
rect 14235 39320 14291 39376
rect 14359 39320 14415 39376
rect 14483 39320 14539 39376
rect 14607 39320 14663 39376
rect 12871 39196 12927 39252
rect 12995 39196 13051 39252
rect 13119 39196 13175 39252
rect 13243 39196 13299 39252
rect 13367 39196 13423 39252
rect 13491 39196 13547 39252
rect 13615 39196 13671 39252
rect 13739 39196 13795 39252
rect 13863 39196 13919 39252
rect 13987 39196 14043 39252
rect 14111 39196 14167 39252
rect 14235 39196 14291 39252
rect 14359 39196 14415 39252
rect 14483 39196 14539 39252
rect 14607 39196 14663 39252
rect 12871 39072 12927 39128
rect 12995 39072 13051 39128
rect 13119 39072 13175 39128
rect 13243 39072 13299 39128
rect 13367 39072 13423 39128
rect 13491 39072 13547 39128
rect 13615 39072 13671 39128
rect 13739 39072 13795 39128
rect 13863 39072 13919 39128
rect 13987 39072 14043 39128
rect 14111 39072 14167 39128
rect 14235 39072 14291 39128
rect 14359 39072 14415 39128
rect 14483 39072 14539 39128
rect 14607 39072 14663 39128
rect 12871 38948 12927 39004
rect 12995 38948 13051 39004
rect 13119 38948 13175 39004
rect 13243 38948 13299 39004
rect 13367 38948 13423 39004
rect 13491 38948 13547 39004
rect 13615 38948 13671 39004
rect 13739 38948 13795 39004
rect 13863 38948 13919 39004
rect 13987 38948 14043 39004
rect 14111 38948 14167 39004
rect 14235 38948 14291 39004
rect 14359 38948 14415 39004
rect 14483 38948 14539 39004
rect 14607 38948 14663 39004
rect 12871 38824 12927 38880
rect 12995 38824 13051 38880
rect 13119 38824 13175 38880
rect 13243 38824 13299 38880
rect 13367 38824 13423 38880
rect 13491 38824 13547 38880
rect 13615 38824 13671 38880
rect 13739 38824 13795 38880
rect 13863 38824 13919 38880
rect 13987 38824 14043 38880
rect 14111 38824 14167 38880
rect 14235 38824 14291 38880
rect 14359 38824 14415 38880
rect 14483 38824 14539 38880
rect 14607 38824 14663 38880
rect 12871 38700 12927 38756
rect 12995 38700 13051 38756
rect 13119 38700 13175 38756
rect 13243 38700 13299 38756
rect 13367 38700 13423 38756
rect 13491 38700 13547 38756
rect 13615 38700 13671 38756
rect 13739 38700 13795 38756
rect 13863 38700 13919 38756
rect 13987 38700 14043 38756
rect 14111 38700 14167 38756
rect 14235 38700 14291 38756
rect 14359 38700 14415 38756
rect 14483 38700 14539 38756
rect 14607 38700 14663 38756
rect 12871 38576 12927 38632
rect 12995 38576 13051 38632
rect 13119 38576 13175 38632
rect 13243 38576 13299 38632
rect 13367 38576 13423 38632
rect 13491 38576 13547 38632
rect 13615 38576 13671 38632
rect 13739 38576 13795 38632
rect 13863 38576 13919 38632
rect 13987 38576 14043 38632
rect 14111 38576 14167 38632
rect 14235 38576 14291 38632
rect 14359 38576 14415 38632
rect 14483 38576 14539 38632
rect 14607 38576 14663 38632
rect 12871 38452 12927 38508
rect 12995 38452 13051 38508
rect 13119 38452 13175 38508
rect 13243 38452 13299 38508
rect 13367 38452 13423 38508
rect 13491 38452 13547 38508
rect 13615 38452 13671 38508
rect 13739 38452 13795 38508
rect 13863 38452 13919 38508
rect 13987 38452 14043 38508
rect 14111 38452 14167 38508
rect 14235 38452 14291 38508
rect 14359 38452 14415 38508
rect 14483 38452 14539 38508
rect 14607 38452 14663 38508
rect 2289 38079 2345 38135
rect 2289 37947 2345 38003
rect 2289 37815 2345 37871
rect 2289 37683 2345 37739
rect 2289 37551 2345 37607
rect 2289 37419 2345 37475
rect 2289 37287 2345 37343
rect 2289 37155 2345 37211
rect 2289 37023 2345 37079
rect 2289 36891 2345 36947
rect 14902 38174 14958 38176
rect 14902 38122 14904 38174
rect 14904 38122 14956 38174
rect 14956 38122 14958 38174
rect 14902 38066 14958 38122
rect 14902 38014 14904 38066
rect 14904 38014 14956 38066
rect 14956 38014 14958 38066
rect 14902 37958 14958 38014
rect 14902 37906 14904 37958
rect 14904 37906 14956 37958
rect 14956 37906 14958 37958
rect 14902 37850 14958 37906
rect 14902 37798 14904 37850
rect 14904 37798 14956 37850
rect 14956 37798 14958 37850
rect 14902 37742 14958 37798
rect 14902 37690 14904 37742
rect 14904 37690 14956 37742
rect 14956 37690 14958 37742
rect 14902 37634 14958 37690
rect 14902 37582 14904 37634
rect 14904 37582 14956 37634
rect 14956 37582 14958 37634
rect 14902 37526 14958 37582
rect 14902 37474 14904 37526
rect 14904 37474 14956 37526
rect 14956 37474 14958 37526
rect 14902 37418 14958 37474
rect 14902 37366 14904 37418
rect 14904 37366 14956 37418
rect 14956 37366 14958 37418
rect 14902 37310 14958 37366
rect 14902 37258 14904 37310
rect 14904 37258 14956 37310
rect 14956 37258 14958 37310
rect 14902 37202 14958 37258
rect 14902 37150 14904 37202
rect 14904 37150 14956 37202
rect 14956 37150 14958 37202
rect 14902 37094 14958 37150
rect 14902 37042 14904 37094
rect 14904 37042 14956 37094
rect 14956 37042 14958 37094
rect 14902 36986 14958 37042
rect 14902 36934 14904 36986
rect 14904 36934 14956 36986
rect 14956 36934 14958 36986
rect 14902 36878 14958 36934
rect 14902 36826 14904 36878
rect 14904 36826 14956 36878
rect 14956 36826 14958 36878
rect 14902 36824 14958 36826
rect 2491 36498 2547 36554
rect 2615 36498 2671 36554
rect 2491 36374 2547 36430
rect 2615 36374 2671 36430
rect 2491 36250 2547 36306
rect 2615 36250 2671 36306
rect 2491 36126 2547 36182
rect 2615 36126 2671 36182
rect 2491 36002 2547 36058
rect 2615 36002 2671 36058
rect 2491 35878 2547 35934
rect 2615 35878 2671 35934
rect 2491 35754 2547 35810
rect 2615 35754 2671 35810
rect 2491 35630 2547 35686
rect 2615 35630 2671 35686
rect 2491 35506 2547 35562
rect 2615 35506 2671 35562
rect 2491 35382 2547 35438
rect 2615 35382 2671 35438
rect 2491 35258 2547 35314
rect 2615 35258 2671 35314
rect 2491 35134 2547 35190
rect 2615 35134 2671 35190
rect 2491 35010 2547 35066
rect 2615 35010 2671 35066
rect 2491 34886 2547 34942
rect 2615 34886 2671 34942
rect 2491 34762 2547 34818
rect 2615 34762 2671 34818
rect 2491 34638 2547 34694
rect 2615 34638 2671 34694
rect 2491 34514 2547 34570
rect 2615 34514 2671 34570
rect 2491 34390 2547 34446
rect 2615 34390 2671 34446
rect 2491 34266 2547 34322
rect 2615 34266 2671 34322
rect 2491 34142 2547 34198
rect 2615 34142 2671 34198
rect 2491 34018 2547 34074
rect 2615 34018 2671 34074
rect 2491 33894 2547 33950
rect 2615 33894 2671 33950
rect 2491 33770 2547 33826
rect 2615 33770 2671 33826
rect 2491 33646 2547 33702
rect 2615 33646 2671 33702
rect 4861 36498 4917 36554
rect 4985 36498 5041 36554
rect 4861 36374 4917 36430
rect 4985 36374 5041 36430
rect 4861 36250 4917 36306
rect 4985 36250 5041 36306
rect 4861 36126 4917 36182
rect 4985 36126 5041 36182
rect 4861 36002 4917 36058
rect 4985 36002 5041 36058
rect 4861 35878 4917 35934
rect 4985 35878 5041 35934
rect 4861 35754 4917 35810
rect 4985 35754 5041 35810
rect 4861 35630 4917 35686
rect 4985 35630 5041 35686
rect 4861 35506 4917 35562
rect 4985 35506 5041 35562
rect 4861 35382 4917 35438
rect 4985 35382 5041 35438
rect 4861 35258 4917 35314
rect 4985 35258 5041 35314
rect 4861 35134 4917 35190
rect 4985 35134 5041 35190
rect 4861 35010 4917 35066
rect 4985 35010 5041 35066
rect 4861 34886 4917 34942
rect 4985 34886 5041 34942
rect 4861 34762 4917 34818
rect 4985 34762 5041 34818
rect 4861 34638 4917 34694
rect 4985 34638 5041 34694
rect 4861 34514 4917 34570
rect 4985 34514 5041 34570
rect 4861 34390 4917 34446
rect 4985 34390 5041 34446
rect 4861 34266 4917 34322
rect 4985 34266 5041 34322
rect 4861 34142 4917 34198
rect 4985 34142 5041 34198
rect 4861 34018 4917 34074
rect 4985 34018 5041 34074
rect 4861 33894 4917 33950
rect 4985 33894 5041 33950
rect 4861 33770 4917 33826
rect 4985 33770 5041 33826
rect 4861 33646 4917 33702
rect 4985 33646 5041 33702
rect 7275 36498 7331 36554
rect 7399 36498 7455 36554
rect 7523 36498 7579 36554
rect 7647 36498 7703 36554
rect 7275 36374 7331 36430
rect 7399 36374 7455 36430
rect 7523 36374 7579 36430
rect 7647 36374 7703 36430
rect 7275 36250 7331 36306
rect 7399 36250 7455 36306
rect 7523 36250 7579 36306
rect 7647 36250 7703 36306
rect 7275 36126 7331 36182
rect 7399 36126 7455 36182
rect 7523 36126 7579 36182
rect 7647 36126 7703 36182
rect 7275 36002 7331 36058
rect 7399 36002 7455 36058
rect 7523 36002 7579 36058
rect 7647 36002 7703 36058
rect 7275 35878 7331 35934
rect 7399 35878 7455 35934
rect 7523 35878 7579 35934
rect 7647 35878 7703 35934
rect 7275 35754 7331 35810
rect 7399 35754 7455 35810
rect 7523 35754 7579 35810
rect 7647 35754 7703 35810
rect 7275 35630 7331 35686
rect 7399 35630 7455 35686
rect 7523 35630 7579 35686
rect 7647 35630 7703 35686
rect 7275 35506 7331 35562
rect 7399 35506 7455 35562
rect 7523 35506 7579 35562
rect 7647 35506 7703 35562
rect 7275 35382 7331 35438
rect 7399 35382 7455 35438
rect 7523 35382 7579 35438
rect 7647 35382 7703 35438
rect 7275 35258 7331 35314
rect 7399 35258 7455 35314
rect 7523 35258 7579 35314
rect 7647 35258 7703 35314
rect 7275 35134 7331 35190
rect 7399 35134 7455 35190
rect 7523 35134 7579 35190
rect 7647 35134 7703 35190
rect 7275 35010 7331 35066
rect 7399 35010 7455 35066
rect 7523 35010 7579 35066
rect 7647 35010 7703 35066
rect 7275 34886 7331 34942
rect 7399 34886 7455 34942
rect 7523 34886 7579 34942
rect 7647 34886 7703 34942
rect 7275 34762 7331 34818
rect 7399 34762 7455 34818
rect 7523 34762 7579 34818
rect 7647 34762 7703 34818
rect 7275 34638 7331 34694
rect 7399 34638 7455 34694
rect 7523 34638 7579 34694
rect 7647 34638 7703 34694
rect 7275 34514 7331 34570
rect 7399 34514 7455 34570
rect 7523 34514 7579 34570
rect 7647 34514 7703 34570
rect 7275 34390 7331 34446
rect 7399 34390 7455 34446
rect 7523 34390 7579 34446
rect 7647 34390 7703 34446
rect 7275 34266 7331 34322
rect 7399 34266 7455 34322
rect 7523 34266 7579 34322
rect 7647 34266 7703 34322
rect 7275 34142 7331 34198
rect 7399 34142 7455 34198
rect 7523 34142 7579 34198
rect 7647 34142 7703 34198
rect 7275 34018 7331 34074
rect 7399 34018 7455 34074
rect 7523 34018 7579 34074
rect 7647 34018 7703 34074
rect 7275 33894 7331 33950
rect 7399 33894 7455 33950
rect 7523 33894 7579 33950
rect 7647 33894 7703 33950
rect 7275 33770 7331 33826
rect 7399 33770 7455 33826
rect 7523 33770 7579 33826
rect 7647 33770 7703 33826
rect 7275 33646 7331 33702
rect 7399 33646 7455 33702
rect 7523 33646 7579 33702
rect 7647 33646 7703 33702
rect 9937 36498 9993 36554
rect 10061 36498 10117 36554
rect 9937 36374 9993 36430
rect 10061 36374 10117 36430
rect 9937 36250 9993 36306
rect 10061 36250 10117 36306
rect 9937 36126 9993 36182
rect 10061 36126 10117 36182
rect 9937 36002 9993 36058
rect 10061 36002 10117 36058
rect 9937 35878 9993 35934
rect 10061 35878 10117 35934
rect 9937 35754 9993 35810
rect 10061 35754 10117 35810
rect 9937 35630 9993 35686
rect 10061 35630 10117 35686
rect 9937 35506 9993 35562
rect 10061 35506 10117 35562
rect 9937 35382 9993 35438
rect 10061 35382 10117 35438
rect 9937 35258 9993 35314
rect 10061 35258 10117 35314
rect 9937 35134 9993 35190
rect 10061 35134 10117 35190
rect 9937 35010 9993 35066
rect 10061 35010 10117 35066
rect 9937 34886 9993 34942
rect 10061 34886 10117 34942
rect 9937 34762 9993 34818
rect 10061 34762 10117 34818
rect 9937 34638 9993 34694
rect 10061 34638 10117 34694
rect 9937 34514 9993 34570
rect 10061 34514 10117 34570
rect 9937 34390 9993 34446
rect 10061 34390 10117 34446
rect 9937 34266 9993 34322
rect 10061 34266 10117 34322
rect 9937 34142 9993 34198
rect 10061 34142 10117 34198
rect 9937 34018 9993 34074
rect 10061 34018 10117 34074
rect 9937 33894 9993 33950
rect 10061 33894 10117 33950
rect 9937 33770 9993 33826
rect 10061 33770 10117 33826
rect 9937 33646 9993 33702
rect 10061 33646 10117 33702
rect 12307 36498 12363 36554
rect 12431 36498 12487 36554
rect 12307 36374 12363 36430
rect 12431 36374 12487 36430
rect 12307 36250 12363 36306
rect 12431 36250 12487 36306
rect 12307 36126 12363 36182
rect 12431 36126 12487 36182
rect 12307 36002 12363 36058
rect 12431 36002 12487 36058
rect 12307 35878 12363 35934
rect 12431 35878 12487 35934
rect 12307 35754 12363 35810
rect 12431 35754 12487 35810
rect 12307 35630 12363 35686
rect 12431 35630 12487 35686
rect 12307 35506 12363 35562
rect 12431 35506 12487 35562
rect 12307 35382 12363 35438
rect 12431 35382 12487 35438
rect 12307 35258 12363 35314
rect 12431 35258 12487 35314
rect 12307 35134 12363 35190
rect 12431 35134 12487 35190
rect 12307 35010 12363 35066
rect 12431 35010 12487 35066
rect 12307 34886 12363 34942
rect 12431 34886 12487 34942
rect 12307 34762 12363 34818
rect 12431 34762 12487 34818
rect 12307 34638 12363 34694
rect 12431 34638 12487 34694
rect 12307 34514 12363 34570
rect 12431 34514 12487 34570
rect 12307 34390 12363 34446
rect 12431 34390 12487 34446
rect 12307 34266 12363 34322
rect 12431 34266 12487 34322
rect 12307 34142 12363 34198
rect 12431 34142 12487 34198
rect 12307 34018 12363 34074
rect 12431 34018 12487 34074
rect 12307 33894 12363 33950
rect 12431 33894 12487 33950
rect 12307 33770 12363 33826
rect 12431 33770 12487 33826
rect 12307 33646 12363 33702
rect 12431 33646 12487 33702
rect 315 33298 371 33354
rect 439 33298 495 33354
rect 563 33298 619 33354
rect 687 33298 743 33354
rect 811 33298 867 33354
rect 935 33298 991 33354
rect 1059 33298 1115 33354
rect 1183 33298 1239 33354
rect 1307 33298 1363 33354
rect 1431 33298 1487 33354
rect 1555 33298 1611 33354
rect 1679 33298 1735 33354
rect 1803 33298 1859 33354
rect 1927 33298 1983 33354
rect 2051 33298 2107 33354
rect 315 33174 371 33230
rect 439 33174 495 33230
rect 563 33174 619 33230
rect 687 33174 743 33230
rect 811 33174 867 33230
rect 935 33174 991 33230
rect 1059 33174 1115 33230
rect 1183 33174 1239 33230
rect 1307 33174 1363 33230
rect 1431 33174 1487 33230
rect 1555 33174 1611 33230
rect 1679 33174 1735 33230
rect 1803 33174 1859 33230
rect 1927 33174 1983 33230
rect 2051 33174 2107 33230
rect 315 33050 371 33106
rect 439 33050 495 33106
rect 563 33050 619 33106
rect 687 33050 743 33106
rect 811 33050 867 33106
rect 935 33050 991 33106
rect 1059 33050 1115 33106
rect 1183 33050 1239 33106
rect 1307 33050 1363 33106
rect 1431 33050 1487 33106
rect 1555 33050 1611 33106
rect 1679 33050 1735 33106
rect 1803 33050 1859 33106
rect 1927 33050 1983 33106
rect 2051 33050 2107 33106
rect 315 32926 371 32982
rect 439 32926 495 32982
rect 563 32926 619 32982
rect 687 32926 743 32982
rect 811 32926 867 32982
rect 935 32926 991 32982
rect 1059 32926 1115 32982
rect 1183 32926 1239 32982
rect 1307 32926 1363 32982
rect 1431 32926 1487 32982
rect 1555 32926 1611 32982
rect 1679 32926 1735 32982
rect 1803 32926 1859 32982
rect 1927 32926 1983 32982
rect 2051 32926 2107 32982
rect 315 32802 371 32858
rect 439 32802 495 32858
rect 563 32802 619 32858
rect 687 32802 743 32858
rect 811 32802 867 32858
rect 935 32802 991 32858
rect 1059 32802 1115 32858
rect 1183 32802 1239 32858
rect 1307 32802 1363 32858
rect 1431 32802 1487 32858
rect 1555 32802 1611 32858
rect 1679 32802 1735 32858
rect 1803 32802 1859 32858
rect 1927 32802 1983 32858
rect 2051 32802 2107 32858
rect 315 32678 371 32734
rect 439 32678 495 32734
rect 563 32678 619 32734
rect 687 32678 743 32734
rect 811 32678 867 32734
rect 935 32678 991 32734
rect 1059 32678 1115 32734
rect 1183 32678 1239 32734
rect 1307 32678 1363 32734
rect 1431 32678 1487 32734
rect 1555 32678 1611 32734
rect 1679 32678 1735 32734
rect 1803 32678 1859 32734
rect 1927 32678 1983 32734
rect 2051 32678 2107 32734
rect 315 32554 371 32610
rect 439 32554 495 32610
rect 563 32554 619 32610
rect 687 32554 743 32610
rect 811 32554 867 32610
rect 935 32554 991 32610
rect 1059 32554 1115 32610
rect 1183 32554 1239 32610
rect 1307 32554 1363 32610
rect 1431 32554 1487 32610
rect 1555 32554 1611 32610
rect 1679 32554 1735 32610
rect 1803 32554 1859 32610
rect 1927 32554 1983 32610
rect 2051 32554 2107 32610
rect 315 32430 371 32486
rect 439 32430 495 32486
rect 563 32430 619 32486
rect 687 32430 743 32486
rect 811 32430 867 32486
rect 935 32430 991 32486
rect 1059 32430 1115 32486
rect 1183 32430 1239 32486
rect 1307 32430 1363 32486
rect 1431 32430 1487 32486
rect 1555 32430 1611 32486
rect 1679 32430 1735 32486
rect 1803 32430 1859 32486
rect 1927 32430 1983 32486
rect 2051 32430 2107 32486
rect 315 32306 371 32362
rect 439 32306 495 32362
rect 563 32306 619 32362
rect 687 32306 743 32362
rect 811 32306 867 32362
rect 935 32306 991 32362
rect 1059 32306 1115 32362
rect 1183 32306 1239 32362
rect 1307 32306 1363 32362
rect 1431 32306 1487 32362
rect 1555 32306 1611 32362
rect 1679 32306 1735 32362
rect 1803 32306 1859 32362
rect 1927 32306 1983 32362
rect 2051 32306 2107 32362
rect 315 32182 371 32238
rect 439 32182 495 32238
rect 563 32182 619 32238
rect 687 32182 743 32238
rect 811 32182 867 32238
rect 935 32182 991 32238
rect 1059 32182 1115 32238
rect 1183 32182 1239 32238
rect 1307 32182 1363 32238
rect 1431 32182 1487 32238
rect 1555 32182 1611 32238
rect 1679 32182 1735 32238
rect 1803 32182 1859 32238
rect 1927 32182 1983 32238
rect 2051 32182 2107 32238
rect 315 32058 371 32114
rect 439 32058 495 32114
rect 563 32058 619 32114
rect 687 32058 743 32114
rect 811 32058 867 32114
rect 935 32058 991 32114
rect 1059 32058 1115 32114
rect 1183 32058 1239 32114
rect 1307 32058 1363 32114
rect 1431 32058 1487 32114
rect 1555 32058 1611 32114
rect 1679 32058 1735 32114
rect 1803 32058 1859 32114
rect 1927 32058 1983 32114
rect 2051 32058 2107 32114
rect 315 31934 371 31990
rect 439 31934 495 31990
rect 563 31934 619 31990
rect 687 31934 743 31990
rect 811 31934 867 31990
rect 935 31934 991 31990
rect 1059 31934 1115 31990
rect 1183 31934 1239 31990
rect 1307 31934 1363 31990
rect 1431 31934 1487 31990
rect 1555 31934 1611 31990
rect 1679 31934 1735 31990
rect 1803 31934 1859 31990
rect 1927 31934 1983 31990
rect 2051 31934 2107 31990
rect 315 31810 371 31866
rect 439 31810 495 31866
rect 563 31810 619 31866
rect 687 31810 743 31866
rect 811 31810 867 31866
rect 935 31810 991 31866
rect 1059 31810 1115 31866
rect 1183 31810 1239 31866
rect 1307 31810 1363 31866
rect 1431 31810 1487 31866
rect 1555 31810 1611 31866
rect 1679 31810 1735 31866
rect 1803 31810 1859 31866
rect 1927 31810 1983 31866
rect 2051 31810 2107 31866
rect 315 31686 371 31742
rect 439 31686 495 31742
rect 563 31686 619 31742
rect 687 31686 743 31742
rect 811 31686 867 31742
rect 935 31686 991 31742
rect 1059 31686 1115 31742
rect 1183 31686 1239 31742
rect 1307 31686 1363 31742
rect 1431 31686 1487 31742
rect 1555 31686 1611 31742
rect 1679 31686 1735 31742
rect 1803 31686 1859 31742
rect 1927 31686 1983 31742
rect 2051 31686 2107 31742
rect 315 31562 371 31618
rect 439 31562 495 31618
rect 563 31562 619 31618
rect 687 31562 743 31618
rect 811 31562 867 31618
rect 935 31562 991 31618
rect 1059 31562 1115 31618
rect 1183 31562 1239 31618
rect 1307 31562 1363 31618
rect 1431 31562 1487 31618
rect 1555 31562 1611 31618
rect 1679 31562 1735 31618
rect 1803 31562 1859 31618
rect 1927 31562 1983 31618
rect 2051 31562 2107 31618
rect 315 31438 371 31494
rect 439 31438 495 31494
rect 563 31438 619 31494
rect 687 31438 743 31494
rect 811 31438 867 31494
rect 935 31438 991 31494
rect 1059 31438 1115 31494
rect 1183 31438 1239 31494
rect 1307 31438 1363 31494
rect 1431 31438 1487 31494
rect 1555 31438 1611 31494
rect 1679 31438 1735 31494
rect 1803 31438 1859 31494
rect 1927 31438 1983 31494
rect 2051 31438 2107 31494
rect 315 31314 371 31370
rect 439 31314 495 31370
rect 563 31314 619 31370
rect 687 31314 743 31370
rect 811 31314 867 31370
rect 935 31314 991 31370
rect 1059 31314 1115 31370
rect 1183 31314 1239 31370
rect 1307 31314 1363 31370
rect 1431 31314 1487 31370
rect 1555 31314 1611 31370
rect 1679 31314 1735 31370
rect 1803 31314 1859 31370
rect 1927 31314 1983 31370
rect 2051 31314 2107 31370
rect 315 31190 371 31246
rect 439 31190 495 31246
rect 563 31190 619 31246
rect 687 31190 743 31246
rect 811 31190 867 31246
rect 935 31190 991 31246
rect 1059 31190 1115 31246
rect 1183 31190 1239 31246
rect 1307 31190 1363 31246
rect 1431 31190 1487 31246
rect 1555 31190 1611 31246
rect 1679 31190 1735 31246
rect 1803 31190 1859 31246
rect 1927 31190 1983 31246
rect 2051 31190 2107 31246
rect 315 31066 371 31122
rect 439 31066 495 31122
rect 563 31066 619 31122
rect 687 31066 743 31122
rect 811 31066 867 31122
rect 935 31066 991 31122
rect 1059 31066 1115 31122
rect 1183 31066 1239 31122
rect 1307 31066 1363 31122
rect 1431 31066 1487 31122
rect 1555 31066 1611 31122
rect 1679 31066 1735 31122
rect 1803 31066 1859 31122
rect 1927 31066 1983 31122
rect 2051 31066 2107 31122
rect 315 30942 371 30998
rect 439 30942 495 30998
rect 563 30942 619 30998
rect 687 30942 743 30998
rect 811 30942 867 30998
rect 935 30942 991 30998
rect 1059 30942 1115 30998
rect 1183 30942 1239 30998
rect 1307 30942 1363 30998
rect 1431 30942 1487 30998
rect 1555 30942 1611 30998
rect 1679 30942 1735 30998
rect 1803 30942 1859 30998
rect 1927 30942 1983 30998
rect 2051 30942 2107 30998
rect 315 30818 371 30874
rect 439 30818 495 30874
rect 563 30818 619 30874
rect 687 30818 743 30874
rect 811 30818 867 30874
rect 935 30818 991 30874
rect 1059 30818 1115 30874
rect 1183 30818 1239 30874
rect 1307 30818 1363 30874
rect 1431 30818 1487 30874
rect 1555 30818 1611 30874
rect 1679 30818 1735 30874
rect 1803 30818 1859 30874
rect 1927 30818 1983 30874
rect 2051 30818 2107 30874
rect 315 30694 371 30750
rect 439 30694 495 30750
rect 563 30694 619 30750
rect 687 30694 743 30750
rect 811 30694 867 30750
rect 935 30694 991 30750
rect 1059 30694 1115 30750
rect 1183 30694 1239 30750
rect 1307 30694 1363 30750
rect 1431 30694 1487 30750
rect 1555 30694 1611 30750
rect 1679 30694 1735 30750
rect 1803 30694 1859 30750
rect 1927 30694 1983 30750
rect 2051 30694 2107 30750
rect 315 30570 371 30626
rect 439 30570 495 30626
rect 563 30570 619 30626
rect 687 30570 743 30626
rect 811 30570 867 30626
rect 935 30570 991 30626
rect 1059 30570 1115 30626
rect 1183 30570 1239 30626
rect 1307 30570 1363 30626
rect 1431 30570 1487 30626
rect 1555 30570 1611 30626
rect 1679 30570 1735 30626
rect 1803 30570 1859 30626
rect 1927 30570 1983 30626
rect 2051 30570 2107 30626
rect 315 30446 371 30502
rect 439 30446 495 30502
rect 563 30446 619 30502
rect 687 30446 743 30502
rect 811 30446 867 30502
rect 935 30446 991 30502
rect 1059 30446 1115 30502
rect 1183 30446 1239 30502
rect 1307 30446 1363 30502
rect 1431 30446 1487 30502
rect 1555 30446 1611 30502
rect 1679 30446 1735 30502
rect 1803 30446 1859 30502
rect 1927 30446 1983 30502
rect 2051 30446 2107 30502
rect 2808 33298 2864 33354
rect 2932 33298 2988 33354
rect 3056 33298 3112 33354
rect 3180 33298 3236 33354
rect 3304 33298 3360 33354
rect 3428 33298 3484 33354
rect 3552 33298 3608 33354
rect 3676 33298 3732 33354
rect 3800 33298 3856 33354
rect 3924 33298 3980 33354
rect 4048 33298 4104 33354
rect 4172 33298 4228 33354
rect 4296 33298 4352 33354
rect 4420 33298 4476 33354
rect 4544 33298 4600 33354
rect 4668 33298 4724 33354
rect 2808 33174 2864 33230
rect 2932 33174 2988 33230
rect 3056 33174 3112 33230
rect 3180 33174 3236 33230
rect 3304 33174 3360 33230
rect 3428 33174 3484 33230
rect 3552 33174 3608 33230
rect 3676 33174 3732 33230
rect 3800 33174 3856 33230
rect 3924 33174 3980 33230
rect 4048 33174 4104 33230
rect 4172 33174 4228 33230
rect 4296 33174 4352 33230
rect 4420 33174 4476 33230
rect 4544 33174 4600 33230
rect 4668 33174 4724 33230
rect 2808 33050 2864 33106
rect 2932 33050 2988 33106
rect 3056 33050 3112 33106
rect 3180 33050 3236 33106
rect 3304 33050 3360 33106
rect 3428 33050 3484 33106
rect 3552 33050 3608 33106
rect 3676 33050 3732 33106
rect 3800 33050 3856 33106
rect 3924 33050 3980 33106
rect 4048 33050 4104 33106
rect 4172 33050 4228 33106
rect 4296 33050 4352 33106
rect 4420 33050 4476 33106
rect 4544 33050 4600 33106
rect 4668 33050 4724 33106
rect 2808 32926 2864 32982
rect 2932 32926 2988 32982
rect 3056 32926 3112 32982
rect 3180 32926 3236 32982
rect 3304 32926 3360 32982
rect 3428 32926 3484 32982
rect 3552 32926 3608 32982
rect 3676 32926 3732 32982
rect 3800 32926 3856 32982
rect 3924 32926 3980 32982
rect 4048 32926 4104 32982
rect 4172 32926 4228 32982
rect 4296 32926 4352 32982
rect 4420 32926 4476 32982
rect 4544 32926 4600 32982
rect 4668 32926 4724 32982
rect 2808 32802 2864 32858
rect 2932 32802 2988 32858
rect 3056 32802 3112 32858
rect 3180 32802 3236 32858
rect 3304 32802 3360 32858
rect 3428 32802 3484 32858
rect 3552 32802 3608 32858
rect 3676 32802 3732 32858
rect 3800 32802 3856 32858
rect 3924 32802 3980 32858
rect 4048 32802 4104 32858
rect 4172 32802 4228 32858
rect 4296 32802 4352 32858
rect 4420 32802 4476 32858
rect 4544 32802 4600 32858
rect 4668 32802 4724 32858
rect 2808 32678 2864 32734
rect 2932 32678 2988 32734
rect 3056 32678 3112 32734
rect 3180 32678 3236 32734
rect 3304 32678 3360 32734
rect 3428 32678 3484 32734
rect 3552 32678 3608 32734
rect 3676 32678 3732 32734
rect 3800 32678 3856 32734
rect 3924 32678 3980 32734
rect 4048 32678 4104 32734
rect 4172 32678 4228 32734
rect 4296 32678 4352 32734
rect 4420 32678 4476 32734
rect 4544 32678 4600 32734
rect 4668 32678 4724 32734
rect 2808 32554 2864 32610
rect 2932 32554 2988 32610
rect 3056 32554 3112 32610
rect 3180 32554 3236 32610
rect 3304 32554 3360 32610
rect 3428 32554 3484 32610
rect 3552 32554 3608 32610
rect 3676 32554 3732 32610
rect 3800 32554 3856 32610
rect 3924 32554 3980 32610
rect 4048 32554 4104 32610
rect 4172 32554 4228 32610
rect 4296 32554 4352 32610
rect 4420 32554 4476 32610
rect 4544 32554 4600 32610
rect 4668 32554 4724 32610
rect 2808 32430 2864 32486
rect 2932 32430 2988 32486
rect 3056 32430 3112 32486
rect 3180 32430 3236 32486
rect 3304 32430 3360 32486
rect 3428 32430 3484 32486
rect 3552 32430 3608 32486
rect 3676 32430 3732 32486
rect 3800 32430 3856 32486
rect 3924 32430 3980 32486
rect 4048 32430 4104 32486
rect 4172 32430 4228 32486
rect 4296 32430 4352 32486
rect 4420 32430 4476 32486
rect 4544 32430 4600 32486
rect 4668 32430 4724 32486
rect 2808 32306 2864 32362
rect 2932 32306 2988 32362
rect 3056 32306 3112 32362
rect 3180 32306 3236 32362
rect 3304 32306 3360 32362
rect 3428 32306 3484 32362
rect 3552 32306 3608 32362
rect 3676 32306 3732 32362
rect 3800 32306 3856 32362
rect 3924 32306 3980 32362
rect 4048 32306 4104 32362
rect 4172 32306 4228 32362
rect 4296 32306 4352 32362
rect 4420 32306 4476 32362
rect 4544 32306 4600 32362
rect 4668 32306 4724 32362
rect 2808 32182 2864 32238
rect 2932 32182 2988 32238
rect 3056 32182 3112 32238
rect 3180 32182 3236 32238
rect 3304 32182 3360 32238
rect 3428 32182 3484 32238
rect 3552 32182 3608 32238
rect 3676 32182 3732 32238
rect 3800 32182 3856 32238
rect 3924 32182 3980 32238
rect 4048 32182 4104 32238
rect 4172 32182 4228 32238
rect 4296 32182 4352 32238
rect 4420 32182 4476 32238
rect 4544 32182 4600 32238
rect 4668 32182 4724 32238
rect 2808 32058 2864 32114
rect 2932 32058 2988 32114
rect 3056 32058 3112 32114
rect 3180 32058 3236 32114
rect 3304 32058 3360 32114
rect 3428 32058 3484 32114
rect 3552 32058 3608 32114
rect 3676 32058 3732 32114
rect 3800 32058 3856 32114
rect 3924 32058 3980 32114
rect 4048 32058 4104 32114
rect 4172 32058 4228 32114
rect 4296 32058 4352 32114
rect 4420 32058 4476 32114
rect 4544 32058 4600 32114
rect 4668 32058 4724 32114
rect 2808 31934 2864 31990
rect 2932 31934 2988 31990
rect 3056 31934 3112 31990
rect 3180 31934 3236 31990
rect 3304 31934 3360 31990
rect 3428 31934 3484 31990
rect 3552 31934 3608 31990
rect 3676 31934 3732 31990
rect 3800 31934 3856 31990
rect 3924 31934 3980 31990
rect 4048 31934 4104 31990
rect 4172 31934 4228 31990
rect 4296 31934 4352 31990
rect 4420 31934 4476 31990
rect 4544 31934 4600 31990
rect 4668 31934 4724 31990
rect 2808 31810 2864 31866
rect 2932 31810 2988 31866
rect 3056 31810 3112 31866
rect 3180 31810 3236 31866
rect 3304 31810 3360 31866
rect 3428 31810 3484 31866
rect 3552 31810 3608 31866
rect 3676 31810 3732 31866
rect 3800 31810 3856 31866
rect 3924 31810 3980 31866
rect 4048 31810 4104 31866
rect 4172 31810 4228 31866
rect 4296 31810 4352 31866
rect 4420 31810 4476 31866
rect 4544 31810 4600 31866
rect 4668 31810 4724 31866
rect 2808 31686 2864 31742
rect 2932 31686 2988 31742
rect 3056 31686 3112 31742
rect 3180 31686 3236 31742
rect 3304 31686 3360 31742
rect 3428 31686 3484 31742
rect 3552 31686 3608 31742
rect 3676 31686 3732 31742
rect 3800 31686 3856 31742
rect 3924 31686 3980 31742
rect 4048 31686 4104 31742
rect 4172 31686 4228 31742
rect 4296 31686 4352 31742
rect 4420 31686 4476 31742
rect 4544 31686 4600 31742
rect 4668 31686 4724 31742
rect 2808 31562 2864 31618
rect 2932 31562 2988 31618
rect 3056 31562 3112 31618
rect 3180 31562 3236 31618
rect 3304 31562 3360 31618
rect 3428 31562 3484 31618
rect 3552 31562 3608 31618
rect 3676 31562 3732 31618
rect 3800 31562 3856 31618
rect 3924 31562 3980 31618
rect 4048 31562 4104 31618
rect 4172 31562 4228 31618
rect 4296 31562 4352 31618
rect 4420 31562 4476 31618
rect 4544 31562 4600 31618
rect 4668 31562 4724 31618
rect 2808 31438 2864 31494
rect 2932 31438 2988 31494
rect 3056 31438 3112 31494
rect 3180 31438 3236 31494
rect 3304 31438 3360 31494
rect 3428 31438 3484 31494
rect 3552 31438 3608 31494
rect 3676 31438 3732 31494
rect 3800 31438 3856 31494
rect 3924 31438 3980 31494
rect 4048 31438 4104 31494
rect 4172 31438 4228 31494
rect 4296 31438 4352 31494
rect 4420 31438 4476 31494
rect 4544 31438 4600 31494
rect 4668 31438 4724 31494
rect 2808 31314 2864 31370
rect 2932 31314 2988 31370
rect 3056 31314 3112 31370
rect 3180 31314 3236 31370
rect 3304 31314 3360 31370
rect 3428 31314 3484 31370
rect 3552 31314 3608 31370
rect 3676 31314 3732 31370
rect 3800 31314 3856 31370
rect 3924 31314 3980 31370
rect 4048 31314 4104 31370
rect 4172 31314 4228 31370
rect 4296 31314 4352 31370
rect 4420 31314 4476 31370
rect 4544 31314 4600 31370
rect 4668 31314 4724 31370
rect 2808 31190 2864 31246
rect 2932 31190 2988 31246
rect 3056 31190 3112 31246
rect 3180 31190 3236 31246
rect 3304 31190 3360 31246
rect 3428 31190 3484 31246
rect 3552 31190 3608 31246
rect 3676 31190 3732 31246
rect 3800 31190 3856 31246
rect 3924 31190 3980 31246
rect 4048 31190 4104 31246
rect 4172 31190 4228 31246
rect 4296 31190 4352 31246
rect 4420 31190 4476 31246
rect 4544 31190 4600 31246
rect 4668 31190 4724 31246
rect 2808 31066 2864 31122
rect 2932 31066 2988 31122
rect 3056 31066 3112 31122
rect 3180 31066 3236 31122
rect 3304 31066 3360 31122
rect 3428 31066 3484 31122
rect 3552 31066 3608 31122
rect 3676 31066 3732 31122
rect 3800 31066 3856 31122
rect 3924 31066 3980 31122
rect 4048 31066 4104 31122
rect 4172 31066 4228 31122
rect 4296 31066 4352 31122
rect 4420 31066 4476 31122
rect 4544 31066 4600 31122
rect 4668 31066 4724 31122
rect 2808 30942 2864 30998
rect 2932 30942 2988 30998
rect 3056 30942 3112 30998
rect 3180 30942 3236 30998
rect 3304 30942 3360 30998
rect 3428 30942 3484 30998
rect 3552 30942 3608 30998
rect 3676 30942 3732 30998
rect 3800 30942 3856 30998
rect 3924 30942 3980 30998
rect 4048 30942 4104 30998
rect 4172 30942 4228 30998
rect 4296 30942 4352 30998
rect 4420 30942 4476 30998
rect 4544 30942 4600 30998
rect 4668 30942 4724 30998
rect 2808 30818 2864 30874
rect 2932 30818 2988 30874
rect 3056 30818 3112 30874
rect 3180 30818 3236 30874
rect 3304 30818 3360 30874
rect 3428 30818 3484 30874
rect 3552 30818 3608 30874
rect 3676 30818 3732 30874
rect 3800 30818 3856 30874
rect 3924 30818 3980 30874
rect 4048 30818 4104 30874
rect 4172 30818 4228 30874
rect 4296 30818 4352 30874
rect 4420 30818 4476 30874
rect 4544 30818 4600 30874
rect 4668 30818 4724 30874
rect 2808 30694 2864 30750
rect 2932 30694 2988 30750
rect 3056 30694 3112 30750
rect 3180 30694 3236 30750
rect 3304 30694 3360 30750
rect 3428 30694 3484 30750
rect 3552 30694 3608 30750
rect 3676 30694 3732 30750
rect 3800 30694 3856 30750
rect 3924 30694 3980 30750
rect 4048 30694 4104 30750
rect 4172 30694 4228 30750
rect 4296 30694 4352 30750
rect 4420 30694 4476 30750
rect 4544 30694 4600 30750
rect 4668 30694 4724 30750
rect 2808 30570 2864 30626
rect 2932 30570 2988 30626
rect 3056 30570 3112 30626
rect 3180 30570 3236 30626
rect 3304 30570 3360 30626
rect 3428 30570 3484 30626
rect 3552 30570 3608 30626
rect 3676 30570 3732 30626
rect 3800 30570 3856 30626
rect 3924 30570 3980 30626
rect 4048 30570 4104 30626
rect 4172 30570 4228 30626
rect 4296 30570 4352 30626
rect 4420 30570 4476 30626
rect 4544 30570 4600 30626
rect 4668 30570 4724 30626
rect 2808 30446 2864 30502
rect 2932 30446 2988 30502
rect 3056 30446 3112 30502
rect 3180 30446 3236 30502
rect 3304 30446 3360 30502
rect 3428 30446 3484 30502
rect 3552 30446 3608 30502
rect 3676 30446 3732 30502
rect 3800 30446 3856 30502
rect 3924 30446 3980 30502
rect 4048 30446 4104 30502
rect 4172 30446 4228 30502
rect 4296 30446 4352 30502
rect 4420 30446 4476 30502
rect 4544 30446 4600 30502
rect 4668 30446 4724 30502
rect 5178 33298 5234 33354
rect 5302 33298 5358 33354
rect 5426 33298 5482 33354
rect 5550 33298 5606 33354
rect 5674 33298 5730 33354
rect 5798 33298 5854 33354
rect 5922 33298 5978 33354
rect 6046 33298 6102 33354
rect 6170 33298 6226 33354
rect 6294 33298 6350 33354
rect 6418 33298 6474 33354
rect 6542 33298 6598 33354
rect 6666 33298 6722 33354
rect 6790 33298 6846 33354
rect 6914 33298 6970 33354
rect 7038 33298 7094 33354
rect 5178 33174 5234 33230
rect 5302 33174 5358 33230
rect 5426 33174 5482 33230
rect 5550 33174 5606 33230
rect 5674 33174 5730 33230
rect 5798 33174 5854 33230
rect 5922 33174 5978 33230
rect 6046 33174 6102 33230
rect 6170 33174 6226 33230
rect 6294 33174 6350 33230
rect 6418 33174 6474 33230
rect 6542 33174 6598 33230
rect 6666 33174 6722 33230
rect 6790 33174 6846 33230
rect 6914 33174 6970 33230
rect 7038 33174 7094 33230
rect 5178 33050 5234 33106
rect 5302 33050 5358 33106
rect 5426 33050 5482 33106
rect 5550 33050 5606 33106
rect 5674 33050 5730 33106
rect 5798 33050 5854 33106
rect 5922 33050 5978 33106
rect 6046 33050 6102 33106
rect 6170 33050 6226 33106
rect 6294 33050 6350 33106
rect 6418 33050 6474 33106
rect 6542 33050 6598 33106
rect 6666 33050 6722 33106
rect 6790 33050 6846 33106
rect 6914 33050 6970 33106
rect 7038 33050 7094 33106
rect 5178 32926 5234 32982
rect 5302 32926 5358 32982
rect 5426 32926 5482 32982
rect 5550 32926 5606 32982
rect 5674 32926 5730 32982
rect 5798 32926 5854 32982
rect 5922 32926 5978 32982
rect 6046 32926 6102 32982
rect 6170 32926 6226 32982
rect 6294 32926 6350 32982
rect 6418 32926 6474 32982
rect 6542 32926 6598 32982
rect 6666 32926 6722 32982
rect 6790 32926 6846 32982
rect 6914 32926 6970 32982
rect 7038 32926 7094 32982
rect 5178 32802 5234 32858
rect 5302 32802 5358 32858
rect 5426 32802 5482 32858
rect 5550 32802 5606 32858
rect 5674 32802 5730 32858
rect 5798 32802 5854 32858
rect 5922 32802 5978 32858
rect 6046 32802 6102 32858
rect 6170 32802 6226 32858
rect 6294 32802 6350 32858
rect 6418 32802 6474 32858
rect 6542 32802 6598 32858
rect 6666 32802 6722 32858
rect 6790 32802 6846 32858
rect 6914 32802 6970 32858
rect 7038 32802 7094 32858
rect 5178 32678 5234 32734
rect 5302 32678 5358 32734
rect 5426 32678 5482 32734
rect 5550 32678 5606 32734
rect 5674 32678 5730 32734
rect 5798 32678 5854 32734
rect 5922 32678 5978 32734
rect 6046 32678 6102 32734
rect 6170 32678 6226 32734
rect 6294 32678 6350 32734
rect 6418 32678 6474 32734
rect 6542 32678 6598 32734
rect 6666 32678 6722 32734
rect 6790 32678 6846 32734
rect 6914 32678 6970 32734
rect 7038 32678 7094 32734
rect 5178 32554 5234 32610
rect 5302 32554 5358 32610
rect 5426 32554 5482 32610
rect 5550 32554 5606 32610
rect 5674 32554 5730 32610
rect 5798 32554 5854 32610
rect 5922 32554 5978 32610
rect 6046 32554 6102 32610
rect 6170 32554 6226 32610
rect 6294 32554 6350 32610
rect 6418 32554 6474 32610
rect 6542 32554 6598 32610
rect 6666 32554 6722 32610
rect 6790 32554 6846 32610
rect 6914 32554 6970 32610
rect 7038 32554 7094 32610
rect 5178 32430 5234 32486
rect 5302 32430 5358 32486
rect 5426 32430 5482 32486
rect 5550 32430 5606 32486
rect 5674 32430 5730 32486
rect 5798 32430 5854 32486
rect 5922 32430 5978 32486
rect 6046 32430 6102 32486
rect 6170 32430 6226 32486
rect 6294 32430 6350 32486
rect 6418 32430 6474 32486
rect 6542 32430 6598 32486
rect 6666 32430 6722 32486
rect 6790 32430 6846 32486
rect 6914 32430 6970 32486
rect 7038 32430 7094 32486
rect 5178 32306 5234 32362
rect 5302 32306 5358 32362
rect 5426 32306 5482 32362
rect 5550 32306 5606 32362
rect 5674 32306 5730 32362
rect 5798 32306 5854 32362
rect 5922 32306 5978 32362
rect 6046 32306 6102 32362
rect 6170 32306 6226 32362
rect 6294 32306 6350 32362
rect 6418 32306 6474 32362
rect 6542 32306 6598 32362
rect 6666 32306 6722 32362
rect 6790 32306 6846 32362
rect 6914 32306 6970 32362
rect 7038 32306 7094 32362
rect 5178 32182 5234 32238
rect 5302 32182 5358 32238
rect 5426 32182 5482 32238
rect 5550 32182 5606 32238
rect 5674 32182 5730 32238
rect 5798 32182 5854 32238
rect 5922 32182 5978 32238
rect 6046 32182 6102 32238
rect 6170 32182 6226 32238
rect 6294 32182 6350 32238
rect 6418 32182 6474 32238
rect 6542 32182 6598 32238
rect 6666 32182 6722 32238
rect 6790 32182 6846 32238
rect 6914 32182 6970 32238
rect 7038 32182 7094 32238
rect 5178 32058 5234 32114
rect 5302 32058 5358 32114
rect 5426 32058 5482 32114
rect 5550 32058 5606 32114
rect 5674 32058 5730 32114
rect 5798 32058 5854 32114
rect 5922 32058 5978 32114
rect 6046 32058 6102 32114
rect 6170 32058 6226 32114
rect 6294 32058 6350 32114
rect 6418 32058 6474 32114
rect 6542 32058 6598 32114
rect 6666 32058 6722 32114
rect 6790 32058 6846 32114
rect 6914 32058 6970 32114
rect 7038 32058 7094 32114
rect 5178 31934 5234 31990
rect 5302 31934 5358 31990
rect 5426 31934 5482 31990
rect 5550 31934 5606 31990
rect 5674 31934 5730 31990
rect 5798 31934 5854 31990
rect 5922 31934 5978 31990
rect 6046 31934 6102 31990
rect 6170 31934 6226 31990
rect 6294 31934 6350 31990
rect 6418 31934 6474 31990
rect 6542 31934 6598 31990
rect 6666 31934 6722 31990
rect 6790 31934 6846 31990
rect 6914 31934 6970 31990
rect 7038 31934 7094 31990
rect 5178 31810 5234 31866
rect 5302 31810 5358 31866
rect 5426 31810 5482 31866
rect 5550 31810 5606 31866
rect 5674 31810 5730 31866
rect 5798 31810 5854 31866
rect 5922 31810 5978 31866
rect 6046 31810 6102 31866
rect 6170 31810 6226 31866
rect 6294 31810 6350 31866
rect 6418 31810 6474 31866
rect 6542 31810 6598 31866
rect 6666 31810 6722 31866
rect 6790 31810 6846 31866
rect 6914 31810 6970 31866
rect 7038 31810 7094 31866
rect 5178 31686 5234 31742
rect 5302 31686 5358 31742
rect 5426 31686 5482 31742
rect 5550 31686 5606 31742
rect 5674 31686 5730 31742
rect 5798 31686 5854 31742
rect 5922 31686 5978 31742
rect 6046 31686 6102 31742
rect 6170 31686 6226 31742
rect 6294 31686 6350 31742
rect 6418 31686 6474 31742
rect 6542 31686 6598 31742
rect 6666 31686 6722 31742
rect 6790 31686 6846 31742
rect 6914 31686 6970 31742
rect 7038 31686 7094 31742
rect 5178 31562 5234 31618
rect 5302 31562 5358 31618
rect 5426 31562 5482 31618
rect 5550 31562 5606 31618
rect 5674 31562 5730 31618
rect 5798 31562 5854 31618
rect 5922 31562 5978 31618
rect 6046 31562 6102 31618
rect 6170 31562 6226 31618
rect 6294 31562 6350 31618
rect 6418 31562 6474 31618
rect 6542 31562 6598 31618
rect 6666 31562 6722 31618
rect 6790 31562 6846 31618
rect 6914 31562 6970 31618
rect 7038 31562 7094 31618
rect 5178 31438 5234 31494
rect 5302 31438 5358 31494
rect 5426 31438 5482 31494
rect 5550 31438 5606 31494
rect 5674 31438 5730 31494
rect 5798 31438 5854 31494
rect 5922 31438 5978 31494
rect 6046 31438 6102 31494
rect 6170 31438 6226 31494
rect 6294 31438 6350 31494
rect 6418 31438 6474 31494
rect 6542 31438 6598 31494
rect 6666 31438 6722 31494
rect 6790 31438 6846 31494
rect 6914 31438 6970 31494
rect 7038 31438 7094 31494
rect 5178 31314 5234 31370
rect 5302 31314 5358 31370
rect 5426 31314 5482 31370
rect 5550 31314 5606 31370
rect 5674 31314 5730 31370
rect 5798 31314 5854 31370
rect 5922 31314 5978 31370
rect 6046 31314 6102 31370
rect 6170 31314 6226 31370
rect 6294 31314 6350 31370
rect 6418 31314 6474 31370
rect 6542 31314 6598 31370
rect 6666 31314 6722 31370
rect 6790 31314 6846 31370
rect 6914 31314 6970 31370
rect 7038 31314 7094 31370
rect 5178 31190 5234 31246
rect 5302 31190 5358 31246
rect 5426 31190 5482 31246
rect 5550 31190 5606 31246
rect 5674 31190 5730 31246
rect 5798 31190 5854 31246
rect 5922 31190 5978 31246
rect 6046 31190 6102 31246
rect 6170 31190 6226 31246
rect 6294 31190 6350 31246
rect 6418 31190 6474 31246
rect 6542 31190 6598 31246
rect 6666 31190 6722 31246
rect 6790 31190 6846 31246
rect 6914 31190 6970 31246
rect 7038 31190 7094 31246
rect 5178 31066 5234 31122
rect 5302 31066 5358 31122
rect 5426 31066 5482 31122
rect 5550 31066 5606 31122
rect 5674 31066 5730 31122
rect 5798 31066 5854 31122
rect 5922 31066 5978 31122
rect 6046 31066 6102 31122
rect 6170 31066 6226 31122
rect 6294 31066 6350 31122
rect 6418 31066 6474 31122
rect 6542 31066 6598 31122
rect 6666 31066 6722 31122
rect 6790 31066 6846 31122
rect 6914 31066 6970 31122
rect 7038 31066 7094 31122
rect 5178 30942 5234 30998
rect 5302 30942 5358 30998
rect 5426 30942 5482 30998
rect 5550 30942 5606 30998
rect 5674 30942 5730 30998
rect 5798 30942 5854 30998
rect 5922 30942 5978 30998
rect 6046 30942 6102 30998
rect 6170 30942 6226 30998
rect 6294 30942 6350 30998
rect 6418 30942 6474 30998
rect 6542 30942 6598 30998
rect 6666 30942 6722 30998
rect 6790 30942 6846 30998
rect 6914 30942 6970 30998
rect 7038 30942 7094 30998
rect 5178 30818 5234 30874
rect 5302 30818 5358 30874
rect 5426 30818 5482 30874
rect 5550 30818 5606 30874
rect 5674 30818 5730 30874
rect 5798 30818 5854 30874
rect 5922 30818 5978 30874
rect 6046 30818 6102 30874
rect 6170 30818 6226 30874
rect 6294 30818 6350 30874
rect 6418 30818 6474 30874
rect 6542 30818 6598 30874
rect 6666 30818 6722 30874
rect 6790 30818 6846 30874
rect 6914 30818 6970 30874
rect 7038 30818 7094 30874
rect 5178 30694 5234 30750
rect 5302 30694 5358 30750
rect 5426 30694 5482 30750
rect 5550 30694 5606 30750
rect 5674 30694 5730 30750
rect 5798 30694 5854 30750
rect 5922 30694 5978 30750
rect 6046 30694 6102 30750
rect 6170 30694 6226 30750
rect 6294 30694 6350 30750
rect 6418 30694 6474 30750
rect 6542 30694 6598 30750
rect 6666 30694 6722 30750
rect 6790 30694 6846 30750
rect 6914 30694 6970 30750
rect 7038 30694 7094 30750
rect 5178 30570 5234 30626
rect 5302 30570 5358 30626
rect 5426 30570 5482 30626
rect 5550 30570 5606 30626
rect 5674 30570 5730 30626
rect 5798 30570 5854 30626
rect 5922 30570 5978 30626
rect 6046 30570 6102 30626
rect 6170 30570 6226 30626
rect 6294 30570 6350 30626
rect 6418 30570 6474 30626
rect 6542 30570 6598 30626
rect 6666 30570 6722 30626
rect 6790 30570 6846 30626
rect 6914 30570 6970 30626
rect 7038 30570 7094 30626
rect 5178 30446 5234 30502
rect 5302 30446 5358 30502
rect 5426 30446 5482 30502
rect 5550 30446 5606 30502
rect 5674 30446 5730 30502
rect 5798 30446 5854 30502
rect 5922 30446 5978 30502
rect 6046 30446 6102 30502
rect 6170 30446 6226 30502
rect 6294 30446 6350 30502
rect 6418 30446 6474 30502
rect 6542 30446 6598 30502
rect 6666 30446 6722 30502
rect 6790 30446 6846 30502
rect 6914 30446 6970 30502
rect 7038 30446 7094 30502
rect 7884 33298 7940 33354
rect 8008 33298 8064 33354
rect 8132 33298 8188 33354
rect 8256 33298 8312 33354
rect 8380 33298 8436 33354
rect 8504 33298 8560 33354
rect 8628 33298 8684 33354
rect 8752 33298 8808 33354
rect 8876 33298 8932 33354
rect 9000 33298 9056 33354
rect 9124 33298 9180 33354
rect 9248 33298 9304 33354
rect 9372 33298 9428 33354
rect 9496 33298 9552 33354
rect 9620 33298 9676 33354
rect 9744 33298 9800 33354
rect 7884 33174 7940 33230
rect 8008 33174 8064 33230
rect 8132 33174 8188 33230
rect 8256 33174 8312 33230
rect 8380 33174 8436 33230
rect 8504 33174 8560 33230
rect 8628 33174 8684 33230
rect 8752 33174 8808 33230
rect 8876 33174 8932 33230
rect 9000 33174 9056 33230
rect 9124 33174 9180 33230
rect 9248 33174 9304 33230
rect 9372 33174 9428 33230
rect 9496 33174 9552 33230
rect 9620 33174 9676 33230
rect 9744 33174 9800 33230
rect 7884 33050 7940 33106
rect 8008 33050 8064 33106
rect 8132 33050 8188 33106
rect 8256 33050 8312 33106
rect 8380 33050 8436 33106
rect 8504 33050 8560 33106
rect 8628 33050 8684 33106
rect 8752 33050 8808 33106
rect 8876 33050 8932 33106
rect 9000 33050 9056 33106
rect 9124 33050 9180 33106
rect 9248 33050 9304 33106
rect 9372 33050 9428 33106
rect 9496 33050 9552 33106
rect 9620 33050 9676 33106
rect 9744 33050 9800 33106
rect 7884 32926 7940 32982
rect 8008 32926 8064 32982
rect 8132 32926 8188 32982
rect 8256 32926 8312 32982
rect 8380 32926 8436 32982
rect 8504 32926 8560 32982
rect 8628 32926 8684 32982
rect 8752 32926 8808 32982
rect 8876 32926 8932 32982
rect 9000 32926 9056 32982
rect 9124 32926 9180 32982
rect 9248 32926 9304 32982
rect 9372 32926 9428 32982
rect 9496 32926 9552 32982
rect 9620 32926 9676 32982
rect 9744 32926 9800 32982
rect 7884 32802 7940 32858
rect 8008 32802 8064 32858
rect 8132 32802 8188 32858
rect 8256 32802 8312 32858
rect 8380 32802 8436 32858
rect 8504 32802 8560 32858
rect 8628 32802 8684 32858
rect 8752 32802 8808 32858
rect 8876 32802 8932 32858
rect 9000 32802 9056 32858
rect 9124 32802 9180 32858
rect 9248 32802 9304 32858
rect 9372 32802 9428 32858
rect 9496 32802 9552 32858
rect 9620 32802 9676 32858
rect 9744 32802 9800 32858
rect 7884 32678 7940 32734
rect 8008 32678 8064 32734
rect 8132 32678 8188 32734
rect 8256 32678 8312 32734
rect 8380 32678 8436 32734
rect 8504 32678 8560 32734
rect 8628 32678 8684 32734
rect 8752 32678 8808 32734
rect 8876 32678 8932 32734
rect 9000 32678 9056 32734
rect 9124 32678 9180 32734
rect 9248 32678 9304 32734
rect 9372 32678 9428 32734
rect 9496 32678 9552 32734
rect 9620 32678 9676 32734
rect 9744 32678 9800 32734
rect 7884 32554 7940 32610
rect 8008 32554 8064 32610
rect 8132 32554 8188 32610
rect 8256 32554 8312 32610
rect 8380 32554 8436 32610
rect 8504 32554 8560 32610
rect 8628 32554 8684 32610
rect 8752 32554 8808 32610
rect 8876 32554 8932 32610
rect 9000 32554 9056 32610
rect 9124 32554 9180 32610
rect 9248 32554 9304 32610
rect 9372 32554 9428 32610
rect 9496 32554 9552 32610
rect 9620 32554 9676 32610
rect 9744 32554 9800 32610
rect 7884 32430 7940 32486
rect 8008 32430 8064 32486
rect 8132 32430 8188 32486
rect 8256 32430 8312 32486
rect 8380 32430 8436 32486
rect 8504 32430 8560 32486
rect 8628 32430 8684 32486
rect 8752 32430 8808 32486
rect 8876 32430 8932 32486
rect 9000 32430 9056 32486
rect 9124 32430 9180 32486
rect 9248 32430 9304 32486
rect 9372 32430 9428 32486
rect 9496 32430 9552 32486
rect 9620 32430 9676 32486
rect 9744 32430 9800 32486
rect 7884 32306 7940 32362
rect 8008 32306 8064 32362
rect 8132 32306 8188 32362
rect 8256 32306 8312 32362
rect 8380 32306 8436 32362
rect 8504 32306 8560 32362
rect 8628 32306 8684 32362
rect 8752 32306 8808 32362
rect 8876 32306 8932 32362
rect 9000 32306 9056 32362
rect 9124 32306 9180 32362
rect 9248 32306 9304 32362
rect 9372 32306 9428 32362
rect 9496 32306 9552 32362
rect 9620 32306 9676 32362
rect 9744 32306 9800 32362
rect 7884 32182 7940 32238
rect 8008 32182 8064 32238
rect 8132 32182 8188 32238
rect 8256 32182 8312 32238
rect 8380 32182 8436 32238
rect 8504 32182 8560 32238
rect 8628 32182 8684 32238
rect 8752 32182 8808 32238
rect 8876 32182 8932 32238
rect 9000 32182 9056 32238
rect 9124 32182 9180 32238
rect 9248 32182 9304 32238
rect 9372 32182 9428 32238
rect 9496 32182 9552 32238
rect 9620 32182 9676 32238
rect 9744 32182 9800 32238
rect 7884 32058 7940 32114
rect 8008 32058 8064 32114
rect 8132 32058 8188 32114
rect 8256 32058 8312 32114
rect 8380 32058 8436 32114
rect 8504 32058 8560 32114
rect 8628 32058 8684 32114
rect 8752 32058 8808 32114
rect 8876 32058 8932 32114
rect 9000 32058 9056 32114
rect 9124 32058 9180 32114
rect 9248 32058 9304 32114
rect 9372 32058 9428 32114
rect 9496 32058 9552 32114
rect 9620 32058 9676 32114
rect 9744 32058 9800 32114
rect 7884 31934 7940 31990
rect 8008 31934 8064 31990
rect 8132 31934 8188 31990
rect 8256 31934 8312 31990
rect 8380 31934 8436 31990
rect 8504 31934 8560 31990
rect 8628 31934 8684 31990
rect 8752 31934 8808 31990
rect 8876 31934 8932 31990
rect 9000 31934 9056 31990
rect 9124 31934 9180 31990
rect 9248 31934 9304 31990
rect 9372 31934 9428 31990
rect 9496 31934 9552 31990
rect 9620 31934 9676 31990
rect 9744 31934 9800 31990
rect 7884 31810 7940 31866
rect 8008 31810 8064 31866
rect 8132 31810 8188 31866
rect 8256 31810 8312 31866
rect 8380 31810 8436 31866
rect 8504 31810 8560 31866
rect 8628 31810 8684 31866
rect 8752 31810 8808 31866
rect 8876 31810 8932 31866
rect 9000 31810 9056 31866
rect 9124 31810 9180 31866
rect 9248 31810 9304 31866
rect 9372 31810 9428 31866
rect 9496 31810 9552 31866
rect 9620 31810 9676 31866
rect 9744 31810 9800 31866
rect 7884 31686 7940 31742
rect 8008 31686 8064 31742
rect 8132 31686 8188 31742
rect 8256 31686 8312 31742
rect 8380 31686 8436 31742
rect 8504 31686 8560 31742
rect 8628 31686 8684 31742
rect 8752 31686 8808 31742
rect 8876 31686 8932 31742
rect 9000 31686 9056 31742
rect 9124 31686 9180 31742
rect 9248 31686 9304 31742
rect 9372 31686 9428 31742
rect 9496 31686 9552 31742
rect 9620 31686 9676 31742
rect 9744 31686 9800 31742
rect 7884 31562 7940 31618
rect 8008 31562 8064 31618
rect 8132 31562 8188 31618
rect 8256 31562 8312 31618
rect 8380 31562 8436 31618
rect 8504 31562 8560 31618
rect 8628 31562 8684 31618
rect 8752 31562 8808 31618
rect 8876 31562 8932 31618
rect 9000 31562 9056 31618
rect 9124 31562 9180 31618
rect 9248 31562 9304 31618
rect 9372 31562 9428 31618
rect 9496 31562 9552 31618
rect 9620 31562 9676 31618
rect 9744 31562 9800 31618
rect 7884 31438 7940 31494
rect 8008 31438 8064 31494
rect 8132 31438 8188 31494
rect 8256 31438 8312 31494
rect 8380 31438 8436 31494
rect 8504 31438 8560 31494
rect 8628 31438 8684 31494
rect 8752 31438 8808 31494
rect 8876 31438 8932 31494
rect 9000 31438 9056 31494
rect 9124 31438 9180 31494
rect 9248 31438 9304 31494
rect 9372 31438 9428 31494
rect 9496 31438 9552 31494
rect 9620 31438 9676 31494
rect 9744 31438 9800 31494
rect 7884 31314 7940 31370
rect 8008 31314 8064 31370
rect 8132 31314 8188 31370
rect 8256 31314 8312 31370
rect 8380 31314 8436 31370
rect 8504 31314 8560 31370
rect 8628 31314 8684 31370
rect 8752 31314 8808 31370
rect 8876 31314 8932 31370
rect 9000 31314 9056 31370
rect 9124 31314 9180 31370
rect 9248 31314 9304 31370
rect 9372 31314 9428 31370
rect 9496 31314 9552 31370
rect 9620 31314 9676 31370
rect 9744 31314 9800 31370
rect 7884 31190 7940 31246
rect 8008 31190 8064 31246
rect 8132 31190 8188 31246
rect 8256 31190 8312 31246
rect 8380 31190 8436 31246
rect 8504 31190 8560 31246
rect 8628 31190 8684 31246
rect 8752 31190 8808 31246
rect 8876 31190 8932 31246
rect 9000 31190 9056 31246
rect 9124 31190 9180 31246
rect 9248 31190 9304 31246
rect 9372 31190 9428 31246
rect 9496 31190 9552 31246
rect 9620 31190 9676 31246
rect 9744 31190 9800 31246
rect 7884 31066 7940 31122
rect 8008 31066 8064 31122
rect 8132 31066 8188 31122
rect 8256 31066 8312 31122
rect 8380 31066 8436 31122
rect 8504 31066 8560 31122
rect 8628 31066 8684 31122
rect 8752 31066 8808 31122
rect 8876 31066 8932 31122
rect 9000 31066 9056 31122
rect 9124 31066 9180 31122
rect 9248 31066 9304 31122
rect 9372 31066 9428 31122
rect 9496 31066 9552 31122
rect 9620 31066 9676 31122
rect 9744 31066 9800 31122
rect 7884 30942 7940 30998
rect 8008 30942 8064 30998
rect 8132 30942 8188 30998
rect 8256 30942 8312 30998
rect 8380 30942 8436 30998
rect 8504 30942 8560 30998
rect 8628 30942 8684 30998
rect 8752 30942 8808 30998
rect 8876 30942 8932 30998
rect 9000 30942 9056 30998
rect 9124 30942 9180 30998
rect 9248 30942 9304 30998
rect 9372 30942 9428 30998
rect 9496 30942 9552 30998
rect 9620 30942 9676 30998
rect 9744 30942 9800 30998
rect 7884 30818 7940 30874
rect 8008 30818 8064 30874
rect 8132 30818 8188 30874
rect 8256 30818 8312 30874
rect 8380 30818 8436 30874
rect 8504 30818 8560 30874
rect 8628 30818 8684 30874
rect 8752 30818 8808 30874
rect 8876 30818 8932 30874
rect 9000 30818 9056 30874
rect 9124 30818 9180 30874
rect 9248 30818 9304 30874
rect 9372 30818 9428 30874
rect 9496 30818 9552 30874
rect 9620 30818 9676 30874
rect 9744 30818 9800 30874
rect 7884 30694 7940 30750
rect 8008 30694 8064 30750
rect 8132 30694 8188 30750
rect 8256 30694 8312 30750
rect 8380 30694 8436 30750
rect 8504 30694 8560 30750
rect 8628 30694 8684 30750
rect 8752 30694 8808 30750
rect 8876 30694 8932 30750
rect 9000 30694 9056 30750
rect 9124 30694 9180 30750
rect 9248 30694 9304 30750
rect 9372 30694 9428 30750
rect 9496 30694 9552 30750
rect 9620 30694 9676 30750
rect 9744 30694 9800 30750
rect 7884 30570 7940 30626
rect 8008 30570 8064 30626
rect 8132 30570 8188 30626
rect 8256 30570 8312 30626
rect 8380 30570 8436 30626
rect 8504 30570 8560 30626
rect 8628 30570 8684 30626
rect 8752 30570 8808 30626
rect 8876 30570 8932 30626
rect 9000 30570 9056 30626
rect 9124 30570 9180 30626
rect 9248 30570 9304 30626
rect 9372 30570 9428 30626
rect 9496 30570 9552 30626
rect 9620 30570 9676 30626
rect 9744 30570 9800 30626
rect 7884 30446 7940 30502
rect 8008 30446 8064 30502
rect 8132 30446 8188 30502
rect 8256 30446 8312 30502
rect 8380 30446 8436 30502
rect 8504 30446 8560 30502
rect 8628 30446 8684 30502
rect 8752 30446 8808 30502
rect 8876 30446 8932 30502
rect 9000 30446 9056 30502
rect 9124 30446 9180 30502
rect 9248 30446 9304 30502
rect 9372 30446 9428 30502
rect 9496 30446 9552 30502
rect 9620 30446 9676 30502
rect 9744 30446 9800 30502
rect 10254 33298 10310 33354
rect 10378 33298 10434 33354
rect 10502 33298 10558 33354
rect 10626 33298 10682 33354
rect 10750 33298 10806 33354
rect 10874 33298 10930 33354
rect 10998 33298 11054 33354
rect 11122 33298 11178 33354
rect 11246 33298 11302 33354
rect 11370 33298 11426 33354
rect 11494 33298 11550 33354
rect 11618 33298 11674 33354
rect 11742 33298 11798 33354
rect 11866 33298 11922 33354
rect 11990 33298 12046 33354
rect 12114 33298 12170 33354
rect 10254 33174 10310 33230
rect 10378 33174 10434 33230
rect 10502 33174 10558 33230
rect 10626 33174 10682 33230
rect 10750 33174 10806 33230
rect 10874 33174 10930 33230
rect 10998 33174 11054 33230
rect 11122 33174 11178 33230
rect 11246 33174 11302 33230
rect 11370 33174 11426 33230
rect 11494 33174 11550 33230
rect 11618 33174 11674 33230
rect 11742 33174 11798 33230
rect 11866 33174 11922 33230
rect 11990 33174 12046 33230
rect 12114 33174 12170 33230
rect 10254 33050 10310 33106
rect 10378 33050 10434 33106
rect 10502 33050 10558 33106
rect 10626 33050 10682 33106
rect 10750 33050 10806 33106
rect 10874 33050 10930 33106
rect 10998 33050 11054 33106
rect 11122 33050 11178 33106
rect 11246 33050 11302 33106
rect 11370 33050 11426 33106
rect 11494 33050 11550 33106
rect 11618 33050 11674 33106
rect 11742 33050 11798 33106
rect 11866 33050 11922 33106
rect 11990 33050 12046 33106
rect 12114 33050 12170 33106
rect 10254 32926 10310 32982
rect 10378 32926 10434 32982
rect 10502 32926 10558 32982
rect 10626 32926 10682 32982
rect 10750 32926 10806 32982
rect 10874 32926 10930 32982
rect 10998 32926 11054 32982
rect 11122 32926 11178 32982
rect 11246 32926 11302 32982
rect 11370 32926 11426 32982
rect 11494 32926 11550 32982
rect 11618 32926 11674 32982
rect 11742 32926 11798 32982
rect 11866 32926 11922 32982
rect 11990 32926 12046 32982
rect 12114 32926 12170 32982
rect 10254 32802 10310 32858
rect 10378 32802 10434 32858
rect 10502 32802 10558 32858
rect 10626 32802 10682 32858
rect 10750 32802 10806 32858
rect 10874 32802 10930 32858
rect 10998 32802 11054 32858
rect 11122 32802 11178 32858
rect 11246 32802 11302 32858
rect 11370 32802 11426 32858
rect 11494 32802 11550 32858
rect 11618 32802 11674 32858
rect 11742 32802 11798 32858
rect 11866 32802 11922 32858
rect 11990 32802 12046 32858
rect 12114 32802 12170 32858
rect 10254 32678 10310 32734
rect 10378 32678 10434 32734
rect 10502 32678 10558 32734
rect 10626 32678 10682 32734
rect 10750 32678 10806 32734
rect 10874 32678 10930 32734
rect 10998 32678 11054 32734
rect 11122 32678 11178 32734
rect 11246 32678 11302 32734
rect 11370 32678 11426 32734
rect 11494 32678 11550 32734
rect 11618 32678 11674 32734
rect 11742 32678 11798 32734
rect 11866 32678 11922 32734
rect 11990 32678 12046 32734
rect 12114 32678 12170 32734
rect 10254 32554 10310 32610
rect 10378 32554 10434 32610
rect 10502 32554 10558 32610
rect 10626 32554 10682 32610
rect 10750 32554 10806 32610
rect 10874 32554 10930 32610
rect 10998 32554 11054 32610
rect 11122 32554 11178 32610
rect 11246 32554 11302 32610
rect 11370 32554 11426 32610
rect 11494 32554 11550 32610
rect 11618 32554 11674 32610
rect 11742 32554 11798 32610
rect 11866 32554 11922 32610
rect 11990 32554 12046 32610
rect 12114 32554 12170 32610
rect 10254 32430 10310 32486
rect 10378 32430 10434 32486
rect 10502 32430 10558 32486
rect 10626 32430 10682 32486
rect 10750 32430 10806 32486
rect 10874 32430 10930 32486
rect 10998 32430 11054 32486
rect 11122 32430 11178 32486
rect 11246 32430 11302 32486
rect 11370 32430 11426 32486
rect 11494 32430 11550 32486
rect 11618 32430 11674 32486
rect 11742 32430 11798 32486
rect 11866 32430 11922 32486
rect 11990 32430 12046 32486
rect 12114 32430 12170 32486
rect 10254 32306 10310 32362
rect 10378 32306 10434 32362
rect 10502 32306 10558 32362
rect 10626 32306 10682 32362
rect 10750 32306 10806 32362
rect 10874 32306 10930 32362
rect 10998 32306 11054 32362
rect 11122 32306 11178 32362
rect 11246 32306 11302 32362
rect 11370 32306 11426 32362
rect 11494 32306 11550 32362
rect 11618 32306 11674 32362
rect 11742 32306 11798 32362
rect 11866 32306 11922 32362
rect 11990 32306 12046 32362
rect 12114 32306 12170 32362
rect 10254 32182 10310 32238
rect 10378 32182 10434 32238
rect 10502 32182 10558 32238
rect 10626 32182 10682 32238
rect 10750 32182 10806 32238
rect 10874 32182 10930 32238
rect 10998 32182 11054 32238
rect 11122 32182 11178 32238
rect 11246 32182 11302 32238
rect 11370 32182 11426 32238
rect 11494 32182 11550 32238
rect 11618 32182 11674 32238
rect 11742 32182 11798 32238
rect 11866 32182 11922 32238
rect 11990 32182 12046 32238
rect 12114 32182 12170 32238
rect 10254 32058 10310 32114
rect 10378 32058 10434 32114
rect 10502 32058 10558 32114
rect 10626 32058 10682 32114
rect 10750 32058 10806 32114
rect 10874 32058 10930 32114
rect 10998 32058 11054 32114
rect 11122 32058 11178 32114
rect 11246 32058 11302 32114
rect 11370 32058 11426 32114
rect 11494 32058 11550 32114
rect 11618 32058 11674 32114
rect 11742 32058 11798 32114
rect 11866 32058 11922 32114
rect 11990 32058 12046 32114
rect 12114 32058 12170 32114
rect 10254 31934 10310 31990
rect 10378 31934 10434 31990
rect 10502 31934 10558 31990
rect 10626 31934 10682 31990
rect 10750 31934 10806 31990
rect 10874 31934 10930 31990
rect 10998 31934 11054 31990
rect 11122 31934 11178 31990
rect 11246 31934 11302 31990
rect 11370 31934 11426 31990
rect 11494 31934 11550 31990
rect 11618 31934 11674 31990
rect 11742 31934 11798 31990
rect 11866 31934 11922 31990
rect 11990 31934 12046 31990
rect 12114 31934 12170 31990
rect 10254 31810 10310 31866
rect 10378 31810 10434 31866
rect 10502 31810 10558 31866
rect 10626 31810 10682 31866
rect 10750 31810 10806 31866
rect 10874 31810 10930 31866
rect 10998 31810 11054 31866
rect 11122 31810 11178 31866
rect 11246 31810 11302 31866
rect 11370 31810 11426 31866
rect 11494 31810 11550 31866
rect 11618 31810 11674 31866
rect 11742 31810 11798 31866
rect 11866 31810 11922 31866
rect 11990 31810 12046 31866
rect 12114 31810 12170 31866
rect 10254 31686 10310 31742
rect 10378 31686 10434 31742
rect 10502 31686 10558 31742
rect 10626 31686 10682 31742
rect 10750 31686 10806 31742
rect 10874 31686 10930 31742
rect 10998 31686 11054 31742
rect 11122 31686 11178 31742
rect 11246 31686 11302 31742
rect 11370 31686 11426 31742
rect 11494 31686 11550 31742
rect 11618 31686 11674 31742
rect 11742 31686 11798 31742
rect 11866 31686 11922 31742
rect 11990 31686 12046 31742
rect 12114 31686 12170 31742
rect 10254 31562 10310 31618
rect 10378 31562 10434 31618
rect 10502 31562 10558 31618
rect 10626 31562 10682 31618
rect 10750 31562 10806 31618
rect 10874 31562 10930 31618
rect 10998 31562 11054 31618
rect 11122 31562 11178 31618
rect 11246 31562 11302 31618
rect 11370 31562 11426 31618
rect 11494 31562 11550 31618
rect 11618 31562 11674 31618
rect 11742 31562 11798 31618
rect 11866 31562 11922 31618
rect 11990 31562 12046 31618
rect 12114 31562 12170 31618
rect 10254 31438 10310 31494
rect 10378 31438 10434 31494
rect 10502 31438 10558 31494
rect 10626 31438 10682 31494
rect 10750 31438 10806 31494
rect 10874 31438 10930 31494
rect 10998 31438 11054 31494
rect 11122 31438 11178 31494
rect 11246 31438 11302 31494
rect 11370 31438 11426 31494
rect 11494 31438 11550 31494
rect 11618 31438 11674 31494
rect 11742 31438 11798 31494
rect 11866 31438 11922 31494
rect 11990 31438 12046 31494
rect 12114 31438 12170 31494
rect 10254 31314 10310 31370
rect 10378 31314 10434 31370
rect 10502 31314 10558 31370
rect 10626 31314 10682 31370
rect 10750 31314 10806 31370
rect 10874 31314 10930 31370
rect 10998 31314 11054 31370
rect 11122 31314 11178 31370
rect 11246 31314 11302 31370
rect 11370 31314 11426 31370
rect 11494 31314 11550 31370
rect 11618 31314 11674 31370
rect 11742 31314 11798 31370
rect 11866 31314 11922 31370
rect 11990 31314 12046 31370
rect 12114 31314 12170 31370
rect 10254 31190 10310 31246
rect 10378 31190 10434 31246
rect 10502 31190 10558 31246
rect 10626 31190 10682 31246
rect 10750 31190 10806 31246
rect 10874 31190 10930 31246
rect 10998 31190 11054 31246
rect 11122 31190 11178 31246
rect 11246 31190 11302 31246
rect 11370 31190 11426 31246
rect 11494 31190 11550 31246
rect 11618 31190 11674 31246
rect 11742 31190 11798 31246
rect 11866 31190 11922 31246
rect 11990 31190 12046 31246
rect 12114 31190 12170 31246
rect 10254 31066 10310 31122
rect 10378 31066 10434 31122
rect 10502 31066 10558 31122
rect 10626 31066 10682 31122
rect 10750 31066 10806 31122
rect 10874 31066 10930 31122
rect 10998 31066 11054 31122
rect 11122 31066 11178 31122
rect 11246 31066 11302 31122
rect 11370 31066 11426 31122
rect 11494 31066 11550 31122
rect 11618 31066 11674 31122
rect 11742 31066 11798 31122
rect 11866 31066 11922 31122
rect 11990 31066 12046 31122
rect 12114 31066 12170 31122
rect 10254 30942 10310 30998
rect 10378 30942 10434 30998
rect 10502 30942 10558 30998
rect 10626 30942 10682 30998
rect 10750 30942 10806 30998
rect 10874 30942 10930 30998
rect 10998 30942 11054 30998
rect 11122 30942 11178 30998
rect 11246 30942 11302 30998
rect 11370 30942 11426 30998
rect 11494 30942 11550 30998
rect 11618 30942 11674 30998
rect 11742 30942 11798 30998
rect 11866 30942 11922 30998
rect 11990 30942 12046 30998
rect 12114 30942 12170 30998
rect 10254 30818 10310 30874
rect 10378 30818 10434 30874
rect 10502 30818 10558 30874
rect 10626 30818 10682 30874
rect 10750 30818 10806 30874
rect 10874 30818 10930 30874
rect 10998 30818 11054 30874
rect 11122 30818 11178 30874
rect 11246 30818 11302 30874
rect 11370 30818 11426 30874
rect 11494 30818 11550 30874
rect 11618 30818 11674 30874
rect 11742 30818 11798 30874
rect 11866 30818 11922 30874
rect 11990 30818 12046 30874
rect 12114 30818 12170 30874
rect 10254 30694 10310 30750
rect 10378 30694 10434 30750
rect 10502 30694 10558 30750
rect 10626 30694 10682 30750
rect 10750 30694 10806 30750
rect 10874 30694 10930 30750
rect 10998 30694 11054 30750
rect 11122 30694 11178 30750
rect 11246 30694 11302 30750
rect 11370 30694 11426 30750
rect 11494 30694 11550 30750
rect 11618 30694 11674 30750
rect 11742 30694 11798 30750
rect 11866 30694 11922 30750
rect 11990 30694 12046 30750
rect 12114 30694 12170 30750
rect 10254 30570 10310 30626
rect 10378 30570 10434 30626
rect 10502 30570 10558 30626
rect 10626 30570 10682 30626
rect 10750 30570 10806 30626
rect 10874 30570 10930 30626
rect 10998 30570 11054 30626
rect 11122 30570 11178 30626
rect 11246 30570 11302 30626
rect 11370 30570 11426 30626
rect 11494 30570 11550 30626
rect 11618 30570 11674 30626
rect 11742 30570 11798 30626
rect 11866 30570 11922 30626
rect 11990 30570 12046 30626
rect 12114 30570 12170 30626
rect 10254 30446 10310 30502
rect 10378 30446 10434 30502
rect 10502 30446 10558 30502
rect 10626 30446 10682 30502
rect 10750 30446 10806 30502
rect 10874 30446 10930 30502
rect 10998 30446 11054 30502
rect 11122 30446 11178 30502
rect 11246 30446 11302 30502
rect 11370 30446 11426 30502
rect 11494 30446 11550 30502
rect 11618 30446 11674 30502
rect 11742 30446 11798 30502
rect 11866 30446 11922 30502
rect 11990 30446 12046 30502
rect 12114 30446 12170 30502
rect 12871 33298 12927 33354
rect 12995 33298 13051 33354
rect 13119 33298 13175 33354
rect 13243 33298 13299 33354
rect 13367 33298 13423 33354
rect 13491 33298 13547 33354
rect 13615 33298 13671 33354
rect 13739 33298 13795 33354
rect 13863 33298 13919 33354
rect 13987 33298 14043 33354
rect 14111 33298 14167 33354
rect 14235 33298 14291 33354
rect 14359 33298 14415 33354
rect 14483 33298 14539 33354
rect 14607 33298 14663 33354
rect 12871 33174 12927 33230
rect 12995 33174 13051 33230
rect 13119 33174 13175 33230
rect 13243 33174 13299 33230
rect 13367 33174 13423 33230
rect 13491 33174 13547 33230
rect 13615 33174 13671 33230
rect 13739 33174 13795 33230
rect 13863 33174 13919 33230
rect 13987 33174 14043 33230
rect 14111 33174 14167 33230
rect 14235 33174 14291 33230
rect 14359 33174 14415 33230
rect 14483 33174 14539 33230
rect 14607 33174 14663 33230
rect 12871 33050 12927 33106
rect 12995 33050 13051 33106
rect 13119 33050 13175 33106
rect 13243 33050 13299 33106
rect 13367 33050 13423 33106
rect 13491 33050 13547 33106
rect 13615 33050 13671 33106
rect 13739 33050 13795 33106
rect 13863 33050 13919 33106
rect 13987 33050 14043 33106
rect 14111 33050 14167 33106
rect 14235 33050 14291 33106
rect 14359 33050 14415 33106
rect 14483 33050 14539 33106
rect 14607 33050 14663 33106
rect 12871 32926 12927 32982
rect 12995 32926 13051 32982
rect 13119 32926 13175 32982
rect 13243 32926 13299 32982
rect 13367 32926 13423 32982
rect 13491 32926 13547 32982
rect 13615 32926 13671 32982
rect 13739 32926 13795 32982
rect 13863 32926 13919 32982
rect 13987 32926 14043 32982
rect 14111 32926 14167 32982
rect 14235 32926 14291 32982
rect 14359 32926 14415 32982
rect 14483 32926 14539 32982
rect 14607 32926 14663 32982
rect 12871 32802 12927 32858
rect 12995 32802 13051 32858
rect 13119 32802 13175 32858
rect 13243 32802 13299 32858
rect 13367 32802 13423 32858
rect 13491 32802 13547 32858
rect 13615 32802 13671 32858
rect 13739 32802 13795 32858
rect 13863 32802 13919 32858
rect 13987 32802 14043 32858
rect 14111 32802 14167 32858
rect 14235 32802 14291 32858
rect 14359 32802 14415 32858
rect 14483 32802 14539 32858
rect 14607 32802 14663 32858
rect 12871 32678 12927 32734
rect 12995 32678 13051 32734
rect 13119 32678 13175 32734
rect 13243 32678 13299 32734
rect 13367 32678 13423 32734
rect 13491 32678 13547 32734
rect 13615 32678 13671 32734
rect 13739 32678 13795 32734
rect 13863 32678 13919 32734
rect 13987 32678 14043 32734
rect 14111 32678 14167 32734
rect 14235 32678 14291 32734
rect 14359 32678 14415 32734
rect 14483 32678 14539 32734
rect 14607 32678 14663 32734
rect 12871 32554 12927 32610
rect 12995 32554 13051 32610
rect 13119 32554 13175 32610
rect 13243 32554 13299 32610
rect 13367 32554 13423 32610
rect 13491 32554 13547 32610
rect 13615 32554 13671 32610
rect 13739 32554 13795 32610
rect 13863 32554 13919 32610
rect 13987 32554 14043 32610
rect 14111 32554 14167 32610
rect 14235 32554 14291 32610
rect 14359 32554 14415 32610
rect 14483 32554 14539 32610
rect 14607 32554 14663 32610
rect 12871 32430 12927 32486
rect 12995 32430 13051 32486
rect 13119 32430 13175 32486
rect 13243 32430 13299 32486
rect 13367 32430 13423 32486
rect 13491 32430 13547 32486
rect 13615 32430 13671 32486
rect 13739 32430 13795 32486
rect 13863 32430 13919 32486
rect 13987 32430 14043 32486
rect 14111 32430 14167 32486
rect 14235 32430 14291 32486
rect 14359 32430 14415 32486
rect 14483 32430 14539 32486
rect 14607 32430 14663 32486
rect 12871 32306 12927 32362
rect 12995 32306 13051 32362
rect 13119 32306 13175 32362
rect 13243 32306 13299 32362
rect 13367 32306 13423 32362
rect 13491 32306 13547 32362
rect 13615 32306 13671 32362
rect 13739 32306 13795 32362
rect 13863 32306 13919 32362
rect 13987 32306 14043 32362
rect 14111 32306 14167 32362
rect 14235 32306 14291 32362
rect 14359 32306 14415 32362
rect 14483 32306 14539 32362
rect 14607 32306 14663 32362
rect 12871 32182 12927 32238
rect 12995 32182 13051 32238
rect 13119 32182 13175 32238
rect 13243 32182 13299 32238
rect 13367 32182 13423 32238
rect 13491 32182 13547 32238
rect 13615 32182 13671 32238
rect 13739 32182 13795 32238
rect 13863 32182 13919 32238
rect 13987 32182 14043 32238
rect 14111 32182 14167 32238
rect 14235 32182 14291 32238
rect 14359 32182 14415 32238
rect 14483 32182 14539 32238
rect 14607 32182 14663 32238
rect 12871 32058 12927 32114
rect 12995 32058 13051 32114
rect 13119 32058 13175 32114
rect 13243 32058 13299 32114
rect 13367 32058 13423 32114
rect 13491 32058 13547 32114
rect 13615 32058 13671 32114
rect 13739 32058 13795 32114
rect 13863 32058 13919 32114
rect 13987 32058 14043 32114
rect 14111 32058 14167 32114
rect 14235 32058 14291 32114
rect 14359 32058 14415 32114
rect 14483 32058 14539 32114
rect 14607 32058 14663 32114
rect 12871 31934 12927 31990
rect 12995 31934 13051 31990
rect 13119 31934 13175 31990
rect 13243 31934 13299 31990
rect 13367 31934 13423 31990
rect 13491 31934 13547 31990
rect 13615 31934 13671 31990
rect 13739 31934 13795 31990
rect 13863 31934 13919 31990
rect 13987 31934 14043 31990
rect 14111 31934 14167 31990
rect 14235 31934 14291 31990
rect 14359 31934 14415 31990
rect 14483 31934 14539 31990
rect 14607 31934 14663 31990
rect 12871 31810 12927 31866
rect 12995 31810 13051 31866
rect 13119 31810 13175 31866
rect 13243 31810 13299 31866
rect 13367 31810 13423 31866
rect 13491 31810 13547 31866
rect 13615 31810 13671 31866
rect 13739 31810 13795 31866
rect 13863 31810 13919 31866
rect 13987 31810 14043 31866
rect 14111 31810 14167 31866
rect 14235 31810 14291 31866
rect 14359 31810 14415 31866
rect 14483 31810 14539 31866
rect 14607 31810 14663 31866
rect 12871 31686 12927 31742
rect 12995 31686 13051 31742
rect 13119 31686 13175 31742
rect 13243 31686 13299 31742
rect 13367 31686 13423 31742
rect 13491 31686 13547 31742
rect 13615 31686 13671 31742
rect 13739 31686 13795 31742
rect 13863 31686 13919 31742
rect 13987 31686 14043 31742
rect 14111 31686 14167 31742
rect 14235 31686 14291 31742
rect 14359 31686 14415 31742
rect 14483 31686 14539 31742
rect 14607 31686 14663 31742
rect 12871 31562 12927 31618
rect 12995 31562 13051 31618
rect 13119 31562 13175 31618
rect 13243 31562 13299 31618
rect 13367 31562 13423 31618
rect 13491 31562 13547 31618
rect 13615 31562 13671 31618
rect 13739 31562 13795 31618
rect 13863 31562 13919 31618
rect 13987 31562 14043 31618
rect 14111 31562 14167 31618
rect 14235 31562 14291 31618
rect 14359 31562 14415 31618
rect 14483 31562 14539 31618
rect 14607 31562 14663 31618
rect 12871 31438 12927 31494
rect 12995 31438 13051 31494
rect 13119 31438 13175 31494
rect 13243 31438 13299 31494
rect 13367 31438 13423 31494
rect 13491 31438 13547 31494
rect 13615 31438 13671 31494
rect 13739 31438 13795 31494
rect 13863 31438 13919 31494
rect 13987 31438 14043 31494
rect 14111 31438 14167 31494
rect 14235 31438 14291 31494
rect 14359 31438 14415 31494
rect 14483 31438 14539 31494
rect 14607 31438 14663 31494
rect 12871 31314 12927 31370
rect 12995 31314 13051 31370
rect 13119 31314 13175 31370
rect 13243 31314 13299 31370
rect 13367 31314 13423 31370
rect 13491 31314 13547 31370
rect 13615 31314 13671 31370
rect 13739 31314 13795 31370
rect 13863 31314 13919 31370
rect 13987 31314 14043 31370
rect 14111 31314 14167 31370
rect 14235 31314 14291 31370
rect 14359 31314 14415 31370
rect 14483 31314 14539 31370
rect 14607 31314 14663 31370
rect 12871 31190 12927 31246
rect 12995 31190 13051 31246
rect 13119 31190 13175 31246
rect 13243 31190 13299 31246
rect 13367 31190 13423 31246
rect 13491 31190 13547 31246
rect 13615 31190 13671 31246
rect 13739 31190 13795 31246
rect 13863 31190 13919 31246
rect 13987 31190 14043 31246
rect 14111 31190 14167 31246
rect 14235 31190 14291 31246
rect 14359 31190 14415 31246
rect 14483 31190 14539 31246
rect 14607 31190 14663 31246
rect 12871 31066 12927 31122
rect 12995 31066 13051 31122
rect 13119 31066 13175 31122
rect 13243 31066 13299 31122
rect 13367 31066 13423 31122
rect 13491 31066 13547 31122
rect 13615 31066 13671 31122
rect 13739 31066 13795 31122
rect 13863 31066 13919 31122
rect 13987 31066 14043 31122
rect 14111 31066 14167 31122
rect 14235 31066 14291 31122
rect 14359 31066 14415 31122
rect 14483 31066 14539 31122
rect 14607 31066 14663 31122
rect 12871 30942 12927 30998
rect 12995 30942 13051 30998
rect 13119 30942 13175 30998
rect 13243 30942 13299 30998
rect 13367 30942 13423 30998
rect 13491 30942 13547 30998
rect 13615 30942 13671 30998
rect 13739 30942 13795 30998
rect 13863 30942 13919 30998
rect 13987 30942 14043 30998
rect 14111 30942 14167 30998
rect 14235 30942 14291 30998
rect 14359 30942 14415 30998
rect 14483 30942 14539 30998
rect 14607 30942 14663 30998
rect 12871 30818 12927 30874
rect 12995 30818 13051 30874
rect 13119 30818 13175 30874
rect 13243 30818 13299 30874
rect 13367 30818 13423 30874
rect 13491 30818 13547 30874
rect 13615 30818 13671 30874
rect 13739 30818 13795 30874
rect 13863 30818 13919 30874
rect 13987 30818 14043 30874
rect 14111 30818 14167 30874
rect 14235 30818 14291 30874
rect 14359 30818 14415 30874
rect 14483 30818 14539 30874
rect 14607 30818 14663 30874
rect 12871 30694 12927 30750
rect 12995 30694 13051 30750
rect 13119 30694 13175 30750
rect 13243 30694 13299 30750
rect 13367 30694 13423 30750
rect 13491 30694 13547 30750
rect 13615 30694 13671 30750
rect 13739 30694 13795 30750
rect 13863 30694 13919 30750
rect 13987 30694 14043 30750
rect 14111 30694 14167 30750
rect 14235 30694 14291 30750
rect 14359 30694 14415 30750
rect 14483 30694 14539 30750
rect 14607 30694 14663 30750
rect 12871 30570 12927 30626
rect 12995 30570 13051 30626
rect 13119 30570 13175 30626
rect 13243 30570 13299 30626
rect 13367 30570 13423 30626
rect 13491 30570 13547 30626
rect 13615 30570 13671 30626
rect 13739 30570 13795 30626
rect 13863 30570 13919 30626
rect 13987 30570 14043 30626
rect 14111 30570 14167 30626
rect 14235 30570 14291 30626
rect 14359 30570 14415 30626
rect 14483 30570 14539 30626
rect 14607 30570 14663 30626
rect 12871 30446 12927 30502
rect 12995 30446 13051 30502
rect 13119 30446 13175 30502
rect 13243 30446 13299 30502
rect 13367 30446 13423 30502
rect 13491 30446 13547 30502
rect 13615 30446 13671 30502
rect 13739 30446 13795 30502
rect 13863 30446 13919 30502
rect 13987 30446 14043 30502
rect 14111 30446 14167 30502
rect 14235 30446 14291 30502
rect 14359 30446 14415 30502
rect 14483 30446 14539 30502
rect 14607 30446 14663 30502
rect 315 30092 371 30148
rect 439 30092 495 30148
rect 563 30092 619 30148
rect 687 30092 743 30148
rect 811 30092 867 30148
rect 935 30092 991 30148
rect 1059 30092 1115 30148
rect 1183 30092 1239 30148
rect 1307 30092 1363 30148
rect 1431 30092 1487 30148
rect 1555 30092 1611 30148
rect 1679 30092 1735 30148
rect 1803 30092 1859 30148
rect 1927 30092 1983 30148
rect 2051 30092 2107 30148
rect 315 29968 371 30024
rect 439 29968 495 30024
rect 563 29968 619 30024
rect 687 29968 743 30024
rect 811 29968 867 30024
rect 935 29968 991 30024
rect 1059 29968 1115 30024
rect 1183 29968 1239 30024
rect 1307 29968 1363 30024
rect 1431 29968 1487 30024
rect 1555 29968 1611 30024
rect 1679 29968 1735 30024
rect 1803 29968 1859 30024
rect 1927 29968 1983 30024
rect 2051 29968 2107 30024
rect 315 29844 371 29900
rect 439 29844 495 29900
rect 563 29844 619 29900
rect 687 29844 743 29900
rect 811 29844 867 29900
rect 935 29844 991 29900
rect 1059 29844 1115 29900
rect 1183 29844 1239 29900
rect 1307 29844 1363 29900
rect 1431 29844 1487 29900
rect 1555 29844 1611 29900
rect 1679 29844 1735 29900
rect 1803 29844 1859 29900
rect 1927 29844 1983 29900
rect 2051 29844 2107 29900
rect 315 29720 371 29776
rect 439 29720 495 29776
rect 563 29720 619 29776
rect 687 29720 743 29776
rect 811 29720 867 29776
rect 935 29720 991 29776
rect 1059 29720 1115 29776
rect 1183 29720 1239 29776
rect 1307 29720 1363 29776
rect 1431 29720 1487 29776
rect 1555 29720 1611 29776
rect 1679 29720 1735 29776
rect 1803 29720 1859 29776
rect 1927 29720 1983 29776
rect 2051 29720 2107 29776
rect 315 29596 371 29652
rect 439 29596 495 29652
rect 563 29596 619 29652
rect 687 29596 743 29652
rect 811 29596 867 29652
rect 935 29596 991 29652
rect 1059 29596 1115 29652
rect 1183 29596 1239 29652
rect 1307 29596 1363 29652
rect 1431 29596 1487 29652
rect 1555 29596 1611 29652
rect 1679 29596 1735 29652
rect 1803 29596 1859 29652
rect 1927 29596 1983 29652
rect 2051 29596 2107 29652
rect 315 29472 371 29528
rect 439 29472 495 29528
rect 563 29472 619 29528
rect 687 29472 743 29528
rect 811 29472 867 29528
rect 935 29472 991 29528
rect 1059 29472 1115 29528
rect 1183 29472 1239 29528
rect 1307 29472 1363 29528
rect 1431 29472 1487 29528
rect 1555 29472 1611 29528
rect 1679 29472 1735 29528
rect 1803 29472 1859 29528
rect 1927 29472 1983 29528
rect 2051 29472 2107 29528
rect 315 29348 371 29404
rect 439 29348 495 29404
rect 563 29348 619 29404
rect 687 29348 743 29404
rect 811 29348 867 29404
rect 935 29348 991 29404
rect 1059 29348 1115 29404
rect 1183 29348 1239 29404
rect 1307 29348 1363 29404
rect 1431 29348 1487 29404
rect 1555 29348 1611 29404
rect 1679 29348 1735 29404
rect 1803 29348 1859 29404
rect 1927 29348 1983 29404
rect 2051 29348 2107 29404
rect 315 29224 371 29280
rect 439 29224 495 29280
rect 563 29224 619 29280
rect 687 29224 743 29280
rect 811 29224 867 29280
rect 935 29224 991 29280
rect 1059 29224 1115 29280
rect 1183 29224 1239 29280
rect 1307 29224 1363 29280
rect 1431 29224 1487 29280
rect 1555 29224 1611 29280
rect 1679 29224 1735 29280
rect 1803 29224 1859 29280
rect 1927 29224 1983 29280
rect 2051 29224 2107 29280
rect 315 29100 371 29156
rect 439 29100 495 29156
rect 563 29100 619 29156
rect 687 29100 743 29156
rect 811 29100 867 29156
rect 935 29100 991 29156
rect 1059 29100 1115 29156
rect 1183 29100 1239 29156
rect 1307 29100 1363 29156
rect 1431 29100 1487 29156
rect 1555 29100 1611 29156
rect 1679 29100 1735 29156
rect 1803 29100 1859 29156
rect 1927 29100 1983 29156
rect 2051 29100 2107 29156
rect 315 28976 371 29032
rect 439 28976 495 29032
rect 563 28976 619 29032
rect 687 28976 743 29032
rect 811 28976 867 29032
rect 935 28976 991 29032
rect 1059 28976 1115 29032
rect 1183 28976 1239 29032
rect 1307 28976 1363 29032
rect 1431 28976 1487 29032
rect 1555 28976 1611 29032
rect 1679 28976 1735 29032
rect 1803 28976 1859 29032
rect 1927 28976 1983 29032
rect 2051 28976 2107 29032
rect 315 28852 371 28908
rect 439 28852 495 28908
rect 563 28852 619 28908
rect 687 28852 743 28908
rect 811 28852 867 28908
rect 935 28852 991 28908
rect 1059 28852 1115 28908
rect 1183 28852 1239 28908
rect 1307 28852 1363 28908
rect 1431 28852 1487 28908
rect 1555 28852 1611 28908
rect 1679 28852 1735 28908
rect 1803 28852 1859 28908
rect 1927 28852 1983 28908
rect 2051 28852 2107 28908
rect 2808 30092 2864 30148
rect 2932 30092 2988 30148
rect 3056 30092 3112 30148
rect 3180 30092 3236 30148
rect 3304 30092 3360 30148
rect 3428 30092 3484 30148
rect 3552 30092 3608 30148
rect 3676 30092 3732 30148
rect 3800 30092 3856 30148
rect 3924 30092 3980 30148
rect 4048 30092 4104 30148
rect 4172 30092 4228 30148
rect 4296 30092 4352 30148
rect 4420 30092 4476 30148
rect 4544 30092 4600 30148
rect 4668 30092 4724 30148
rect 2808 29968 2864 30024
rect 2932 29968 2988 30024
rect 3056 29968 3112 30024
rect 3180 29968 3236 30024
rect 3304 29968 3360 30024
rect 3428 29968 3484 30024
rect 3552 29968 3608 30024
rect 3676 29968 3732 30024
rect 3800 29968 3856 30024
rect 3924 29968 3980 30024
rect 4048 29968 4104 30024
rect 4172 29968 4228 30024
rect 4296 29968 4352 30024
rect 4420 29968 4476 30024
rect 4544 29968 4600 30024
rect 4668 29968 4724 30024
rect 2808 29844 2864 29900
rect 2932 29844 2988 29900
rect 3056 29844 3112 29900
rect 3180 29844 3236 29900
rect 3304 29844 3360 29900
rect 3428 29844 3484 29900
rect 3552 29844 3608 29900
rect 3676 29844 3732 29900
rect 3800 29844 3856 29900
rect 3924 29844 3980 29900
rect 4048 29844 4104 29900
rect 4172 29844 4228 29900
rect 4296 29844 4352 29900
rect 4420 29844 4476 29900
rect 4544 29844 4600 29900
rect 4668 29844 4724 29900
rect 2808 29720 2864 29776
rect 2932 29720 2988 29776
rect 3056 29720 3112 29776
rect 3180 29720 3236 29776
rect 3304 29720 3360 29776
rect 3428 29720 3484 29776
rect 3552 29720 3608 29776
rect 3676 29720 3732 29776
rect 3800 29720 3856 29776
rect 3924 29720 3980 29776
rect 4048 29720 4104 29776
rect 4172 29720 4228 29776
rect 4296 29720 4352 29776
rect 4420 29720 4476 29776
rect 4544 29720 4600 29776
rect 4668 29720 4724 29776
rect 2808 29596 2864 29652
rect 2932 29596 2988 29652
rect 3056 29596 3112 29652
rect 3180 29596 3236 29652
rect 3304 29596 3360 29652
rect 3428 29596 3484 29652
rect 3552 29596 3608 29652
rect 3676 29596 3732 29652
rect 3800 29596 3856 29652
rect 3924 29596 3980 29652
rect 4048 29596 4104 29652
rect 4172 29596 4228 29652
rect 4296 29596 4352 29652
rect 4420 29596 4476 29652
rect 4544 29596 4600 29652
rect 4668 29596 4724 29652
rect 2808 29472 2864 29528
rect 2932 29472 2988 29528
rect 3056 29472 3112 29528
rect 3180 29472 3236 29528
rect 3304 29472 3360 29528
rect 3428 29472 3484 29528
rect 3552 29472 3608 29528
rect 3676 29472 3732 29528
rect 3800 29472 3856 29528
rect 3924 29472 3980 29528
rect 4048 29472 4104 29528
rect 4172 29472 4228 29528
rect 4296 29472 4352 29528
rect 4420 29472 4476 29528
rect 4544 29472 4600 29528
rect 4668 29472 4724 29528
rect 2808 29348 2864 29404
rect 2932 29348 2988 29404
rect 3056 29348 3112 29404
rect 3180 29348 3236 29404
rect 3304 29348 3360 29404
rect 3428 29348 3484 29404
rect 3552 29348 3608 29404
rect 3676 29348 3732 29404
rect 3800 29348 3856 29404
rect 3924 29348 3980 29404
rect 4048 29348 4104 29404
rect 4172 29348 4228 29404
rect 4296 29348 4352 29404
rect 4420 29348 4476 29404
rect 4544 29348 4600 29404
rect 4668 29348 4724 29404
rect 2808 29224 2864 29280
rect 2932 29224 2988 29280
rect 3056 29224 3112 29280
rect 3180 29224 3236 29280
rect 3304 29224 3360 29280
rect 3428 29224 3484 29280
rect 3552 29224 3608 29280
rect 3676 29224 3732 29280
rect 3800 29224 3856 29280
rect 3924 29224 3980 29280
rect 4048 29224 4104 29280
rect 4172 29224 4228 29280
rect 4296 29224 4352 29280
rect 4420 29224 4476 29280
rect 4544 29224 4600 29280
rect 4668 29224 4724 29280
rect 2808 29100 2864 29156
rect 2932 29100 2988 29156
rect 3056 29100 3112 29156
rect 3180 29100 3236 29156
rect 3304 29100 3360 29156
rect 3428 29100 3484 29156
rect 3552 29100 3608 29156
rect 3676 29100 3732 29156
rect 3800 29100 3856 29156
rect 3924 29100 3980 29156
rect 4048 29100 4104 29156
rect 4172 29100 4228 29156
rect 4296 29100 4352 29156
rect 4420 29100 4476 29156
rect 4544 29100 4600 29156
rect 4668 29100 4724 29156
rect 2808 28976 2864 29032
rect 2932 28976 2988 29032
rect 3056 28976 3112 29032
rect 3180 28976 3236 29032
rect 3304 28976 3360 29032
rect 3428 28976 3484 29032
rect 3552 28976 3608 29032
rect 3676 28976 3732 29032
rect 3800 28976 3856 29032
rect 3924 28976 3980 29032
rect 4048 28976 4104 29032
rect 4172 28976 4228 29032
rect 4296 28976 4352 29032
rect 4420 28976 4476 29032
rect 4544 28976 4600 29032
rect 4668 28976 4724 29032
rect 2808 28852 2864 28908
rect 2932 28852 2988 28908
rect 3056 28852 3112 28908
rect 3180 28852 3236 28908
rect 3304 28852 3360 28908
rect 3428 28852 3484 28908
rect 3552 28852 3608 28908
rect 3676 28852 3732 28908
rect 3800 28852 3856 28908
rect 3924 28852 3980 28908
rect 4048 28852 4104 28908
rect 4172 28852 4228 28908
rect 4296 28852 4352 28908
rect 4420 28852 4476 28908
rect 4544 28852 4600 28908
rect 4668 28852 4724 28908
rect 5178 30092 5234 30148
rect 5302 30092 5358 30148
rect 5426 30092 5482 30148
rect 5550 30092 5606 30148
rect 5674 30092 5730 30148
rect 5798 30092 5854 30148
rect 5922 30092 5978 30148
rect 6046 30092 6102 30148
rect 6170 30092 6226 30148
rect 6294 30092 6350 30148
rect 6418 30092 6474 30148
rect 6542 30092 6598 30148
rect 6666 30092 6722 30148
rect 6790 30092 6846 30148
rect 6914 30092 6970 30148
rect 7038 30092 7094 30148
rect 5178 29968 5234 30024
rect 5302 29968 5358 30024
rect 5426 29968 5482 30024
rect 5550 29968 5606 30024
rect 5674 29968 5730 30024
rect 5798 29968 5854 30024
rect 5922 29968 5978 30024
rect 6046 29968 6102 30024
rect 6170 29968 6226 30024
rect 6294 29968 6350 30024
rect 6418 29968 6474 30024
rect 6542 29968 6598 30024
rect 6666 29968 6722 30024
rect 6790 29968 6846 30024
rect 6914 29968 6970 30024
rect 7038 29968 7094 30024
rect 5178 29844 5234 29900
rect 5302 29844 5358 29900
rect 5426 29844 5482 29900
rect 5550 29844 5606 29900
rect 5674 29844 5730 29900
rect 5798 29844 5854 29900
rect 5922 29844 5978 29900
rect 6046 29844 6102 29900
rect 6170 29844 6226 29900
rect 6294 29844 6350 29900
rect 6418 29844 6474 29900
rect 6542 29844 6598 29900
rect 6666 29844 6722 29900
rect 6790 29844 6846 29900
rect 6914 29844 6970 29900
rect 7038 29844 7094 29900
rect 5178 29720 5234 29776
rect 5302 29720 5358 29776
rect 5426 29720 5482 29776
rect 5550 29720 5606 29776
rect 5674 29720 5730 29776
rect 5798 29720 5854 29776
rect 5922 29720 5978 29776
rect 6046 29720 6102 29776
rect 6170 29720 6226 29776
rect 6294 29720 6350 29776
rect 6418 29720 6474 29776
rect 6542 29720 6598 29776
rect 6666 29720 6722 29776
rect 6790 29720 6846 29776
rect 6914 29720 6970 29776
rect 7038 29720 7094 29776
rect 5178 29596 5234 29652
rect 5302 29596 5358 29652
rect 5426 29596 5482 29652
rect 5550 29596 5606 29652
rect 5674 29596 5730 29652
rect 5798 29596 5854 29652
rect 5922 29596 5978 29652
rect 6046 29596 6102 29652
rect 6170 29596 6226 29652
rect 6294 29596 6350 29652
rect 6418 29596 6474 29652
rect 6542 29596 6598 29652
rect 6666 29596 6722 29652
rect 6790 29596 6846 29652
rect 6914 29596 6970 29652
rect 7038 29596 7094 29652
rect 5178 29472 5234 29528
rect 5302 29472 5358 29528
rect 5426 29472 5482 29528
rect 5550 29472 5606 29528
rect 5674 29472 5730 29528
rect 5798 29472 5854 29528
rect 5922 29472 5978 29528
rect 6046 29472 6102 29528
rect 6170 29472 6226 29528
rect 6294 29472 6350 29528
rect 6418 29472 6474 29528
rect 6542 29472 6598 29528
rect 6666 29472 6722 29528
rect 6790 29472 6846 29528
rect 6914 29472 6970 29528
rect 7038 29472 7094 29528
rect 5178 29348 5234 29404
rect 5302 29348 5358 29404
rect 5426 29348 5482 29404
rect 5550 29348 5606 29404
rect 5674 29348 5730 29404
rect 5798 29348 5854 29404
rect 5922 29348 5978 29404
rect 6046 29348 6102 29404
rect 6170 29348 6226 29404
rect 6294 29348 6350 29404
rect 6418 29348 6474 29404
rect 6542 29348 6598 29404
rect 6666 29348 6722 29404
rect 6790 29348 6846 29404
rect 6914 29348 6970 29404
rect 7038 29348 7094 29404
rect 5178 29224 5234 29280
rect 5302 29224 5358 29280
rect 5426 29224 5482 29280
rect 5550 29224 5606 29280
rect 5674 29224 5730 29280
rect 5798 29224 5854 29280
rect 5922 29224 5978 29280
rect 6046 29224 6102 29280
rect 6170 29224 6226 29280
rect 6294 29224 6350 29280
rect 6418 29224 6474 29280
rect 6542 29224 6598 29280
rect 6666 29224 6722 29280
rect 6790 29224 6846 29280
rect 6914 29224 6970 29280
rect 7038 29224 7094 29280
rect 5178 29100 5234 29156
rect 5302 29100 5358 29156
rect 5426 29100 5482 29156
rect 5550 29100 5606 29156
rect 5674 29100 5730 29156
rect 5798 29100 5854 29156
rect 5922 29100 5978 29156
rect 6046 29100 6102 29156
rect 6170 29100 6226 29156
rect 6294 29100 6350 29156
rect 6418 29100 6474 29156
rect 6542 29100 6598 29156
rect 6666 29100 6722 29156
rect 6790 29100 6846 29156
rect 6914 29100 6970 29156
rect 7038 29100 7094 29156
rect 5178 28976 5234 29032
rect 5302 28976 5358 29032
rect 5426 28976 5482 29032
rect 5550 28976 5606 29032
rect 5674 28976 5730 29032
rect 5798 28976 5854 29032
rect 5922 28976 5978 29032
rect 6046 28976 6102 29032
rect 6170 28976 6226 29032
rect 6294 28976 6350 29032
rect 6418 28976 6474 29032
rect 6542 28976 6598 29032
rect 6666 28976 6722 29032
rect 6790 28976 6846 29032
rect 6914 28976 6970 29032
rect 7038 28976 7094 29032
rect 5178 28852 5234 28908
rect 5302 28852 5358 28908
rect 5426 28852 5482 28908
rect 5550 28852 5606 28908
rect 5674 28852 5730 28908
rect 5798 28852 5854 28908
rect 5922 28852 5978 28908
rect 6046 28852 6102 28908
rect 6170 28852 6226 28908
rect 6294 28852 6350 28908
rect 6418 28852 6474 28908
rect 6542 28852 6598 28908
rect 6666 28852 6722 28908
rect 6790 28852 6846 28908
rect 6914 28852 6970 28908
rect 7038 28852 7094 28908
rect 7884 30092 7940 30148
rect 8008 30092 8064 30148
rect 8132 30092 8188 30148
rect 8256 30092 8312 30148
rect 8380 30092 8436 30148
rect 8504 30092 8560 30148
rect 8628 30092 8684 30148
rect 8752 30092 8808 30148
rect 8876 30092 8932 30148
rect 9000 30092 9056 30148
rect 9124 30092 9180 30148
rect 9248 30092 9304 30148
rect 9372 30092 9428 30148
rect 9496 30092 9552 30148
rect 9620 30092 9676 30148
rect 9744 30092 9800 30148
rect 7884 29968 7940 30024
rect 8008 29968 8064 30024
rect 8132 29968 8188 30024
rect 8256 29968 8312 30024
rect 8380 29968 8436 30024
rect 8504 29968 8560 30024
rect 8628 29968 8684 30024
rect 8752 29968 8808 30024
rect 8876 29968 8932 30024
rect 9000 29968 9056 30024
rect 9124 29968 9180 30024
rect 9248 29968 9304 30024
rect 9372 29968 9428 30024
rect 9496 29968 9552 30024
rect 9620 29968 9676 30024
rect 9744 29968 9800 30024
rect 7884 29844 7940 29900
rect 8008 29844 8064 29900
rect 8132 29844 8188 29900
rect 8256 29844 8312 29900
rect 8380 29844 8436 29900
rect 8504 29844 8560 29900
rect 8628 29844 8684 29900
rect 8752 29844 8808 29900
rect 8876 29844 8932 29900
rect 9000 29844 9056 29900
rect 9124 29844 9180 29900
rect 9248 29844 9304 29900
rect 9372 29844 9428 29900
rect 9496 29844 9552 29900
rect 9620 29844 9676 29900
rect 9744 29844 9800 29900
rect 7884 29720 7940 29776
rect 8008 29720 8064 29776
rect 8132 29720 8188 29776
rect 8256 29720 8312 29776
rect 8380 29720 8436 29776
rect 8504 29720 8560 29776
rect 8628 29720 8684 29776
rect 8752 29720 8808 29776
rect 8876 29720 8932 29776
rect 9000 29720 9056 29776
rect 9124 29720 9180 29776
rect 9248 29720 9304 29776
rect 9372 29720 9428 29776
rect 9496 29720 9552 29776
rect 9620 29720 9676 29776
rect 9744 29720 9800 29776
rect 7884 29596 7940 29652
rect 8008 29596 8064 29652
rect 8132 29596 8188 29652
rect 8256 29596 8312 29652
rect 8380 29596 8436 29652
rect 8504 29596 8560 29652
rect 8628 29596 8684 29652
rect 8752 29596 8808 29652
rect 8876 29596 8932 29652
rect 9000 29596 9056 29652
rect 9124 29596 9180 29652
rect 9248 29596 9304 29652
rect 9372 29596 9428 29652
rect 9496 29596 9552 29652
rect 9620 29596 9676 29652
rect 9744 29596 9800 29652
rect 7884 29472 7940 29528
rect 8008 29472 8064 29528
rect 8132 29472 8188 29528
rect 8256 29472 8312 29528
rect 8380 29472 8436 29528
rect 8504 29472 8560 29528
rect 8628 29472 8684 29528
rect 8752 29472 8808 29528
rect 8876 29472 8932 29528
rect 9000 29472 9056 29528
rect 9124 29472 9180 29528
rect 9248 29472 9304 29528
rect 9372 29472 9428 29528
rect 9496 29472 9552 29528
rect 9620 29472 9676 29528
rect 9744 29472 9800 29528
rect 7884 29348 7940 29404
rect 8008 29348 8064 29404
rect 8132 29348 8188 29404
rect 8256 29348 8312 29404
rect 8380 29348 8436 29404
rect 8504 29348 8560 29404
rect 8628 29348 8684 29404
rect 8752 29348 8808 29404
rect 8876 29348 8932 29404
rect 9000 29348 9056 29404
rect 9124 29348 9180 29404
rect 9248 29348 9304 29404
rect 9372 29348 9428 29404
rect 9496 29348 9552 29404
rect 9620 29348 9676 29404
rect 9744 29348 9800 29404
rect 7884 29224 7940 29280
rect 8008 29224 8064 29280
rect 8132 29224 8188 29280
rect 8256 29224 8312 29280
rect 8380 29224 8436 29280
rect 8504 29224 8560 29280
rect 8628 29224 8684 29280
rect 8752 29224 8808 29280
rect 8876 29224 8932 29280
rect 9000 29224 9056 29280
rect 9124 29224 9180 29280
rect 9248 29224 9304 29280
rect 9372 29224 9428 29280
rect 9496 29224 9552 29280
rect 9620 29224 9676 29280
rect 9744 29224 9800 29280
rect 7884 29100 7940 29156
rect 8008 29100 8064 29156
rect 8132 29100 8188 29156
rect 8256 29100 8312 29156
rect 8380 29100 8436 29156
rect 8504 29100 8560 29156
rect 8628 29100 8684 29156
rect 8752 29100 8808 29156
rect 8876 29100 8932 29156
rect 9000 29100 9056 29156
rect 9124 29100 9180 29156
rect 9248 29100 9304 29156
rect 9372 29100 9428 29156
rect 9496 29100 9552 29156
rect 9620 29100 9676 29156
rect 9744 29100 9800 29156
rect 7884 28976 7940 29032
rect 8008 28976 8064 29032
rect 8132 28976 8188 29032
rect 8256 28976 8312 29032
rect 8380 28976 8436 29032
rect 8504 28976 8560 29032
rect 8628 28976 8684 29032
rect 8752 28976 8808 29032
rect 8876 28976 8932 29032
rect 9000 28976 9056 29032
rect 9124 28976 9180 29032
rect 9248 28976 9304 29032
rect 9372 28976 9428 29032
rect 9496 28976 9552 29032
rect 9620 28976 9676 29032
rect 9744 28976 9800 29032
rect 7884 28852 7940 28908
rect 8008 28852 8064 28908
rect 8132 28852 8188 28908
rect 8256 28852 8312 28908
rect 8380 28852 8436 28908
rect 8504 28852 8560 28908
rect 8628 28852 8684 28908
rect 8752 28852 8808 28908
rect 8876 28852 8932 28908
rect 9000 28852 9056 28908
rect 9124 28852 9180 28908
rect 9248 28852 9304 28908
rect 9372 28852 9428 28908
rect 9496 28852 9552 28908
rect 9620 28852 9676 28908
rect 9744 28852 9800 28908
rect 10254 30092 10310 30148
rect 10378 30092 10434 30148
rect 10502 30092 10558 30148
rect 10626 30092 10682 30148
rect 10750 30092 10806 30148
rect 10874 30092 10930 30148
rect 10998 30092 11054 30148
rect 11122 30092 11178 30148
rect 11246 30092 11302 30148
rect 11370 30092 11426 30148
rect 11494 30092 11550 30148
rect 11618 30092 11674 30148
rect 11742 30092 11798 30148
rect 11866 30092 11922 30148
rect 11990 30092 12046 30148
rect 12114 30092 12170 30148
rect 10254 29968 10310 30024
rect 10378 29968 10434 30024
rect 10502 29968 10558 30024
rect 10626 29968 10682 30024
rect 10750 29968 10806 30024
rect 10874 29968 10930 30024
rect 10998 29968 11054 30024
rect 11122 29968 11178 30024
rect 11246 29968 11302 30024
rect 11370 29968 11426 30024
rect 11494 29968 11550 30024
rect 11618 29968 11674 30024
rect 11742 29968 11798 30024
rect 11866 29968 11922 30024
rect 11990 29968 12046 30024
rect 12114 29968 12170 30024
rect 10254 29844 10310 29900
rect 10378 29844 10434 29900
rect 10502 29844 10558 29900
rect 10626 29844 10682 29900
rect 10750 29844 10806 29900
rect 10874 29844 10930 29900
rect 10998 29844 11054 29900
rect 11122 29844 11178 29900
rect 11246 29844 11302 29900
rect 11370 29844 11426 29900
rect 11494 29844 11550 29900
rect 11618 29844 11674 29900
rect 11742 29844 11798 29900
rect 11866 29844 11922 29900
rect 11990 29844 12046 29900
rect 12114 29844 12170 29900
rect 10254 29720 10310 29776
rect 10378 29720 10434 29776
rect 10502 29720 10558 29776
rect 10626 29720 10682 29776
rect 10750 29720 10806 29776
rect 10874 29720 10930 29776
rect 10998 29720 11054 29776
rect 11122 29720 11178 29776
rect 11246 29720 11302 29776
rect 11370 29720 11426 29776
rect 11494 29720 11550 29776
rect 11618 29720 11674 29776
rect 11742 29720 11798 29776
rect 11866 29720 11922 29776
rect 11990 29720 12046 29776
rect 12114 29720 12170 29776
rect 10254 29596 10310 29652
rect 10378 29596 10434 29652
rect 10502 29596 10558 29652
rect 10626 29596 10682 29652
rect 10750 29596 10806 29652
rect 10874 29596 10930 29652
rect 10998 29596 11054 29652
rect 11122 29596 11178 29652
rect 11246 29596 11302 29652
rect 11370 29596 11426 29652
rect 11494 29596 11550 29652
rect 11618 29596 11674 29652
rect 11742 29596 11798 29652
rect 11866 29596 11922 29652
rect 11990 29596 12046 29652
rect 12114 29596 12170 29652
rect 10254 29472 10310 29528
rect 10378 29472 10434 29528
rect 10502 29472 10558 29528
rect 10626 29472 10682 29528
rect 10750 29472 10806 29528
rect 10874 29472 10930 29528
rect 10998 29472 11054 29528
rect 11122 29472 11178 29528
rect 11246 29472 11302 29528
rect 11370 29472 11426 29528
rect 11494 29472 11550 29528
rect 11618 29472 11674 29528
rect 11742 29472 11798 29528
rect 11866 29472 11922 29528
rect 11990 29472 12046 29528
rect 12114 29472 12170 29528
rect 10254 29348 10310 29404
rect 10378 29348 10434 29404
rect 10502 29348 10558 29404
rect 10626 29348 10682 29404
rect 10750 29348 10806 29404
rect 10874 29348 10930 29404
rect 10998 29348 11054 29404
rect 11122 29348 11178 29404
rect 11246 29348 11302 29404
rect 11370 29348 11426 29404
rect 11494 29348 11550 29404
rect 11618 29348 11674 29404
rect 11742 29348 11798 29404
rect 11866 29348 11922 29404
rect 11990 29348 12046 29404
rect 12114 29348 12170 29404
rect 10254 29224 10310 29280
rect 10378 29224 10434 29280
rect 10502 29224 10558 29280
rect 10626 29224 10682 29280
rect 10750 29224 10806 29280
rect 10874 29224 10930 29280
rect 10998 29224 11054 29280
rect 11122 29224 11178 29280
rect 11246 29224 11302 29280
rect 11370 29224 11426 29280
rect 11494 29224 11550 29280
rect 11618 29224 11674 29280
rect 11742 29224 11798 29280
rect 11866 29224 11922 29280
rect 11990 29224 12046 29280
rect 12114 29224 12170 29280
rect 10254 29100 10310 29156
rect 10378 29100 10434 29156
rect 10502 29100 10558 29156
rect 10626 29100 10682 29156
rect 10750 29100 10806 29156
rect 10874 29100 10930 29156
rect 10998 29100 11054 29156
rect 11122 29100 11178 29156
rect 11246 29100 11302 29156
rect 11370 29100 11426 29156
rect 11494 29100 11550 29156
rect 11618 29100 11674 29156
rect 11742 29100 11798 29156
rect 11866 29100 11922 29156
rect 11990 29100 12046 29156
rect 12114 29100 12170 29156
rect 10254 28976 10310 29032
rect 10378 28976 10434 29032
rect 10502 28976 10558 29032
rect 10626 28976 10682 29032
rect 10750 28976 10806 29032
rect 10874 28976 10930 29032
rect 10998 28976 11054 29032
rect 11122 28976 11178 29032
rect 11246 28976 11302 29032
rect 11370 28976 11426 29032
rect 11494 28976 11550 29032
rect 11618 28976 11674 29032
rect 11742 28976 11798 29032
rect 11866 28976 11922 29032
rect 11990 28976 12046 29032
rect 12114 28976 12170 29032
rect 10254 28852 10310 28908
rect 10378 28852 10434 28908
rect 10502 28852 10558 28908
rect 10626 28852 10682 28908
rect 10750 28852 10806 28908
rect 10874 28852 10930 28908
rect 10998 28852 11054 28908
rect 11122 28852 11178 28908
rect 11246 28852 11302 28908
rect 11370 28852 11426 28908
rect 11494 28852 11550 28908
rect 11618 28852 11674 28908
rect 11742 28852 11798 28908
rect 11866 28852 11922 28908
rect 11990 28852 12046 28908
rect 12114 28852 12170 28908
rect 12871 30092 12927 30148
rect 12995 30092 13051 30148
rect 13119 30092 13175 30148
rect 13243 30092 13299 30148
rect 13367 30092 13423 30148
rect 13491 30092 13547 30148
rect 13615 30092 13671 30148
rect 13739 30092 13795 30148
rect 13863 30092 13919 30148
rect 13987 30092 14043 30148
rect 14111 30092 14167 30148
rect 14235 30092 14291 30148
rect 14359 30092 14415 30148
rect 14483 30092 14539 30148
rect 14607 30092 14663 30148
rect 12871 29968 12927 30024
rect 12995 29968 13051 30024
rect 13119 29968 13175 30024
rect 13243 29968 13299 30024
rect 13367 29968 13423 30024
rect 13491 29968 13547 30024
rect 13615 29968 13671 30024
rect 13739 29968 13795 30024
rect 13863 29968 13919 30024
rect 13987 29968 14043 30024
rect 14111 29968 14167 30024
rect 14235 29968 14291 30024
rect 14359 29968 14415 30024
rect 14483 29968 14539 30024
rect 14607 29968 14663 30024
rect 12871 29844 12927 29900
rect 12995 29844 13051 29900
rect 13119 29844 13175 29900
rect 13243 29844 13299 29900
rect 13367 29844 13423 29900
rect 13491 29844 13547 29900
rect 13615 29844 13671 29900
rect 13739 29844 13795 29900
rect 13863 29844 13919 29900
rect 13987 29844 14043 29900
rect 14111 29844 14167 29900
rect 14235 29844 14291 29900
rect 14359 29844 14415 29900
rect 14483 29844 14539 29900
rect 14607 29844 14663 29900
rect 12871 29720 12927 29776
rect 12995 29720 13051 29776
rect 13119 29720 13175 29776
rect 13243 29720 13299 29776
rect 13367 29720 13423 29776
rect 13491 29720 13547 29776
rect 13615 29720 13671 29776
rect 13739 29720 13795 29776
rect 13863 29720 13919 29776
rect 13987 29720 14043 29776
rect 14111 29720 14167 29776
rect 14235 29720 14291 29776
rect 14359 29720 14415 29776
rect 14483 29720 14539 29776
rect 14607 29720 14663 29776
rect 12871 29596 12927 29652
rect 12995 29596 13051 29652
rect 13119 29596 13175 29652
rect 13243 29596 13299 29652
rect 13367 29596 13423 29652
rect 13491 29596 13547 29652
rect 13615 29596 13671 29652
rect 13739 29596 13795 29652
rect 13863 29596 13919 29652
rect 13987 29596 14043 29652
rect 14111 29596 14167 29652
rect 14235 29596 14291 29652
rect 14359 29596 14415 29652
rect 14483 29596 14539 29652
rect 14607 29596 14663 29652
rect 12871 29472 12927 29528
rect 12995 29472 13051 29528
rect 13119 29472 13175 29528
rect 13243 29472 13299 29528
rect 13367 29472 13423 29528
rect 13491 29472 13547 29528
rect 13615 29472 13671 29528
rect 13739 29472 13795 29528
rect 13863 29472 13919 29528
rect 13987 29472 14043 29528
rect 14111 29472 14167 29528
rect 14235 29472 14291 29528
rect 14359 29472 14415 29528
rect 14483 29472 14539 29528
rect 14607 29472 14663 29528
rect 12871 29348 12927 29404
rect 12995 29348 13051 29404
rect 13119 29348 13175 29404
rect 13243 29348 13299 29404
rect 13367 29348 13423 29404
rect 13491 29348 13547 29404
rect 13615 29348 13671 29404
rect 13739 29348 13795 29404
rect 13863 29348 13919 29404
rect 13987 29348 14043 29404
rect 14111 29348 14167 29404
rect 14235 29348 14291 29404
rect 14359 29348 14415 29404
rect 14483 29348 14539 29404
rect 14607 29348 14663 29404
rect 12871 29224 12927 29280
rect 12995 29224 13051 29280
rect 13119 29224 13175 29280
rect 13243 29224 13299 29280
rect 13367 29224 13423 29280
rect 13491 29224 13547 29280
rect 13615 29224 13671 29280
rect 13739 29224 13795 29280
rect 13863 29224 13919 29280
rect 13987 29224 14043 29280
rect 14111 29224 14167 29280
rect 14235 29224 14291 29280
rect 14359 29224 14415 29280
rect 14483 29224 14539 29280
rect 14607 29224 14663 29280
rect 12871 29100 12927 29156
rect 12995 29100 13051 29156
rect 13119 29100 13175 29156
rect 13243 29100 13299 29156
rect 13367 29100 13423 29156
rect 13491 29100 13547 29156
rect 13615 29100 13671 29156
rect 13739 29100 13795 29156
rect 13863 29100 13919 29156
rect 13987 29100 14043 29156
rect 14111 29100 14167 29156
rect 14235 29100 14291 29156
rect 14359 29100 14415 29156
rect 14483 29100 14539 29156
rect 14607 29100 14663 29156
rect 12871 28976 12927 29032
rect 12995 28976 13051 29032
rect 13119 28976 13175 29032
rect 13243 28976 13299 29032
rect 13367 28976 13423 29032
rect 13491 28976 13547 29032
rect 13615 28976 13671 29032
rect 13739 28976 13795 29032
rect 13863 28976 13919 29032
rect 13987 28976 14043 29032
rect 14111 28976 14167 29032
rect 14235 28976 14291 29032
rect 14359 28976 14415 29032
rect 14483 28976 14539 29032
rect 14607 28976 14663 29032
rect 12871 28852 12927 28908
rect 12995 28852 13051 28908
rect 13119 28852 13175 28908
rect 13243 28852 13299 28908
rect 13367 28852 13423 28908
rect 13491 28852 13547 28908
rect 13615 28852 13671 28908
rect 13739 28852 13795 28908
rect 13863 28852 13919 28908
rect 13987 28852 14043 28908
rect 14111 28852 14167 28908
rect 14235 28852 14291 28908
rect 14359 28852 14415 28908
rect 14483 28852 14539 28908
rect 14607 28852 14663 28908
rect 2491 28492 2547 28548
rect 2615 28492 2671 28548
rect 2491 28368 2547 28424
rect 2615 28368 2671 28424
rect 2491 28244 2547 28300
rect 2615 28244 2671 28300
rect 2491 28120 2547 28176
rect 2615 28120 2671 28176
rect 2491 27996 2547 28052
rect 2615 27996 2671 28052
rect 2491 27872 2547 27928
rect 2615 27872 2671 27928
rect 2491 27748 2547 27804
rect 2615 27748 2671 27804
rect 2491 27624 2547 27680
rect 2615 27624 2671 27680
rect 2491 27500 2547 27556
rect 2615 27500 2671 27556
rect 2491 27376 2547 27432
rect 2615 27376 2671 27432
rect 2491 27252 2547 27308
rect 2615 27252 2671 27308
rect 4861 28492 4917 28548
rect 4985 28492 5041 28548
rect 4861 28368 4917 28424
rect 4985 28368 5041 28424
rect 4861 28244 4917 28300
rect 4985 28244 5041 28300
rect 4861 28120 4917 28176
rect 4985 28120 5041 28176
rect 4861 27996 4917 28052
rect 4985 27996 5041 28052
rect 4861 27872 4917 27928
rect 4985 27872 5041 27928
rect 4861 27748 4917 27804
rect 4985 27748 5041 27804
rect 4861 27624 4917 27680
rect 4985 27624 5041 27680
rect 4861 27500 4917 27556
rect 4985 27500 5041 27556
rect 4861 27376 4917 27432
rect 4985 27376 5041 27432
rect 4861 27252 4917 27308
rect 4985 27252 5041 27308
rect 7275 28492 7331 28548
rect 7399 28492 7455 28548
rect 7523 28492 7579 28548
rect 7647 28492 7703 28548
rect 7275 28368 7331 28424
rect 7399 28368 7455 28424
rect 7523 28368 7579 28424
rect 7647 28368 7703 28424
rect 7275 28244 7331 28300
rect 7399 28244 7455 28300
rect 7523 28244 7579 28300
rect 7647 28244 7703 28300
rect 7275 28120 7331 28176
rect 7399 28120 7455 28176
rect 7523 28120 7579 28176
rect 7647 28120 7703 28176
rect 7275 27996 7331 28052
rect 7399 27996 7455 28052
rect 7523 27996 7579 28052
rect 7647 27996 7703 28052
rect 7275 27872 7331 27928
rect 7399 27872 7455 27928
rect 7523 27872 7579 27928
rect 7647 27872 7703 27928
rect 7275 27748 7331 27804
rect 7399 27748 7455 27804
rect 7523 27748 7579 27804
rect 7647 27748 7703 27804
rect 7275 27624 7331 27680
rect 7399 27624 7455 27680
rect 7523 27624 7579 27680
rect 7647 27624 7703 27680
rect 7275 27500 7331 27556
rect 7399 27500 7455 27556
rect 7523 27500 7579 27556
rect 7647 27500 7703 27556
rect 7275 27376 7331 27432
rect 7399 27376 7455 27432
rect 7523 27376 7579 27432
rect 7647 27376 7703 27432
rect 7275 27252 7331 27308
rect 7399 27252 7455 27308
rect 7523 27252 7579 27308
rect 7647 27252 7703 27308
rect 9937 28492 9993 28548
rect 10061 28492 10117 28548
rect 9937 28368 9993 28424
rect 10061 28368 10117 28424
rect 9937 28244 9993 28300
rect 10061 28244 10117 28300
rect 9937 28120 9993 28176
rect 10061 28120 10117 28176
rect 9937 27996 9993 28052
rect 10061 27996 10117 28052
rect 9937 27872 9993 27928
rect 10061 27872 10117 27928
rect 9937 27748 9993 27804
rect 10061 27748 10117 27804
rect 9937 27624 9993 27680
rect 10061 27624 10117 27680
rect 9937 27500 9993 27556
rect 10061 27500 10117 27556
rect 9937 27376 9993 27432
rect 10061 27376 10117 27432
rect 9937 27252 9993 27308
rect 10061 27252 10117 27308
rect 12307 28492 12363 28548
rect 12431 28492 12487 28548
rect 12307 28368 12363 28424
rect 12431 28368 12487 28424
rect 12307 28244 12363 28300
rect 12431 28244 12487 28300
rect 12307 28120 12363 28176
rect 12431 28120 12487 28176
rect 12307 27996 12363 28052
rect 12431 27996 12487 28052
rect 12307 27872 12363 27928
rect 12431 27872 12487 27928
rect 12307 27748 12363 27804
rect 12431 27748 12487 27804
rect 12307 27624 12363 27680
rect 12431 27624 12487 27680
rect 12307 27500 12363 27556
rect 12431 27500 12487 27556
rect 12307 27376 12363 27432
rect 12431 27376 12487 27432
rect 12307 27252 12363 27308
rect 12431 27252 12487 27308
rect 315 26898 371 26954
rect 439 26898 495 26954
rect 563 26898 619 26954
rect 687 26898 743 26954
rect 811 26898 867 26954
rect 935 26898 991 26954
rect 1059 26898 1115 26954
rect 1183 26898 1239 26954
rect 1307 26898 1363 26954
rect 1431 26898 1487 26954
rect 1555 26898 1611 26954
rect 1679 26898 1735 26954
rect 1803 26898 1859 26954
rect 1927 26898 1983 26954
rect 2051 26898 2107 26954
rect 315 26774 371 26830
rect 439 26774 495 26830
rect 563 26774 619 26830
rect 687 26774 743 26830
rect 811 26774 867 26830
rect 935 26774 991 26830
rect 1059 26774 1115 26830
rect 1183 26774 1239 26830
rect 1307 26774 1363 26830
rect 1431 26774 1487 26830
rect 1555 26774 1611 26830
rect 1679 26774 1735 26830
rect 1803 26774 1859 26830
rect 1927 26774 1983 26830
rect 2051 26774 2107 26830
rect 315 26650 371 26706
rect 439 26650 495 26706
rect 563 26650 619 26706
rect 687 26650 743 26706
rect 811 26650 867 26706
rect 935 26650 991 26706
rect 1059 26650 1115 26706
rect 1183 26650 1239 26706
rect 1307 26650 1363 26706
rect 1431 26650 1487 26706
rect 1555 26650 1611 26706
rect 1679 26650 1735 26706
rect 1803 26650 1859 26706
rect 1927 26650 1983 26706
rect 2051 26650 2107 26706
rect 315 26526 371 26582
rect 439 26526 495 26582
rect 563 26526 619 26582
rect 687 26526 743 26582
rect 811 26526 867 26582
rect 935 26526 991 26582
rect 1059 26526 1115 26582
rect 1183 26526 1239 26582
rect 1307 26526 1363 26582
rect 1431 26526 1487 26582
rect 1555 26526 1611 26582
rect 1679 26526 1735 26582
rect 1803 26526 1859 26582
rect 1927 26526 1983 26582
rect 2051 26526 2107 26582
rect 315 26402 371 26458
rect 439 26402 495 26458
rect 563 26402 619 26458
rect 687 26402 743 26458
rect 811 26402 867 26458
rect 935 26402 991 26458
rect 1059 26402 1115 26458
rect 1183 26402 1239 26458
rect 1307 26402 1363 26458
rect 1431 26402 1487 26458
rect 1555 26402 1611 26458
rect 1679 26402 1735 26458
rect 1803 26402 1859 26458
rect 1927 26402 1983 26458
rect 2051 26402 2107 26458
rect 315 26278 371 26334
rect 439 26278 495 26334
rect 563 26278 619 26334
rect 687 26278 743 26334
rect 811 26278 867 26334
rect 935 26278 991 26334
rect 1059 26278 1115 26334
rect 1183 26278 1239 26334
rect 1307 26278 1363 26334
rect 1431 26278 1487 26334
rect 1555 26278 1611 26334
rect 1679 26278 1735 26334
rect 1803 26278 1859 26334
rect 1927 26278 1983 26334
rect 2051 26278 2107 26334
rect 315 26154 371 26210
rect 439 26154 495 26210
rect 563 26154 619 26210
rect 687 26154 743 26210
rect 811 26154 867 26210
rect 935 26154 991 26210
rect 1059 26154 1115 26210
rect 1183 26154 1239 26210
rect 1307 26154 1363 26210
rect 1431 26154 1487 26210
rect 1555 26154 1611 26210
rect 1679 26154 1735 26210
rect 1803 26154 1859 26210
rect 1927 26154 1983 26210
rect 2051 26154 2107 26210
rect 315 26030 371 26086
rect 439 26030 495 26086
rect 563 26030 619 26086
rect 687 26030 743 26086
rect 811 26030 867 26086
rect 935 26030 991 26086
rect 1059 26030 1115 26086
rect 1183 26030 1239 26086
rect 1307 26030 1363 26086
rect 1431 26030 1487 26086
rect 1555 26030 1611 26086
rect 1679 26030 1735 26086
rect 1803 26030 1859 26086
rect 1927 26030 1983 26086
rect 2051 26030 2107 26086
rect 315 25906 371 25962
rect 439 25906 495 25962
rect 563 25906 619 25962
rect 687 25906 743 25962
rect 811 25906 867 25962
rect 935 25906 991 25962
rect 1059 25906 1115 25962
rect 1183 25906 1239 25962
rect 1307 25906 1363 25962
rect 1431 25906 1487 25962
rect 1555 25906 1611 25962
rect 1679 25906 1735 25962
rect 1803 25906 1859 25962
rect 1927 25906 1983 25962
rect 2051 25906 2107 25962
rect 315 25782 371 25838
rect 439 25782 495 25838
rect 563 25782 619 25838
rect 687 25782 743 25838
rect 811 25782 867 25838
rect 935 25782 991 25838
rect 1059 25782 1115 25838
rect 1183 25782 1239 25838
rect 1307 25782 1363 25838
rect 1431 25782 1487 25838
rect 1555 25782 1611 25838
rect 1679 25782 1735 25838
rect 1803 25782 1859 25838
rect 1927 25782 1983 25838
rect 2051 25782 2107 25838
rect 315 25658 371 25714
rect 439 25658 495 25714
rect 563 25658 619 25714
rect 687 25658 743 25714
rect 811 25658 867 25714
rect 935 25658 991 25714
rect 1059 25658 1115 25714
rect 1183 25658 1239 25714
rect 1307 25658 1363 25714
rect 1431 25658 1487 25714
rect 1555 25658 1611 25714
rect 1679 25658 1735 25714
rect 1803 25658 1859 25714
rect 1927 25658 1983 25714
rect 2051 25658 2107 25714
rect 315 25534 371 25590
rect 439 25534 495 25590
rect 563 25534 619 25590
rect 687 25534 743 25590
rect 811 25534 867 25590
rect 935 25534 991 25590
rect 1059 25534 1115 25590
rect 1183 25534 1239 25590
rect 1307 25534 1363 25590
rect 1431 25534 1487 25590
rect 1555 25534 1611 25590
rect 1679 25534 1735 25590
rect 1803 25534 1859 25590
rect 1927 25534 1983 25590
rect 2051 25534 2107 25590
rect 315 25410 371 25466
rect 439 25410 495 25466
rect 563 25410 619 25466
rect 687 25410 743 25466
rect 811 25410 867 25466
rect 935 25410 991 25466
rect 1059 25410 1115 25466
rect 1183 25410 1239 25466
rect 1307 25410 1363 25466
rect 1431 25410 1487 25466
rect 1555 25410 1611 25466
rect 1679 25410 1735 25466
rect 1803 25410 1859 25466
rect 1927 25410 1983 25466
rect 2051 25410 2107 25466
rect 315 25286 371 25342
rect 439 25286 495 25342
rect 563 25286 619 25342
rect 687 25286 743 25342
rect 811 25286 867 25342
rect 935 25286 991 25342
rect 1059 25286 1115 25342
rect 1183 25286 1239 25342
rect 1307 25286 1363 25342
rect 1431 25286 1487 25342
rect 1555 25286 1611 25342
rect 1679 25286 1735 25342
rect 1803 25286 1859 25342
rect 1927 25286 1983 25342
rect 2051 25286 2107 25342
rect 315 25162 371 25218
rect 439 25162 495 25218
rect 563 25162 619 25218
rect 687 25162 743 25218
rect 811 25162 867 25218
rect 935 25162 991 25218
rect 1059 25162 1115 25218
rect 1183 25162 1239 25218
rect 1307 25162 1363 25218
rect 1431 25162 1487 25218
rect 1555 25162 1611 25218
rect 1679 25162 1735 25218
rect 1803 25162 1859 25218
rect 1927 25162 1983 25218
rect 2051 25162 2107 25218
rect 315 25038 371 25094
rect 439 25038 495 25094
rect 563 25038 619 25094
rect 687 25038 743 25094
rect 811 25038 867 25094
rect 935 25038 991 25094
rect 1059 25038 1115 25094
rect 1183 25038 1239 25094
rect 1307 25038 1363 25094
rect 1431 25038 1487 25094
rect 1555 25038 1611 25094
rect 1679 25038 1735 25094
rect 1803 25038 1859 25094
rect 1927 25038 1983 25094
rect 2051 25038 2107 25094
rect 315 24914 371 24970
rect 439 24914 495 24970
rect 563 24914 619 24970
rect 687 24914 743 24970
rect 811 24914 867 24970
rect 935 24914 991 24970
rect 1059 24914 1115 24970
rect 1183 24914 1239 24970
rect 1307 24914 1363 24970
rect 1431 24914 1487 24970
rect 1555 24914 1611 24970
rect 1679 24914 1735 24970
rect 1803 24914 1859 24970
rect 1927 24914 1983 24970
rect 2051 24914 2107 24970
rect 315 24790 371 24846
rect 439 24790 495 24846
rect 563 24790 619 24846
rect 687 24790 743 24846
rect 811 24790 867 24846
rect 935 24790 991 24846
rect 1059 24790 1115 24846
rect 1183 24790 1239 24846
rect 1307 24790 1363 24846
rect 1431 24790 1487 24846
rect 1555 24790 1611 24846
rect 1679 24790 1735 24846
rect 1803 24790 1859 24846
rect 1927 24790 1983 24846
rect 2051 24790 2107 24846
rect 315 24666 371 24722
rect 439 24666 495 24722
rect 563 24666 619 24722
rect 687 24666 743 24722
rect 811 24666 867 24722
rect 935 24666 991 24722
rect 1059 24666 1115 24722
rect 1183 24666 1239 24722
rect 1307 24666 1363 24722
rect 1431 24666 1487 24722
rect 1555 24666 1611 24722
rect 1679 24666 1735 24722
rect 1803 24666 1859 24722
rect 1927 24666 1983 24722
rect 2051 24666 2107 24722
rect 315 24542 371 24598
rect 439 24542 495 24598
rect 563 24542 619 24598
rect 687 24542 743 24598
rect 811 24542 867 24598
rect 935 24542 991 24598
rect 1059 24542 1115 24598
rect 1183 24542 1239 24598
rect 1307 24542 1363 24598
rect 1431 24542 1487 24598
rect 1555 24542 1611 24598
rect 1679 24542 1735 24598
rect 1803 24542 1859 24598
rect 1927 24542 1983 24598
rect 2051 24542 2107 24598
rect 315 24418 371 24474
rect 439 24418 495 24474
rect 563 24418 619 24474
rect 687 24418 743 24474
rect 811 24418 867 24474
rect 935 24418 991 24474
rect 1059 24418 1115 24474
rect 1183 24418 1239 24474
rect 1307 24418 1363 24474
rect 1431 24418 1487 24474
rect 1555 24418 1611 24474
rect 1679 24418 1735 24474
rect 1803 24418 1859 24474
rect 1927 24418 1983 24474
rect 2051 24418 2107 24474
rect 315 24294 371 24350
rect 439 24294 495 24350
rect 563 24294 619 24350
rect 687 24294 743 24350
rect 811 24294 867 24350
rect 935 24294 991 24350
rect 1059 24294 1115 24350
rect 1183 24294 1239 24350
rect 1307 24294 1363 24350
rect 1431 24294 1487 24350
rect 1555 24294 1611 24350
rect 1679 24294 1735 24350
rect 1803 24294 1859 24350
rect 1927 24294 1983 24350
rect 2051 24294 2107 24350
rect 315 24170 371 24226
rect 439 24170 495 24226
rect 563 24170 619 24226
rect 687 24170 743 24226
rect 811 24170 867 24226
rect 935 24170 991 24226
rect 1059 24170 1115 24226
rect 1183 24170 1239 24226
rect 1307 24170 1363 24226
rect 1431 24170 1487 24226
rect 1555 24170 1611 24226
rect 1679 24170 1735 24226
rect 1803 24170 1859 24226
rect 1927 24170 1983 24226
rect 2051 24170 2107 24226
rect 315 24046 371 24102
rect 439 24046 495 24102
rect 563 24046 619 24102
rect 687 24046 743 24102
rect 811 24046 867 24102
rect 935 24046 991 24102
rect 1059 24046 1115 24102
rect 1183 24046 1239 24102
rect 1307 24046 1363 24102
rect 1431 24046 1487 24102
rect 1555 24046 1611 24102
rect 1679 24046 1735 24102
rect 1803 24046 1859 24102
rect 1927 24046 1983 24102
rect 2051 24046 2107 24102
rect 2808 26898 2864 26954
rect 2932 26898 2988 26954
rect 3056 26898 3112 26954
rect 3180 26898 3236 26954
rect 3304 26898 3360 26954
rect 3428 26898 3484 26954
rect 3552 26898 3608 26954
rect 3676 26898 3732 26954
rect 3800 26898 3856 26954
rect 3924 26898 3980 26954
rect 4048 26898 4104 26954
rect 4172 26898 4228 26954
rect 4296 26898 4352 26954
rect 4420 26898 4476 26954
rect 4544 26898 4600 26954
rect 4668 26898 4724 26954
rect 2808 26774 2864 26830
rect 2932 26774 2988 26830
rect 3056 26774 3112 26830
rect 3180 26774 3236 26830
rect 3304 26774 3360 26830
rect 3428 26774 3484 26830
rect 3552 26774 3608 26830
rect 3676 26774 3732 26830
rect 3800 26774 3856 26830
rect 3924 26774 3980 26830
rect 4048 26774 4104 26830
rect 4172 26774 4228 26830
rect 4296 26774 4352 26830
rect 4420 26774 4476 26830
rect 4544 26774 4600 26830
rect 4668 26774 4724 26830
rect 2808 26650 2864 26706
rect 2932 26650 2988 26706
rect 3056 26650 3112 26706
rect 3180 26650 3236 26706
rect 3304 26650 3360 26706
rect 3428 26650 3484 26706
rect 3552 26650 3608 26706
rect 3676 26650 3732 26706
rect 3800 26650 3856 26706
rect 3924 26650 3980 26706
rect 4048 26650 4104 26706
rect 4172 26650 4228 26706
rect 4296 26650 4352 26706
rect 4420 26650 4476 26706
rect 4544 26650 4600 26706
rect 4668 26650 4724 26706
rect 2808 26526 2864 26582
rect 2932 26526 2988 26582
rect 3056 26526 3112 26582
rect 3180 26526 3236 26582
rect 3304 26526 3360 26582
rect 3428 26526 3484 26582
rect 3552 26526 3608 26582
rect 3676 26526 3732 26582
rect 3800 26526 3856 26582
rect 3924 26526 3980 26582
rect 4048 26526 4104 26582
rect 4172 26526 4228 26582
rect 4296 26526 4352 26582
rect 4420 26526 4476 26582
rect 4544 26526 4600 26582
rect 4668 26526 4724 26582
rect 2808 26402 2864 26458
rect 2932 26402 2988 26458
rect 3056 26402 3112 26458
rect 3180 26402 3236 26458
rect 3304 26402 3360 26458
rect 3428 26402 3484 26458
rect 3552 26402 3608 26458
rect 3676 26402 3732 26458
rect 3800 26402 3856 26458
rect 3924 26402 3980 26458
rect 4048 26402 4104 26458
rect 4172 26402 4228 26458
rect 4296 26402 4352 26458
rect 4420 26402 4476 26458
rect 4544 26402 4600 26458
rect 4668 26402 4724 26458
rect 2808 26278 2864 26334
rect 2932 26278 2988 26334
rect 3056 26278 3112 26334
rect 3180 26278 3236 26334
rect 3304 26278 3360 26334
rect 3428 26278 3484 26334
rect 3552 26278 3608 26334
rect 3676 26278 3732 26334
rect 3800 26278 3856 26334
rect 3924 26278 3980 26334
rect 4048 26278 4104 26334
rect 4172 26278 4228 26334
rect 4296 26278 4352 26334
rect 4420 26278 4476 26334
rect 4544 26278 4600 26334
rect 4668 26278 4724 26334
rect 2808 26154 2864 26210
rect 2932 26154 2988 26210
rect 3056 26154 3112 26210
rect 3180 26154 3236 26210
rect 3304 26154 3360 26210
rect 3428 26154 3484 26210
rect 3552 26154 3608 26210
rect 3676 26154 3732 26210
rect 3800 26154 3856 26210
rect 3924 26154 3980 26210
rect 4048 26154 4104 26210
rect 4172 26154 4228 26210
rect 4296 26154 4352 26210
rect 4420 26154 4476 26210
rect 4544 26154 4600 26210
rect 4668 26154 4724 26210
rect 2808 26030 2864 26086
rect 2932 26030 2988 26086
rect 3056 26030 3112 26086
rect 3180 26030 3236 26086
rect 3304 26030 3360 26086
rect 3428 26030 3484 26086
rect 3552 26030 3608 26086
rect 3676 26030 3732 26086
rect 3800 26030 3856 26086
rect 3924 26030 3980 26086
rect 4048 26030 4104 26086
rect 4172 26030 4228 26086
rect 4296 26030 4352 26086
rect 4420 26030 4476 26086
rect 4544 26030 4600 26086
rect 4668 26030 4724 26086
rect 2808 25906 2864 25962
rect 2932 25906 2988 25962
rect 3056 25906 3112 25962
rect 3180 25906 3236 25962
rect 3304 25906 3360 25962
rect 3428 25906 3484 25962
rect 3552 25906 3608 25962
rect 3676 25906 3732 25962
rect 3800 25906 3856 25962
rect 3924 25906 3980 25962
rect 4048 25906 4104 25962
rect 4172 25906 4228 25962
rect 4296 25906 4352 25962
rect 4420 25906 4476 25962
rect 4544 25906 4600 25962
rect 4668 25906 4724 25962
rect 2808 25782 2864 25838
rect 2932 25782 2988 25838
rect 3056 25782 3112 25838
rect 3180 25782 3236 25838
rect 3304 25782 3360 25838
rect 3428 25782 3484 25838
rect 3552 25782 3608 25838
rect 3676 25782 3732 25838
rect 3800 25782 3856 25838
rect 3924 25782 3980 25838
rect 4048 25782 4104 25838
rect 4172 25782 4228 25838
rect 4296 25782 4352 25838
rect 4420 25782 4476 25838
rect 4544 25782 4600 25838
rect 4668 25782 4724 25838
rect 2808 25658 2864 25714
rect 2932 25658 2988 25714
rect 3056 25658 3112 25714
rect 3180 25658 3236 25714
rect 3304 25658 3360 25714
rect 3428 25658 3484 25714
rect 3552 25658 3608 25714
rect 3676 25658 3732 25714
rect 3800 25658 3856 25714
rect 3924 25658 3980 25714
rect 4048 25658 4104 25714
rect 4172 25658 4228 25714
rect 4296 25658 4352 25714
rect 4420 25658 4476 25714
rect 4544 25658 4600 25714
rect 4668 25658 4724 25714
rect 2808 25534 2864 25590
rect 2932 25534 2988 25590
rect 3056 25534 3112 25590
rect 3180 25534 3236 25590
rect 3304 25534 3360 25590
rect 3428 25534 3484 25590
rect 3552 25534 3608 25590
rect 3676 25534 3732 25590
rect 3800 25534 3856 25590
rect 3924 25534 3980 25590
rect 4048 25534 4104 25590
rect 4172 25534 4228 25590
rect 4296 25534 4352 25590
rect 4420 25534 4476 25590
rect 4544 25534 4600 25590
rect 4668 25534 4724 25590
rect 2808 25410 2864 25466
rect 2932 25410 2988 25466
rect 3056 25410 3112 25466
rect 3180 25410 3236 25466
rect 3304 25410 3360 25466
rect 3428 25410 3484 25466
rect 3552 25410 3608 25466
rect 3676 25410 3732 25466
rect 3800 25410 3856 25466
rect 3924 25410 3980 25466
rect 4048 25410 4104 25466
rect 4172 25410 4228 25466
rect 4296 25410 4352 25466
rect 4420 25410 4476 25466
rect 4544 25410 4600 25466
rect 4668 25410 4724 25466
rect 2808 25286 2864 25342
rect 2932 25286 2988 25342
rect 3056 25286 3112 25342
rect 3180 25286 3236 25342
rect 3304 25286 3360 25342
rect 3428 25286 3484 25342
rect 3552 25286 3608 25342
rect 3676 25286 3732 25342
rect 3800 25286 3856 25342
rect 3924 25286 3980 25342
rect 4048 25286 4104 25342
rect 4172 25286 4228 25342
rect 4296 25286 4352 25342
rect 4420 25286 4476 25342
rect 4544 25286 4600 25342
rect 4668 25286 4724 25342
rect 2808 25162 2864 25218
rect 2932 25162 2988 25218
rect 3056 25162 3112 25218
rect 3180 25162 3236 25218
rect 3304 25162 3360 25218
rect 3428 25162 3484 25218
rect 3552 25162 3608 25218
rect 3676 25162 3732 25218
rect 3800 25162 3856 25218
rect 3924 25162 3980 25218
rect 4048 25162 4104 25218
rect 4172 25162 4228 25218
rect 4296 25162 4352 25218
rect 4420 25162 4476 25218
rect 4544 25162 4600 25218
rect 4668 25162 4724 25218
rect 2808 25038 2864 25094
rect 2932 25038 2988 25094
rect 3056 25038 3112 25094
rect 3180 25038 3236 25094
rect 3304 25038 3360 25094
rect 3428 25038 3484 25094
rect 3552 25038 3608 25094
rect 3676 25038 3732 25094
rect 3800 25038 3856 25094
rect 3924 25038 3980 25094
rect 4048 25038 4104 25094
rect 4172 25038 4228 25094
rect 4296 25038 4352 25094
rect 4420 25038 4476 25094
rect 4544 25038 4600 25094
rect 4668 25038 4724 25094
rect 2808 24914 2864 24970
rect 2932 24914 2988 24970
rect 3056 24914 3112 24970
rect 3180 24914 3236 24970
rect 3304 24914 3360 24970
rect 3428 24914 3484 24970
rect 3552 24914 3608 24970
rect 3676 24914 3732 24970
rect 3800 24914 3856 24970
rect 3924 24914 3980 24970
rect 4048 24914 4104 24970
rect 4172 24914 4228 24970
rect 4296 24914 4352 24970
rect 4420 24914 4476 24970
rect 4544 24914 4600 24970
rect 4668 24914 4724 24970
rect 2808 24790 2864 24846
rect 2932 24790 2988 24846
rect 3056 24790 3112 24846
rect 3180 24790 3236 24846
rect 3304 24790 3360 24846
rect 3428 24790 3484 24846
rect 3552 24790 3608 24846
rect 3676 24790 3732 24846
rect 3800 24790 3856 24846
rect 3924 24790 3980 24846
rect 4048 24790 4104 24846
rect 4172 24790 4228 24846
rect 4296 24790 4352 24846
rect 4420 24790 4476 24846
rect 4544 24790 4600 24846
rect 4668 24790 4724 24846
rect 2808 24666 2864 24722
rect 2932 24666 2988 24722
rect 3056 24666 3112 24722
rect 3180 24666 3236 24722
rect 3304 24666 3360 24722
rect 3428 24666 3484 24722
rect 3552 24666 3608 24722
rect 3676 24666 3732 24722
rect 3800 24666 3856 24722
rect 3924 24666 3980 24722
rect 4048 24666 4104 24722
rect 4172 24666 4228 24722
rect 4296 24666 4352 24722
rect 4420 24666 4476 24722
rect 4544 24666 4600 24722
rect 4668 24666 4724 24722
rect 2808 24542 2864 24598
rect 2932 24542 2988 24598
rect 3056 24542 3112 24598
rect 3180 24542 3236 24598
rect 3304 24542 3360 24598
rect 3428 24542 3484 24598
rect 3552 24542 3608 24598
rect 3676 24542 3732 24598
rect 3800 24542 3856 24598
rect 3924 24542 3980 24598
rect 4048 24542 4104 24598
rect 4172 24542 4228 24598
rect 4296 24542 4352 24598
rect 4420 24542 4476 24598
rect 4544 24542 4600 24598
rect 4668 24542 4724 24598
rect 2808 24418 2864 24474
rect 2932 24418 2988 24474
rect 3056 24418 3112 24474
rect 3180 24418 3236 24474
rect 3304 24418 3360 24474
rect 3428 24418 3484 24474
rect 3552 24418 3608 24474
rect 3676 24418 3732 24474
rect 3800 24418 3856 24474
rect 3924 24418 3980 24474
rect 4048 24418 4104 24474
rect 4172 24418 4228 24474
rect 4296 24418 4352 24474
rect 4420 24418 4476 24474
rect 4544 24418 4600 24474
rect 4668 24418 4724 24474
rect 2808 24294 2864 24350
rect 2932 24294 2988 24350
rect 3056 24294 3112 24350
rect 3180 24294 3236 24350
rect 3304 24294 3360 24350
rect 3428 24294 3484 24350
rect 3552 24294 3608 24350
rect 3676 24294 3732 24350
rect 3800 24294 3856 24350
rect 3924 24294 3980 24350
rect 4048 24294 4104 24350
rect 4172 24294 4228 24350
rect 4296 24294 4352 24350
rect 4420 24294 4476 24350
rect 4544 24294 4600 24350
rect 4668 24294 4724 24350
rect 2808 24170 2864 24226
rect 2932 24170 2988 24226
rect 3056 24170 3112 24226
rect 3180 24170 3236 24226
rect 3304 24170 3360 24226
rect 3428 24170 3484 24226
rect 3552 24170 3608 24226
rect 3676 24170 3732 24226
rect 3800 24170 3856 24226
rect 3924 24170 3980 24226
rect 4048 24170 4104 24226
rect 4172 24170 4228 24226
rect 4296 24170 4352 24226
rect 4420 24170 4476 24226
rect 4544 24170 4600 24226
rect 4668 24170 4724 24226
rect 2808 24046 2864 24102
rect 2932 24046 2988 24102
rect 3056 24046 3112 24102
rect 3180 24046 3236 24102
rect 3304 24046 3360 24102
rect 3428 24046 3484 24102
rect 3552 24046 3608 24102
rect 3676 24046 3732 24102
rect 3800 24046 3856 24102
rect 3924 24046 3980 24102
rect 4048 24046 4104 24102
rect 4172 24046 4228 24102
rect 4296 24046 4352 24102
rect 4420 24046 4476 24102
rect 4544 24046 4600 24102
rect 4668 24046 4724 24102
rect 5178 26898 5234 26954
rect 5302 26898 5358 26954
rect 5426 26898 5482 26954
rect 5550 26898 5606 26954
rect 5674 26898 5730 26954
rect 5798 26898 5854 26954
rect 5922 26898 5978 26954
rect 6046 26898 6102 26954
rect 6170 26898 6226 26954
rect 6294 26898 6350 26954
rect 6418 26898 6474 26954
rect 6542 26898 6598 26954
rect 6666 26898 6722 26954
rect 6790 26898 6846 26954
rect 6914 26898 6970 26954
rect 7038 26898 7094 26954
rect 5178 26774 5234 26830
rect 5302 26774 5358 26830
rect 5426 26774 5482 26830
rect 5550 26774 5606 26830
rect 5674 26774 5730 26830
rect 5798 26774 5854 26830
rect 5922 26774 5978 26830
rect 6046 26774 6102 26830
rect 6170 26774 6226 26830
rect 6294 26774 6350 26830
rect 6418 26774 6474 26830
rect 6542 26774 6598 26830
rect 6666 26774 6722 26830
rect 6790 26774 6846 26830
rect 6914 26774 6970 26830
rect 7038 26774 7094 26830
rect 5178 26650 5234 26706
rect 5302 26650 5358 26706
rect 5426 26650 5482 26706
rect 5550 26650 5606 26706
rect 5674 26650 5730 26706
rect 5798 26650 5854 26706
rect 5922 26650 5978 26706
rect 6046 26650 6102 26706
rect 6170 26650 6226 26706
rect 6294 26650 6350 26706
rect 6418 26650 6474 26706
rect 6542 26650 6598 26706
rect 6666 26650 6722 26706
rect 6790 26650 6846 26706
rect 6914 26650 6970 26706
rect 7038 26650 7094 26706
rect 5178 26526 5234 26582
rect 5302 26526 5358 26582
rect 5426 26526 5482 26582
rect 5550 26526 5606 26582
rect 5674 26526 5730 26582
rect 5798 26526 5854 26582
rect 5922 26526 5978 26582
rect 6046 26526 6102 26582
rect 6170 26526 6226 26582
rect 6294 26526 6350 26582
rect 6418 26526 6474 26582
rect 6542 26526 6598 26582
rect 6666 26526 6722 26582
rect 6790 26526 6846 26582
rect 6914 26526 6970 26582
rect 7038 26526 7094 26582
rect 5178 26402 5234 26458
rect 5302 26402 5358 26458
rect 5426 26402 5482 26458
rect 5550 26402 5606 26458
rect 5674 26402 5730 26458
rect 5798 26402 5854 26458
rect 5922 26402 5978 26458
rect 6046 26402 6102 26458
rect 6170 26402 6226 26458
rect 6294 26402 6350 26458
rect 6418 26402 6474 26458
rect 6542 26402 6598 26458
rect 6666 26402 6722 26458
rect 6790 26402 6846 26458
rect 6914 26402 6970 26458
rect 7038 26402 7094 26458
rect 5178 26278 5234 26334
rect 5302 26278 5358 26334
rect 5426 26278 5482 26334
rect 5550 26278 5606 26334
rect 5674 26278 5730 26334
rect 5798 26278 5854 26334
rect 5922 26278 5978 26334
rect 6046 26278 6102 26334
rect 6170 26278 6226 26334
rect 6294 26278 6350 26334
rect 6418 26278 6474 26334
rect 6542 26278 6598 26334
rect 6666 26278 6722 26334
rect 6790 26278 6846 26334
rect 6914 26278 6970 26334
rect 7038 26278 7094 26334
rect 5178 26154 5234 26210
rect 5302 26154 5358 26210
rect 5426 26154 5482 26210
rect 5550 26154 5606 26210
rect 5674 26154 5730 26210
rect 5798 26154 5854 26210
rect 5922 26154 5978 26210
rect 6046 26154 6102 26210
rect 6170 26154 6226 26210
rect 6294 26154 6350 26210
rect 6418 26154 6474 26210
rect 6542 26154 6598 26210
rect 6666 26154 6722 26210
rect 6790 26154 6846 26210
rect 6914 26154 6970 26210
rect 7038 26154 7094 26210
rect 5178 26030 5234 26086
rect 5302 26030 5358 26086
rect 5426 26030 5482 26086
rect 5550 26030 5606 26086
rect 5674 26030 5730 26086
rect 5798 26030 5854 26086
rect 5922 26030 5978 26086
rect 6046 26030 6102 26086
rect 6170 26030 6226 26086
rect 6294 26030 6350 26086
rect 6418 26030 6474 26086
rect 6542 26030 6598 26086
rect 6666 26030 6722 26086
rect 6790 26030 6846 26086
rect 6914 26030 6970 26086
rect 7038 26030 7094 26086
rect 5178 25906 5234 25962
rect 5302 25906 5358 25962
rect 5426 25906 5482 25962
rect 5550 25906 5606 25962
rect 5674 25906 5730 25962
rect 5798 25906 5854 25962
rect 5922 25906 5978 25962
rect 6046 25906 6102 25962
rect 6170 25906 6226 25962
rect 6294 25906 6350 25962
rect 6418 25906 6474 25962
rect 6542 25906 6598 25962
rect 6666 25906 6722 25962
rect 6790 25906 6846 25962
rect 6914 25906 6970 25962
rect 7038 25906 7094 25962
rect 5178 25782 5234 25838
rect 5302 25782 5358 25838
rect 5426 25782 5482 25838
rect 5550 25782 5606 25838
rect 5674 25782 5730 25838
rect 5798 25782 5854 25838
rect 5922 25782 5978 25838
rect 6046 25782 6102 25838
rect 6170 25782 6226 25838
rect 6294 25782 6350 25838
rect 6418 25782 6474 25838
rect 6542 25782 6598 25838
rect 6666 25782 6722 25838
rect 6790 25782 6846 25838
rect 6914 25782 6970 25838
rect 7038 25782 7094 25838
rect 5178 25658 5234 25714
rect 5302 25658 5358 25714
rect 5426 25658 5482 25714
rect 5550 25658 5606 25714
rect 5674 25658 5730 25714
rect 5798 25658 5854 25714
rect 5922 25658 5978 25714
rect 6046 25658 6102 25714
rect 6170 25658 6226 25714
rect 6294 25658 6350 25714
rect 6418 25658 6474 25714
rect 6542 25658 6598 25714
rect 6666 25658 6722 25714
rect 6790 25658 6846 25714
rect 6914 25658 6970 25714
rect 7038 25658 7094 25714
rect 5178 25534 5234 25590
rect 5302 25534 5358 25590
rect 5426 25534 5482 25590
rect 5550 25534 5606 25590
rect 5674 25534 5730 25590
rect 5798 25534 5854 25590
rect 5922 25534 5978 25590
rect 6046 25534 6102 25590
rect 6170 25534 6226 25590
rect 6294 25534 6350 25590
rect 6418 25534 6474 25590
rect 6542 25534 6598 25590
rect 6666 25534 6722 25590
rect 6790 25534 6846 25590
rect 6914 25534 6970 25590
rect 7038 25534 7094 25590
rect 5178 25410 5234 25466
rect 5302 25410 5358 25466
rect 5426 25410 5482 25466
rect 5550 25410 5606 25466
rect 5674 25410 5730 25466
rect 5798 25410 5854 25466
rect 5922 25410 5978 25466
rect 6046 25410 6102 25466
rect 6170 25410 6226 25466
rect 6294 25410 6350 25466
rect 6418 25410 6474 25466
rect 6542 25410 6598 25466
rect 6666 25410 6722 25466
rect 6790 25410 6846 25466
rect 6914 25410 6970 25466
rect 7038 25410 7094 25466
rect 5178 25286 5234 25342
rect 5302 25286 5358 25342
rect 5426 25286 5482 25342
rect 5550 25286 5606 25342
rect 5674 25286 5730 25342
rect 5798 25286 5854 25342
rect 5922 25286 5978 25342
rect 6046 25286 6102 25342
rect 6170 25286 6226 25342
rect 6294 25286 6350 25342
rect 6418 25286 6474 25342
rect 6542 25286 6598 25342
rect 6666 25286 6722 25342
rect 6790 25286 6846 25342
rect 6914 25286 6970 25342
rect 7038 25286 7094 25342
rect 5178 25162 5234 25218
rect 5302 25162 5358 25218
rect 5426 25162 5482 25218
rect 5550 25162 5606 25218
rect 5674 25162 5730 25218
rect 5798 25162 5854 25218
rect 5922 25162 5978 25218
rect 6046 25162 6102 25218
rect 6170 25162 6226 25218
rect 6294 25162 6350 25218
rect 6418 25162 6474 25218
rect 6542 25162 6598 25218
rect 6666 25162 6722 25218
rect 6790 25162 6846 25218
rect 6914 25162 6970 25218
rect 7038 25162 7094 25218
rect 5178 25038 5234 25094
rect 5302 25038 5358 25094
rect 5426 25038 5482 25094
rect 5550 25038 5606 25094
rect 5674 25038 5730 25094
rect 5798 25038 5854 25094
rect 5922 25038 5978 25094
rect 6046 25038 6102 25094
rect 6170 25038 6226 25094
rect 6294 25038 6350 25094
rect 6418 25038 6474 25094
rect 6542 25038 6598 25094
rect 6666 25038 6722 25094
rect 6790 25038 6846 25094
rect 6914 25038 6970 25094
rect 7038 25038 7094 25094
rect 5178 24914 5234 24970
rect 5302 24914 5358 24970
rect 5426 24914 5482 24970
rect 5550 24914 5606 24970
rect 5674 24914 5730 24970
rect 5798 24914 5854 24970
rect 5922 24914 5978 24970
rect 6046 24914 6102 24970
rect 6170 24914 6226 24970
rect 6294 24914 6350 24970
rect 6418 24914 6474 24970
rect 6542 24914 6598 24970
rect 6666 24914 6722 24970
rect 6790 24914 6846 24970
rect 6914 24914 6970 24970
rect 7038 24914 7094 24970
rect 5178 24790 5234 24846
rect 5302 24790 5358 24846
rect 5426 24790 5482 24846
rect 5550 24790 5606 24846
rect 5674 24790 5730 24846
rect 5798 24790 5854 24846
rect 5922 24790 5978 24846
rect 6046 24790 6102 24846
rect 6170 24790 6226 24846
rect 6294 24790 6350 24846
rect 6418 24790 6474 24846
rect 6542 24790 6598 24846
rect 6666 24790 6722 24846
rect 6790 24790 6846 24846
rect 6914 24790 6970 24846
rect 7038 24790 7094 24846
rect 5178 24666 5234 24722
rect 5302 24666 5358 24722
rect 5426 24666 5482 24722
rect 5550 24666 5606 24722
rect 5674 24666 5730 24722
rect 5798 24666 5854 24722
rect 5922 24666 5978 24722
rect 6046 24666 6102 24722
rect 6170 24666 6226 24722
rect 6294 24666 6350 24722
rect 6418 24666 6474 24722
rect 6542 24666 6598 24722
rect 6666 24666 6722 24722
rect 6790 24666 6846 24722
rect 6914 24666 6970 24722
rect 7038 24666 7094 24722
rect 5178 24542 5234 24598
rect 5302 24542 5358 24598
rect 5426 24542 5482 24598
rect 5550 24542 5606 24598
rect 5674 24542 5730 24598
rect 5798 24542 5854 24598
rect 5922 24542 5978 24598
rect 6046 24542 6102 24598
rect 6170 24542 6226 24598
rect 6294 24542 6350 24598
rect 6418 24542 6474 24598
rect 6542 24542 6598 24598
rect 6666 24542 6722 24598
rect 6790 24542 6846 24598
rect 6914 24542 6970 24598
rect 7038 24542 7094 24598
rect 5178 24418 5234 24474
rect 5302 24418 5358 24474
rect 5426 24418 5482 24474
rect 5550 24418 5606 24474
rect 5674 24418 5730 24474
rect 5798 24418 5854 24474
rect 5922 24418 5978 24474
rect 6046 24418 6102 24474
rect 6170 24418 6226 24474
rect 6294 24418 6350 24474
rect 6418 24418 6474 24474
rect 6542 24418 6598 24474
rect 6666 24418 6722 24474
rect 6790 24418 6846 24474
rect 6914 24418 6970 24474
rect 7038 24418 7094 24474
rect 5178 24294 5234 24350
rect 5302 24294 5358 24350
rect 5426 24294 5482 24350
rect 5550 24294 5606 24350
rect 5674 24294 5730 24350
rect 5798 24294 5854 24350
rect 5922 24294 5978 24350
rect 6046 24294 6102 24350
rect 6170 24294 6226 24350
rect 6294 24294 6350 24350
rect 6418 24294 6474 24350
rect 6542 24294 6598 24350
rect 6666 24294 6722 24350
rect 6790 24294 6846 24350
rect 6914 24294 6970 24350
rect 7038 24294 7094 24350
rect 5178 24170 5234 24226
rect 5302 24170 5358 24226
rect 5426 24170 5482 24226
rect 5550 24170 5606 24226
rect 5674 24170 5730 24226
rect 5798 24170 5854 24226
rect 5922 24170 5978 24226
rect 6046 24170 6102 24226
rect 6170 24170 6226 24226
rect 6294 24170 6350 24226
rect 6418 24170 6474 24226
rect 6542 24170 6598 24226
rect 6666 24170 6722 24226
rect 6790 24170 6846 24226
rect 6914 24170 6970 24226
rect 7038 24170 7094 24226
rect 5178 24046 5234 24102
rect 5302 24046 5358 24102
rect 5426 24046 5482 24102
rect 5550 24046 5606 24102
rect 5674 24046 5730 24102
rect 5798 24046 5854 24102
rect 5922 24046 5978 24102
rect 6046 24046 6102 24102
rect 6170 24046 6226 24102
rect 6294 24046 6350 24102
rect 6418 24046 6474 24102
rect 6542 24046 6598 24102
rect 6666 24046 6722 24102
rect 6790 24046 6846 24102
rect 6914 24046 6970 24102
rect 7038 24046 7094 24102
rect 7884 26898 7940 26954
rect 8008 26898 8064 26954
rect 8132 26898 8188 26954
rect 8256 26898 8312 26954
rect 8380 26898 8436 26954
rect 8504 26898 8560 26954
rect 8628 26898 8684 26954
rect 8752 26898 8808 26954
rect 8876 26898 8932 26954
rect 9000 26898 9056 26954
rect 9124 26898 9180 26954
rect 9248 26898 9304 26954
rect 9372 26898 9428 26954
rect 9496 26898 9552 26954
rect 9620 26898 9676 26954
rect 9744 26898 9800 26954
rect 7884 26774 7940 26830
rect 8008 26774 8064 26830
rect 8132 26774 8188 26830
rect 8256 26774 8312 26830
rect 8380 26774 8436 26830
rect 8504 26774 8560 26830
rect 8628 26774 8684 26830
rect 8752 26774 8808 26830
rect 8876 26774 8932 26830
rect 9000 26774 9056 26830
rect 9124 26774 9180 26830
rect 9248 26774 9304 26830
rect 9372 26774 9428 26830
rect 9496 26774 9552 26830
rect 9620 26774 9676 26830
rect 9744 26774 9800 26830
rect 7884 26650 7940 26706
rect 8008 26650 8064 26706
rect 8132 26650 8188 26706
rect 8256 26650 8312 26706
rect 8380 26650 8436 26706
rect 8504 26650 8560 26706
rect 8628 26650 8684 26706
rect 8752 26650 8808 26706
rect 8876 26650 8932 26706
rect 9000 26650 9056 26706
rect 9124 26650 9180 26706
rect 9248 26650 9304 26706
rect 9372 26650 9428 26706
rect 9496 26650 9552 26706
rect 9620 26650 9676 26706
rect 9744 26650 9800 26706
rect 7884 26526 7940 26582
rect 8008 26526 8064 26582
rect 8132 26526 8188 26582
rect 8256 26526 8312 26582
rect 8380 26526 8436 26582
rect 8504 26526 8560 26582
rect 8628 26526 8684 26582
rect 8752 26526 8808 26582
rect 8876 26526 8932 26582
rect 9000 26526 9056 26582
rect 9124 26526 9180 26582
rect 9248 26526 9304 26582
rect 9372 26526 9428 26582
rect 9496 26526 9552 26582
rect 9620 26526 9676 26582
rect 9744 26526 9800 26582
rect 7884 26402 7940 26458
rect 8008 26402 8064 26458
rect 8132 26402 8188 26458
rect 8256 26402 8312 26458
rect 8380 26402 8436 26458
rect 8504 26402 8560 26458
rect 8628 26402 8684 26458
rect 8752 26402 8808 26458
rect 8876 26402 8932 26458
rect 9000 26402 9056 26458
rect 9124 26402 9180 26458
rect 9248 26402 9304 26458
rect 9372 26402 9428 26458
rect 9496 26402 9552 26458
rect 9620 26402 9676 26458
rect 9744 26402 9800 26458
rect 7884 26278 7940 26334
rect 8008 26278 8064 26334
rect 8132 26278 8188 26334
rect 8256 26278 8312 26334
rect 8380 26278 8436 26334
rect 8504 26278 8560 26334
rect 8628 26278 8684 26334
rect 8752 26278 8808 26334
rect 8876 26278 8932 26334
rect 9000 26278 9056 26334
rect 9124 26278 9180 26334
rect 9248 26278 9304 26334
rect 9372 26278 9428 26334
rect 9496 26278 9552 26334
rect 9620 26278 9676 26334
rect 9744 26278 9800 26334
rect 7884 26154 7940 26210
rect 8008 26154 8064 26210
rect 8132 26154 8188 26210
rect 8256 26154 8312 26210
rect 8380 26154 8436 26210
rect 8504 26154 8560 26210
rect 8628 26154 8684 26210
rect 8752 26154 8808 26210
rect 8876 26154 8932 26210
rect 9000 26154 9056 26210
rect 9124 26154 9180 26210
rect 9248 26154 9304 26210
rect 9372 26154 9428 26210
rect 9496 26154 9552 26210
rect 9620 26154 9676 26210
rect 9744 26154 9800 26210
rect 7884 26030 7940 26086
rect 8008 26030 8064 26086
rect 8132 26030 8188 26086
rect 8256 26030 8312 26086
rect 8380 26030 8436 26086
rect 8504 26030 8560 26086
rect 8628 26030 8684 26086
rect 8752 26030 8808 26086
rect 8876 26030 8932 26086
rect 9000 26030 9056 26086
rect 9124 26030 9180 26086
rect 9248 26030 9304 26086
rect 9372 26030 9428 26086
rect 9496 26030 9552 26086
rect 9620 26030 9676 26086
rect 9744 26030 9800 26086
rect 7884 25906 7940 25962
rect 8008 25906 8064 25962
rect 8132 25906 8188 25962
rect 8256 25906 8312 25962
rect 8380 25906 8436 25962
rect 8504 25906 8560 25962
rect 8628 25906 8684 25962
rect 8752 25906 8808 25962
rect 8876 25906 8932 25962
rect 9000 25906 9056 25962
rect 9124 25906 9180 25962
rect 9248 25906 9304 25962
rect 9372 25906 9428 25962
rect 9496 25906 9552 25962
rect 9620 25906 9676 25962
rect 9744 25906 9800 25962
rect 7884 25782 7940 25838
rect 8008 25782 8064 25838
rect 8132 25782 8188 25838
rect 8256 25782 8312 25838
rect 8380 25782 8436 25838
rect 8504 25782 8560 25838
rect 8628 25782 8684 25838
rect 8752 25782 8808 25838
rect 8876 25782 8932 25838
rect 9000 25782 9056 25838
rect 9124 25782 9180 25838
rect 9248 25782 9304 25838
rect 9372 25782 9428 25838
rect 9496 25782 9552 25838
rect 9620 25782 9676 25838
rect 9744 25782 9800 25838
rect 7884 25658 7940 25714
rect 8008 25658 8064 25714
rect 8132 25658 8188 25714
rect 8256 25658 8312 25714
rect 8380 25658 8436 25714
rect 8504 25658 8560 25714
rect 8628 25658 8684 25714
rect 8752 25658 8808 25714
rect 8876 25658 8932 25714
rect 9000 25658 9056 25714
rect 9124 25658 9180 25714
rect 9248 25658 9304 25714
rect 9372 25658 9428 25714
rect 9496 25658 9552 25714
rect 9620 25658 9676 25714
rect 9744 25658 9800 25714
rect 7884 25534 7940 25590
rect 8008 25534 8064 25590
rect 8132 25534 8188 25590
rect 8256 25534 8312 25590
rect 8380 25534 8436 25590
rect 8504 25534 8560 25590
rect 8628 25534 8684 25590
rect 8752 25534 8808 25590
rect 8876 25534 8932 25590
rect 9000 25534 9056 25590
rect 9124 25534 9180 25590
rect 9248 25534 9304 25590
rect 9372 25534 9428 25590
rect 9496 25534 9552 25590
rect 9620 25534 9676 25590
rect 9744 25534 9800 25590
rect 7884 25410 7940 25466
rect 8008 25410 8064 25466
rect 8132 25410 8188 25466
rect 8256 25410 8312 25466
rect 8380 25410 8436 25466
rect 8504 25410 8560 25466
rect 8628 25410 8684 25466
rect 8752 25410 8808 25466
rect 8876 25410 8932 25466
rect 9000 25410 9056 25466
rect 9124 25410 9180 25466
rect 9248 25410 9304 25466
rect 9372 25410 9428 25466
rect 9496 25410 9552 25466
rect 9620 25410 9676 25466
rect 9744 25410 9800 25466
rect 7884 25286 7940 25342
rect 8008 25286 8064 25342
rect 8132 25286 8188 25342
rect 8256 25286 8312 25342
rect 8380 25286 8436 25342
rect 8504 25286 8560 25342
rect 8628 25286 8684 25342
rect 8752 25286 8808 25342
rect 8876 25286 8932 25342
rect 9000 25286 9056 25342
rect 9124 25286 9180 25342
rect 9248 25286 9304 25342
rect 9372 25286 9428 25342
rect 9496 25286 9552 25342
rect 9620 25286 9676 25342
rect 9744 25286 9800 25342
rect 7884 25162 7940 25218
rect 8008 25162 8064 25218
rect 8132 25162 8188 25218
rect 8256 25162 8312 25218
rect 8380 25162 8436 25218
rect 8504 25162 8560 25218
rect 8628 25162 8684 25218
rect 8752 25162 8808 25218
rect 8876 25162 8932 25218
rect 9000 25162 9056 25218
rect 9124 25162 9180 25218
rect 9248 25162 9304 25218
rect 9372 25162 9428 25218
rect 9496 25162 9552 25218
rect 9620 25162 9676 25218
rect 9744 25162 9800 25218
rect 7884 25038 7940 25094
rect 8008 25038 8064 25094
rect 8132 25038 8188 25094
rect 8256 25038 8312 25094
rect 8380 25038 8436 25094
rect 8504 25038 8560 25094
rect 8628 25038 8684 25094
rect 8752 25038 8808 25094
rect 8876 25038 8932 25094
rect 9000 25038 9056 25094
rect 9124 25038 9180 25094
rect 9248 25038 9304 25094
rect 9372 25038 9428 25094
rect 9496 25038 9552 25094
rect 9620 25038 9676 25094
rect 9744 25038 9800 25094
rect 7884 24914 7940 24970
rect 8008 24914 8064 24970
rect 8132 24914 8188 24970
rect 8256 24914 8312 24970
rect 8380 24914 8436 24970
rect 8504 24914 8560 24970
rect 8628 24914 8684 24970
rect 8752 24914 8808 24970
rect 8876 24914 8932 24970
rect 9000 24914 9056 24970
rect 9124 24914 9180 24970
rect 9248 24914 9304 24970
rect 9372 24914 9428 24970
rect 9496 24914 9552 24970
rect 9620 24914 9676 24970
rect 9744 24914 9800 24970
rect 7884 24790 7940 24846
rect 8008 24790 8064 24846
rect 8132 24790 8188 24846
rect 8256 24790 8312 24846
rect 8380 24790 8436 24846
rect 8504 24790 8560 24846
rect 8628 24790 8684 24846
rect 8752 24790 8808 24846
rect 8876 24790 8932 24846
rect 9000 24790 9056 24846
rect 9124 24790 9180 24846
rect 9248 24790 9304 24846
rect 9372 24790 9428 24846
rect 9496 24790 9552 24846
rect 9620 24790 9676 24846
rect 9744 24790 9800 24846
rect 7884 24666 7940 24722
rect 8008 24666 8064 24722
rect 8132 24666 8188 24722
rect 8256 24666 8312 24722
rect 8380 24666 8436 24722
rect 8504 24666 8560 24722
rect 8628 24666 8684 24722
rect 8752 24666 8808 24722
rect 8876 24666 8932 24722
rect 9000 24666 9056 24722
rect 9124 24666 9180 24722
rect 9248 24666 9304 24722
rect 9372 24666 9428 24722
rect 9496 24666 9552 24722
rect 9620 24666 9676 24722
rect 9744 24666 9800 24722
rect 7884 24542 7940 24598
rect 8008 24542 8064 24598
rect 8132 24542 8188 24598
rect 8256 24542 8312 24598
rect 8380 24542 8436 24598
rect 8504 24542 8560 24598
rect 8628 24542 8684 24598
rect 8752 24542 8808 24598
rect 8876 24542 8932 24598
rect 9000 24542 9056 24598
rect 9124 24542 9180 24598
rect 9248 24542 9304 24598
rect 9372 24542 9428 24598
rect 9496 24542 9552 24598
rect 9620 24542 9676 24598
rect 9744 24542 9800 24598
rect 7884 24418 7940 24474
rect 8008 24418 8064 24474
rect 8132 24418 8188 24474
rect 8256 24418 8312 24474
rect 8380 24418 8436 24474
rect 8504 24418 8560 24474
rect 8628 24418 8684 24474
rect 8752 24418 8808 24474
rect 8876 24418 8932 24474
rect 9000 24418 9056 24474
rect 9124 24418 9180 24474
rect 9248 24418 9304 24474
rect 9372 24418 9428 24474
rect 9496 24418 9552 24474
rect 9620 24418 9676 24474
rect 9744 24418 9800 24474
rect 7884 24294 7940 24350
rect 8008 24294 8064 24350
rect 8132 24294 8188 24350
rect 8256 24294 8312 24350
rect 8380 24294 8436 24350
rect 8504 24294 8560 24350
rect 8628 24294 8684 24350
rect 8752 24294 8808 24350
rect 8876 24294 8932 24350
rect 9000 24294 9056 24350
rect 9124 24294 9180 24350
rect 9248 24294 9304 24350
rect 9372 24294 9428 24350
rect 9496 24294 9552 24350
rect 9620 24294 9676 24350
rect 9744 24294 9800 24350
rect 7884 24170 7940 24226
rect 8008 24170 8064 24226
rect 8132 24170 8188 24226
rect 8256 24170 8312 24226
rect 8380 24170 8436 24226
rect 8504 24170 8560 24226
rect 8628 24170 8684 24226
rect 8752 24170 8808 24226
rect 8876 24170 8932 24226
rect 9000 24170 9056 24226
rect 9124 24170 9180 24226
rect 9248 24170 9304 24226
rect 9372 24170 9428 24226
rect 9496 24170 9552 24226
rect 9620 24170 9676 24226
rect 9744 24170 9800 24226
rect 7884 24046 7940 24102
rect 8008 24046 8064 24102
rect 8132 24046 8188 24102
rect 8256 24046 8312 24102
rect 8380 24046 8436 24102
rect 8504 24046 8560 24102
rect 8628 24046 8684 24102
rect 8752 24046 8808 24102
rect 8876 24046 8932 24102
rect 9000 24046 9056 24102
rect 9124 24046 9180 24102
rect 9248 24046 9304 24102
rect 9372 24046 9428 24102
rect 9496 24046 9552 24102
rect 9620 24046 9676 24102
rect 9744 24046 9800 24102
rect 10254 26898 10310 26954
rect 10378 26898 10434 26954
rect 10502 26898 10558 26954
rect 10626 26898 10682 26954
rect 10750 26898 10806 26954
rect 10874 26898 10930 26954
rect 10998 26898 11054 26954
rect 11122 26898 11178 26954
rect 11246 26898 11302 26954
rect 11370 26898 11426 26954
rect 11494 26898 11550 26954
rect 11618 26898 11674 26954
rect 11742 26898 11798 26954
rect 11866 26898 11922 26954
rect 11990 26898 12046 26954
rect 12114 26898 12170 26954
rect 10254 26774 10310 26830
rect 10378 26774 10434 26830
rect 10502 26774 10558 26830
rect 10626 26774 10682 26830
rect 10750 26774 10806 26830
rect 10874 26774 10930 26830
rect 10998 26774 11054 26830
rect 11122 26774 11178 26830
rect 11246 26774 11302 26830
rect 11370 26774 11426 26830
rect 11494 26774 11550 26830
rect 11618 26774 11674 26830
rect 11742 26774 11798 26830
rect 11866 26774 11922 26830
rect 11990 26774 12046 26830
rect 12114 26774 12170 26830
rect 10254 26650 10310 26706
rect 10378 26650 10434 26706
rect 10502 26650 10558 26706
rect 10626 26650 10682 26706
rect 10750 26650 10806 26706
rect 10874 26650 10930 26706
rect 10998 26650 11054 26706
rect 11122 26650 11178 26706
rect 11246 26650 11302 26706
rect 11370 26650 11426 26706
rect 11494 26650 11550 26706
rect 11618 26650 11674 26706
rect 11742 26650 11798 26706
rect 11866 26650 11922 26706
rect 11990 26650 12046 26706
rect 12114 26650 12170 26706
rect 10254 26526 10310 26582
rect 10378 26526 10434 26582
rect 10502 26526 10558 26582
rect 10626 26526 10682 26582
rect 10750 26526 10806 26582
rect 10874 26526 10930 26582
rect 10998 26526 11054 26582
rect 11122 26526 11178 26582
rect 11246 26526 11302 26582
rect 11370 26526 11426 26582
rect 11494 26526 11550 26582
rect 11618 26526 11674 26582
rect 11742 26526 11798 26582
rect 11866 26526 11922 26582
rect 11990 26526 12046 26582
rect 12114 26526 12170 26582
rect 10254 26402 10310 26458
rect 10378 26402 10434 26458
rect 10502 26402 10558 26458
rect 10626 26402 10682 26458
rect 10750 26402 10806 26458
rect 10874 26402 10930 26458
rect 10998 26402 11054 26458
rect 11122 26402 11178 26458
rect 11246 26402 11302 26458
rect 11370 26402 11426 26458
rect 11494 26402 11550 26458
rect 11618 26402 11674 26458
rect 11742 26402 11798 26458
rect 11866 26402 11922 26458
rect 11990 26402 12046 26458
rect 12114 26402 12170 26458
rect 10254 26278 10310 26334
rect 10378 26278 10434 26334
rect 10502 26278 10558 26334
rect 10626 26278 10682 26334
rect 10750 26278 10806 26334
rect 10874 26278 10930 26334
rect 10998 26278 11054 26334
rect 11122 26278 11178 26334
rect 11246 26278 11302 26334
rect 11370 26278 11426 26334
rect 11494 26278 11550 26334
rect 11618 26278 11674 26334
rect 11742 26278 11798 26334
rect 11866 26278 11922 26334
rect 11990 26278 12046 26334
rect 12114 26278 12170 26334
rect 10254 26154 10310 26210
rect 10378 26154 10434 26210
rect 10502 26154 10558 26210
rect 10626 26154 10682 26210
rect 10750 26154 10806 26210
rect 10874 26154 10930 26210
rect 10998 26154 11054 26210
rect 11122 26154 11178 26210
rect 11246 26154 11302 26210
rect 11370 26154 11426 26210
rect 11494 26154 11550 26210
rect 11618 26154 11674 26210
rect 11742 26154 11798 26210
rect 11866 26154 11922 26210
rect 11990 26154 12046 26210
rect 12114 26154 12170 26210
rect 10254 26030 10310 26086
rect 10378 26030 10434 26086
rect 10502 26030 10558 26086
rect 10626 26030 10682 26086
rect 10750 26030 10806 26086
rect 10874 26030 10930 26086
rect 10998 26030 11054 26086
rect 11122 26030 11178 26086
rect 11246 26030 11302 26086
rect 11370 26030 11426 26086
rect 11494 26030 11550 26086
rect 11618 26030 11674 26086
rect 11742 26030 11798 26086
rect 11866 26030 11922 26086
rect 11990 26030 12046 26086
rect 12114 26030 12170 26086
rect 10254 25906 10310 25962
rect 10378 25906 10434 25962
rect 10502 25906 10558 25962
rect 10626 25906 10682 25962
rect 10750 25906 10806 25962
rect 10874 25906 10930 25962
rect 10998 25906 11054 25962
rect 11122 25906 11178 25962
rect 11246 25906 11302 25962
rect 11370 25906 11426 25962
rect 11494 25906 11550 25962
rect 11618 25906 11674 25962
rect 11742 25906 11798 25962
rect 11866 25906 11922 25962
rect 11990 25906 12046 25962
rect 12114 25906 12170 25962
rect 10254 25782 10310 25838
rect 10378 25782 10434 25838
rect 10502 25782 10558 25838
rect 10626 25782 10682 25838
rect 10750 25782 10806 25838
rect 10874 25782 10930 25838
rect 10998 25782 11054 25838
rect 11122 25782 11178 25838
rect 11246 25782 11302 25838
rect 11370 25782 11426 25838
rect 11494 25782 11550 25838
rect 11618 25782 11674 25838
rect 11742 25782 11798 25838
rect 11866 25782 11922 25838
rect 11990 25782 12046 25838
rect 12114 25782 12170 25838
rect 10254 25658 10310 25714
rect 10378 25658 10434 25714
rect 10502 25658 10558 25714
rect 10626 25658 10682 25714
rect 10750 25658 10806 25714
rect 10874 25658 10930 25714
rect 10998 25658 11054 25714
rect 11122 25658 11178 25714
rect 11246 25658 11302 25714
rect 11370 25658 11426 25714
rect 11494 25658 11550 25714
rect 11618 25658 11674 25714
rect 11742 25658 11798 25714
rect 11866 25658 11922 25714
rect 11990 25658 12046 25714
rect 12114 25658 12170 25714
rect 10254 25534 10310 25590
rect 10378 25534 10434 25590
rect 10502 25534 10558 25590
rect 10626 25534 10682 25590
rect 10750 25534 10806 25590
rect 10874 25534 10930 25590
rect 10998 25534 11054 25590
rect 11122 25534 11178 25590
rect 11246 25534 11302 25590
rect 11370 25534 11426 25590
rect 11494 25534 11550 25590
rect 11618 25534 11674 25590
rect 11742 25534 11798 25590
rect 11866 25534 11922 25590
rect 11990 25534 12046 25590
rect 12114 25534 12170 25590
rect 10254 25410 10310 25466
rect 10378 25410 10434 25466
rect 10502 25410 10558 25466
rect 10626 25410 10682 25466
rect 10750 25410 10806 25466
rect 10874 25410 10930 25466
rect 10998 25410 11054 25466
rect 11122 25410 11178 25466
rect 11246 25410 11302 25466
rect 11370 25410 11426 25466
rect 11494 25410 11550 25466
rect 11618 25410 11674 25466
rect 11742 25410 11798 25466
rect 11866 25410 11922 25466
rect 11990 25410 12046 25466
rect 12114 25410 12170 25466
rect 10254 25286 10310 25342
rect 10378 25286 10434 25342
rect 10502 25286 10558 25342
rect 10626 25286 10682 25342
rect 10750 25286 10806 25342
rect 10874 25286 10930 25342
rect 10998 25286 11054 25342
rect 11122 25286 11178 25342
rect 11246 25286 11302 25342
rect 11370 25286 11426 25342
rect 11494 25286 11550 25342
rect 11618 25286 11674 25342
rect 11742 25286 11798 25342
rect 11866 25286 11922 25342
rect 11990 25286 12046 25342
rect 12114 25286 12170 25342
rect 10254 25162 10310 25218
rect 10378 25162 10434 25218
rect 10502 25162 10558 25218
rect 10626 25162 10682 25218
rect 10750 25162 10806 25218
rect 10874 25162 10930 25218
rect 10998 25162 11054 25218
rect 11122 25162 11178 25218
rect 11246 25162 11302 25218
rect 11370 25162 11426 25218
rect 11494 25162 11550 25218
rect 11618 25162 11674 25218
rect 11742 25162 11798 25218
rect 11866 25162 11922 25218
rect 11990 25162 12046 25218
rect 12114 25162 12170 25218
rect 10254 25038 10310 25094
rect 10378 25038 10434 25094
rect 10502 25038 10558 25094
rect 10626 25038 10682 25094
rect 10750 25038 10806 25094
rect 10874 25038 10930 25094
rect 10998 25038 11054 25094
rect 11122 25038 11178 25094
rect 11246 25038 11302 25094
rect 11370 25038 11426 25094
rect 11494 25038 11550 25094
rect 11618 25038 11674 25094
rect 11742 25038 11798 25094
rect 11866 25038 11922 25094
rect 11990 25038 12046 25094
rect 12114 25038 12170 25094
rect 10254 24914 10310 24970
rect 10378 24914 10434 24970
rect 10502 24914 10558 24970
rect 10626 24914 10682 24970
rect 10750 24914 10806 24970
rect 10874 24914 10930 24970
rect 10998 24914 11054 24970
rect 11122 24914 11178 24970
rect 11246 24914 11302 24970
rect 11370 24914 11426 24970
rect 11494 24914 11550 24970
rect 11618 24914 11674 24970
rect 11742 24914 11798 24970
rect 11866 24914 11922 24970
rect 11990 24914 12046 24970
rect 12114 24914 12170 24970
rect 10254 24790 10310 24846
rect 10378 24790 10434 24846
rect 10502 24790 10558 24846
rect 10626 24790 10682 24846
rect 10750 24790 10806 24846
rect 10874 24790 10930 24846
rect 10998 24790 11054 24846
rect 11122 24790 11178 24846
rect 11246 24790 11302 24846
rect 11370 24790 11426 24846
rect 11494 24790 11550 24846
rect 11618 24790 11674 24846
rect 11742 24790 11798 24846
rect 11866 24790 11922 24846
rect 11990 24790 12046 24846
rect 12114 24790 12170 24846
rect 10254 24666 10310 24722
rect 10378 24666 10434 24722
rect 10502 24666 10558 24722
rect 10626 24666 10682 24722
rect 10750 24666 10806 24722
rect 10874 24666 10930 24722
rect 10998 24666 11054 24722
rect 11122 24666 11178 24722
rect 11246 24666 11302 24722
rect 11370 24666 11426 24722
rect 11494 24666 11550 24722
rect 11618 24666 11674 24722
rect 11742 24666 11798 24722
rect 11866 24666 11922 24722
rect 11990 24666 12046 24722
rect 12114 24666 12170 24722
rect 10254 24542 10310 24598
rect 10378 24542 10434 24598
rect 10502 24542 10558 24598
rect 10626 24542 10682 24598
rect 10750 24542 10806 24598
rect 10874 24542 10930 24598
rect 10998 24542 11054 24598
rect 11122 24542 11178 24598
rect 11246 24542 11302 24598
rect 11370 24542 11426 24598
rect 11494 24542 11550 24598
rect 11618 24542 11674 24598
rect 11742 24542 11798 24598
rect 11866 24542 11922 24598
rect 11990 24542 12046 24598
rect 12114 24542 12170 24598
rect 10254 24418 10310 24474
rect 10378 24418 10434 24474
rect 10502 24418 10558 24474
rect 10626 24418 10682 24474
rect 10750 24418 10806 24474
rect 10874 24418 10930 24474
rect 10998 24418 11054 24474
rect 11122 24418 11178 24474
rect 11246 24418 11302 24474
rect 11370 24418 11426 24474
rect 11494 24418 11550 24474
rect 11618 24418 11674 24474
rect 11742 24418 11798 24474
rect 11866 24418 11922 24474
rect 11990 24418 12046 24474
rect 12114 24418 12170 24474
rect 10254 24294 10310 24350
rect 10378 24294 10434 24350
rect 10502 24294 10558 24350
rect 10626 24294 10682 24350
rect 10750 24294 10806 24350
rect 10874 24294 10930 24350
rect 10998 24294 11054 24350
rect 11122 24294 11178 24350
rect 11246 24294 11302 24350
rect 11370 24294 11426 24350
rect 11494 24294 11550 24350
rect 11618 24294 11674 24350
rect 11742 24294 11798 24350
rect 11866 24294 11922 24350
rect 11990 24294 12046 24350
rect 12114 24294 12170 24350
rect 10254 24170 10310 24226
rect 10378 24170 10434 24226
rect 10502 24170 10558 24226
rect 10626 24170 10682 24226
rect 10750 24170 10806 24226
rect 10874 24170 10930 24226
rect 10998 24170 11054 24226
rect 11122 24170 11178 24226
rect 11246 24170 11302 24226
rect 11370 24170 11426 24226
rect 11494 24170 11550 24226
rect 11618 24170 11674 24226
rect 11742 24170 11798 24226
rect 11866 24170 11922 24226
rect 11990 24170 12046 24226
rect 12114 24170 12170 24226
rect 10254 24046 10310 24102
rect 10378 24046 10434 24102
rect 10502 24046 10558 24102
rect 10626 24046 10682 24102
rect 10750 24046 10806 24102
rect 10874 24046 10930 24102
rect 10998 24046 11054 24102
rect 11122 24046 11178 24102
rect 11246 24046 11302 24102
rect 11370 24046 11426 24102
rect 11494 24046 11550 24102
rect 11618 24046 11674 24102
rect 11742 24046 11798 24102
rect 11866 24046 11922 24102
rect 11990 24046 12046 24102
rect 12114 24046 12170 24102
rect 12871 26898 12927 26954
rect 12995 26898 13051 26954
rect 13119 26898 13175 26954
rect 13243 26898 13299 26954
rect 13367 26898 13423 26954
rect 13491 26898 13547 26954
rect 13615 26898 13671 26954
rect 13739 26898 13795 26954
rect 13863 26898 13919 26954
rect 13987 26898 14043 26954
rect 14111 26898 14167 26954
rect 14235 26898 14291 26954
rect 14359 26898 14415 26954
rect 14483 26898 14539 26954
rect 14607 26898 14663 26954
rect 12871 26774 12927 26830
rect 12995 26774 13051 26830
rect 13119 26774 13175 26830
rect 13243 26774 13299 26830
rect 13367 26774 13423 26830
rect 13491 26774 13547 26830
rect 13615 26774 13671 26830
rect 13739 26774 13795 26830
rect 13863 26774 13919 26830
rect 13987 26774 14043 26830
rect 14111 26774 14167 26830
rect 14235 26774 14291 26830
rect 14359 26774 14415 26830
rect 14483 26774 14539 26830
rect 14607 26774 14663 26830
rect 12871 26650 12927 26706
rect 12995 26650 13051 26706
rect 13119 26650 13175 26706
rect 13243 26650 13299 26706
rect 13367 26650 13423 26706
rect 13491 26650 13547 26706
rect 13615 26650 13671 26706
rect 13739 26650 13795 26706
rect 13863 26650 13919 26706
rect 13987 26650 14043 26706
rect 14111 26650 14167 26706
rect 14235 26650 14291 26706
rect 14359 26650 14415 26706
rect 14483 26650 14539 26706
rect 14607 26650 14663 26706
rect 12871 26526 12927 26582
rect 12995 26526 13051 26582
rect 13119 26526 13175 26582
rect 13243 26526 13299 26582
rect 13367 26526 13423 26582
rect 13491 26526 13547 26582
rect 13615 26526 13671 26582
rect 13739 26526 13795 26582
rect 13863 26526 13919 26582
rect 13987 26526 14043 26582
rect 14111 26526 14167 26582
rect 14235 26526 14291 26582
rect 14359 26526 14415 26582
rect 14483 26526 14539 26582
rect 14607 26526 14663 26582
rect 12871 26402 12927 26458
rect 12995 26402 13051 26458
rect 13119 26402 13175 26458
rect 13243 26402 13299 26458
rect 13367 26402 13423 26458
rect 13491 26402 13547 26458
rect 13615 26402 13671 26458
rect 13739 26402 13795 26458
rect 13863 26402 13919 26458
rect 13987 26402 14043 26458
rect 14111 26402 14167 26458
rect 14235 26402 14291 26458
rect 14359 26402 14415 26458
rect 14483 26402 14539 26458
rect 14607 26402 14663 26458
rect 12871 26278 12927 26334
rect 12995 26278 13051 26334
rect 13119 26278 13175 26334
rect 13243 26278 13299 26334
rect 13367 26278 13423 26334
rect 13491 26278 13547 26334
rect 13615 26278 13671 26334
rect 13739 26278 13795 26334
rect 13863 26278 13919 26334
rect 13987 26278 14043 26334
rect 14111 26278 14167 26334
rect 14235 26278 14291 26334
rect 14359 26278 14415 26334
rect 14483 26278 14539 26334
rect 14607 26278 14663 26334
rect 12871 26154 12927 26210
rect 12995 26154 13051 26210
rect 13119 26154 13175 26210
rect 13243 26154 13299 26210
rect 13367 26154 13423 26210
rect 13491 26154 13547 26210
rect 13615 26154 13671 26210
rect 13739 26154 13795 26210
rect 13863 26154 13919 26210
rect 13987 26154 14043 26210
rect 14111 26154 14167 26210
rect 14235 26154 14291 26210
rect 14359 26154 14415 26210
rect 14483 26154 14539 26210
rect 14607 26154 14663 26210
rect 12871 26030 12927 26086
rect 12995 26030 13051 26086
rect 13119 26030 13175 26086
rect 13243 26030 13299 26086
rect 13367 26030 13423 26086
rect 13491 26030 13547 26086
rect 13615 26030 13671 26086
rect 13739 26030 13795 26086
rect 13863 26030 13919 26086
rect 13987 26030 14043 26086
rect 14111 26030 14167 26086
rect 14235 26030 14291 26086
rect 14359 26030 14415 26086
rect 14483 26030 14539 26086
rect 14607 26030 14663 26086
rect 12871 25906 12927 25962
rect 12995 25906 13051 25962
rect 13119 25906 13175 25962
rect 13243 25906 13299 25962
rect 13367 25906 13423 25962
rect 13491 25906 13547 25962
rect 13615 25906 13671 25962
rect 13739 25906 13795 25962
rect 13863 25906 13919 25962
rect 13987 25906 14043 25962
rect 14111 25906 14167 25962
rect 14235 25906 14291 25962
rect 14359 25906 14415 25962
rect 14483 25906 14539 25962
rect 14607 25906 14663 25962
rect 12871 25782 12927 25838
rect 12995 25782 13051 25838
rect 13119 25782 13175 25838
rect 13243 25782 13299 25838
rect 13367 25782 13423 25838
rect 13491 25782 13547 25838
rect 13615 25782 13671 25838
rect 13739 25782 13795 25838
rect 13863 25782 13919 25838
rect 13987 25782 14043 25838
rect 14111 25782 14167 25838
rect 14235 25782 14291 25838
rect 14359 25782 14415 25838
rect 14483 25782 14539 25838
rect 14607 25782 14663 25838
rect 12871 25658 12927 25714
rect 12995 25658 13051 25714
rect 13119 25658 13175 25714
rect 13243 25658 13299 25714
rect 13367 25658 13423 25714
rect 13491 25658 13547 25714
rect 13615 25658 13671 25714
rect 13739 25658 13795 25714
rect 13863 25658 13919 25714
rect 13987 25658 14043 25714
rect 14111 25658 14167 25714
rect 14235 25658 14291 25714
rect 14359 25658 14415 25714
rect 14483 25658 14539 25714
rect 14607 25658 14663 25714
rect 12871 25534 12927 25590
rect 12995 25534 13051 25590
rect 13119 25534 13175 25590
rect 13243 25534 13299 25590
rect 13367 25534 13423 25590
rect 13491 25534 13547 25590
rect 13615 25534 13671 25590
rect 13739 25534 13795 25590
rect 13863 25534 13919 25590
rect 13987 25534 14043 25590
rect 14111 25534 14167 25590
rect 14235 25534 14291 25590
rect 14359 25534 14415 25590
rect 14483 25534 14539 25590
rect 14607 25534 14663 25590
rect 12871 25410 12927 25466
rect 12995 25410 13051 25466
rect 13119 25410 13175 25466
rect 13243 25410 13299 25466
rect 13367 25410 13423 25466
rect 13491 25410 13547 25466
rect 13615 25410 13671 25466
rect 13739 25410 13795 25466
rect 13863 25410 13919 25466
rect 13987 25410 14043 25466
rect 14111 25410 14167 25466
rect 14235 25410 14291 25466
rect 14359 25410 14415 25466
rect 14483 25410 14539 25466
rect 14607 25410 14663 25466
rect 12871 25286 12927 25342
rect 12995 25286 13051 25342
rect 13119 25286 13175 25342
rect 13243 25286 13299 25342
rect 13367 25286 13423 25342
rect 13491 25286 13547 25342
rect 13615 25286 13671 25342
rect 13739 25286 13795 25342
rect 13863 25286 13919 25342
rect 13987 25286 14043 25342
rect 14111 25286 14167 25342
rect 14235 25286 14291 25342
rect 14359 25286 14415 25342
rect 14483 25286 14539 25342
rect 14607 25286 14663 25342
rect 12871 25162 12927 25218
rect 12995 25162 13051 25218
rect 13119 25162 13175 25218
rect 13243 25162 13299 25218
rect 13367 25162 13423 25218
rect 13491 25162 13547 25218
rect 13615 25162 13671 25218
rect 13739 25162 13795 25218
rect 13863 25162 13919 25218
rect 13987 25162 14043 25218
rect 14111 25162 14167 25218
rect 14235 25162 14291 25218
rect 14359 25162 14415 25218
rect 14483 25162 14539 25218
rect 14607 25162 14663 25218
rect 12871 25038 12927 25094
rect 12995 25038 13051 25094
rect 13119 25038 13175 25094
rect 13243 25038 13299 25094
rect 13367 25038 13423 25094
rect 13491 25038 13547 25094
rect 13615 25038 13671 25094
rect 13739 25038 13795 25094
rect 13863 25038 13919 25094
rect 13987 25038 14043 25094
rect 14111 25038 14167 25094
rect 14235 25038 14291 25094
rect 14359 25038 14415 25094
rect 14483 25038 14539 25094
rect 14607 25038 14663 25094
rect 12871 24914 12927 24970
rect 12995 24914 13051 24970
rect 13119 24914 13175 24970
rect 13243 24914 13299 24970
rect 13367 24914 13423 24970
rect 13491 24914 13547 24970
rect 13615 24914 13671 24970
rect 13739 24914 13795 24970
rect 13863 24914 13919 24970
rect 13987 24914 14043 24970
rect 14111 24914 14167 24970
rect 14235 24914 14291 24970
rect 14359 24914 14415 24970
rect 14483 24914 14539 24970
rect 14607 24914 14663 24970
rect 12871 24790 12927 24846
rect 12995 24790 13051 24846
rect 13119 24790 13175 24846
rect 13243 24790 13299 24846
rect 13367 24790 13423 24846
rect 13491 24790 13547 24846
rect 13615 24790 13671 24846
rect 13739 24790 13795 24846
rect 13863 24790 13919 24846
rect 13987 24790 14043 24846
rect 14111 24790 14167 24846
rect 14235 24790 14291 24846
rect 14359 24790 14415 24846
rect 14483 24790 14539 24846
rect 14607 24790 14663 24846
rect 12871 24666 12927 24722
rect 12995 24666 13051 24722
rect 13119 24666 13175 24722
rect 13243 24666 13299 24722
rect 13367 24666 13423 24722
rect 13491 24666 13547 24722
rect 13615 24666 13671 24722
rect 13739 24666 13795 24722
rect 13863 24666 13919 24722
rect 13987 24666 14043 24722
rect 14111 24666 14167 24722
rect 14235 24666 14291 24722
rect 14359 24666 14415 24722
rect 14483 24666 14539 24722
rect 14607 24666 14663 24722
rect 12871 24542 12927 24598
rect 12995 24542 13051 24598
rect 13119 24542 13175 24598
rect 13243 24542 13299 24598
rect 13367 24542 13423 24598
rect 13491 24542 13547 24598
rect 13615 24542 13671 24598
rect 13739 24542 13795 24598
rect 13863 24542 13919 24598
rect 13987 24542 14043 24598
rect 14111 24542 14167 24598
rect 14235 24542 14291 24598
rect 14359 24542 14415 24598
rect 14483 24542 14539 24598
rect 14607 24542 14663 24598
rect 12871 24418 12927 24474
rect 12995 24418 13051 24474
rect 13119 24418 13175 24474
rect 13243 24418 13299 24474
rect 13367 24418 13423 24474
rect 13491 24418 13547 24474
rect 13615 24418 13671 24474
rect 13739 24418 13795 24474
rect 13863 24418 13919 24474
rect 13987 24418 14043 24474
rect 14111 24418 14167 24474
rect 14235 24418 14291 24474
rect 14359 24418 14415 24474
rect 14483 24418 14539 24474
rect 14607 24418 14663 24474
rect 12871 24294 12927 24350
rect 12995 24294 13051 24350
rect 13119 24294 13175 24350
rect 13243 24294 13299 24350
rect 13367 24294 13423 24350
rect 13491 24294 13547 24350
rect 13615 24294 13671 24350
rect 13739 24294 13795 24350
rect 13863 24294 13919 24350
rect 13987 24294 14043 24350
rect 14111 24294 14167 24350
rect 14235 24294 14291 24350
rect 14359 24294 14415 24350
rect 14483 24294 14539 24350
rect 14607 24294 14663 24350
rect 12871 24170 12927 24226
rect 12995 24170 13051 24226
rect 13119 24170 13175 24226
rect 13243 24170 13299 24226
rect 13367 24170 13423 24226
rect 13491 24170 13547 24226
rect 13615 24170 13671 24226
rect 13739 24170 13795 24226
rect 13863 24170 13919 24226
rect 13987 24170 14043 24226
rect 14111 24170 14167 24226
rect 14235 24170 14291 24226
rect 14359 24170 14415 24226
rect 14483 24170 14539 24226
rect 14607 24170 14663 24226
rect 12871 24046 12927 24102
rect 12995 24046 13051 24102
rect 13119 24046 13175 24102
rect 13243 24046 13299 24102
rect 13367 24046 13423 24102
rect 13491 24046 13547 24102
rect 13615 24046 13671 24102
rect 13739 24046 13795 24102
rect 13863 24046 13919 24102
rect 13987 24046 14043 24102
rect 14111 24046 14167 24102
rect 14235 24046 14291 24102
rect 14359 24046 14415 24102
rect 14483 24046 14539 24102
rect 14607 24046 14663 24102
rect 315 23698 371 23754
rect 439 23698 495 23754
rect 563 23698 619 23754
rect 687 23698 743 23754
rect 811 23698 867 23754
rect 935 23698 991 23754
rect 1059 23698 1115 23754
rect 1183 23698 1239 23754
rect 1307 23698 1363 23754
rect 1431 23698 1487 23754
rect 1555 23698 1611 23754
rect 1679 23698 1735 23754
rect 1803 23698 1859 23754
rect 1927 23698 1983 23754
rect 2051 23698 2107 23754
rect 315 23574 371 23630
rect 439 23574 495 23630
rect 563 23574 619 23630
rect 687 23574 743 23630
rect 811 23574 867 23630
rect 935 23574 991 23630
rect 1059 23574 1115 23630
rect 1183 23574 1239 23630
rect 1307 23574 1363 23630
rect 1431 23574 1487 23630
rect 1555 23574 1611 23630
rect 1679 23574 1735 23630
rect 1803 23574 1859 23630
rect 1927 23574 1983 23630
rect 2051 23574 2107 23630
rect 315 23450 371 23506
rect 439 23450 495 23506
rect 563 23450 619 23506
rect 687 23450 743 23506
rect 811 23450 867 23506
rect 935 23450 991 23506
rect 1059 23450 1115 23506
rect 1183 23450 1239 23506
rect 1307 23450 1363 23506
rect 1431 23450 1487 23506
rect 1555 23450 1611 23506
rect 1679 23450 1735 23506
rect 1803 23450 1859 23506
rect 1927 23450 1983 23506
rect 2051 23450 2107 23506
rect 315 23326 371 23382
rect 439 23326 495 23382
rect 563 23326 619 23382
rect 687 23326 743 23382
rect 811 23326 867 23382
rect 935 23326 991 23382
rect 1059 23326 1115 23382
rect 1183 23326 1239 23382
rect 1307 23326 1363 23382
rect 1431 23326 1487 23382
rect 1555 23326 1611 23382
rect 1679 23326 1735 23382
rect 1803 23326 1859 23382
rect 1927 23326 1983 23382
rect 2051 23326 2107 23382
rect 315 23202 371 23258
rect 439 23202 495 23258
rect 563 23202 619 23258
rect 687 23202 743 23258
rect 811 23202 867 23258
rect 935 23202 991 23258
rect 1059 23202 1115 23258
rect 1183 23202 1239 23258
rect 1307 23202 1363 23258
rect 1431 23202 1487 23258
rect 1555 23202 1611 23258
rect 1679 23202 1735 23258
rect 1803 23202 1859 23258
rect 1927 23202 1983 23258
rect 2051 23202 2107 23258
rect 315 23078 371 23134
rect 439 23078 495 23134
rect 563 23078 619 23134
rect 687 23078 743 23134
rect 811 23078 867 23134
rect 935 23078 991 23134
rect 1059 23078 1115 23134
rect 1183 23078 1239 23134
rect 1307 23078 1363 23134
rect 1431 23078 1487 23134
rect 1555 23078 1611 23134
rect 1679 23078 1735 23134
rect 1803 23078 1859 23134
rect 1927 23078 1983 23134
rect 2051 23078 2107 23134
rect 315 22954 371 23010
rect 439 22954 495 23010
rect 563 22954 619 23010
rect 687 22954 743 23010
rect 811 22954 867 23010
rect 935 22954 991 23010
rect 1059 22954 1115 23010
rect 1183 22954 1239 23010
rect 1307 22954 1363 23010
rect 1431 22954 1487 23010
rect 1555 22954 1611 23010
rect 1679 22954 1735 23010
rect 1803 22954 1859 23010
rect 1927 22954 1983 23010
rect 2051 22954 2107 23010
rect 315 22830 371 22886
rect 439 22830 495 22886
rect 563 22830 619 22886
rect 687 22830 743 22886
rect 811 22830 867 22886
rect 935 22830 991 22886
rect 1059 22830 1115 22886
rect 1183 22830 1239 22886
rect 1307 22830 1363 22886
rect 1431 22830 1487 22886
rect 1555 22830 1611 22886
rect 1679 22830 1735 22886
rect 1803 22830 1859 22886
rect 1927 22830 1983 22886
rect 2051 22830 2107 22886
rect 315 22706 371 22762
rect 439 22706 495 22762
rect 563 22706 619 22762
rect 687 22706 743 22762
rect 811 22706 867 22762
rect 935 22706 991 22762
rect 1059 22706 1115 22762
rect 1183 22706 1239 22762
rect 1307 22706 1363 22762
rect 1431 22706 1487 22762
rect 1555 22706 1611 22762
rect 1679 22706 1735 22762
rect 1803 22706 1859 22762
rect 1927 22706 1983 22762
rect 2051 22706 2107 22762
rect 315 22582 371 22638
rect 439 22582 495 22638
rect 563 22582 619 22638
rect 687 22582 743 22638
rect 811 22582 867 22638
rect 935 22582 991 22638
rect 1059 22582 1115 22638
rect 1183 22582 1239 22638
rect 1307 22582 1363 22638
rect 1431 22582 1487 22638
rect 1555 22582 1611 22638
rect 1679 22582 1735 22638
rect 1803 22582 1859 22638
rect 1927 22582 1983 22638
rect 2051 22582 2107 22638
rect 315 22458 371 22514
rect 439 22458 495 22514
rect 563 22458 619 22514
rect 687 22458 743 22514
rect 811 22458 867 22514
rect 935 22458 991 22514
rect 1059 22458 1115 22514
rect 1183 22458 1239 22514
rect 1307 22458 1363 22514
rect 1431 22458 1487 22514
rect 1555 22458 1611 22514
rect 1679 22458 1735 22514
rect 1803 22458 1859 22514
rect 1927 22458 1983 22514
rect 2051 22458 2107 22514
rect 315 22334 371 22390
rect 439 22334 495 22390
rect 563 22334 619 22390
rect 687 22334 743 22390
rect 811 22334 867 22390
rect 935 22334 991 22390
rect 1059 22334 1115 22390
rect 1183 22334 1239 22390
rect 1307 22334 1363 22390
rect 1431 22334 1487 22390
rect 1555 22334 1611 22390
rect 1679 22334 1735 22390
rect 1803 22334 1859 22390
rect 1927 22334 1983 22390
rect 2051 22334 2107 22390
rect 315 22210 371 22266
rect 439 22210 495 22266
rect 563 22210 619 22266
rect 687 22210 743 22266
rect 811 22210 867 22266
rect 935 22210 991 22266
rect 1059 22210 1115 22266
rect 1183 22210 1239 22266
rect 1307 22210 1363 22266
rect 1431 22210 1487 22266
rect 1555 22210 1611 22266
rect 1679 22210 1735 22266
rect 1803 22210 1859 22266
rect 1927 22210 1983 22266
rect 2051 22210 2107 22266
rect 315 22086 371 22142
rect 439 22086 495 22142
rect 563 22086 619 22142
rect 687 22086 743 22142
rect 811 22086 867 22142
rect 935 22086 991 22142
rect 1059 22086 1115 22142
rect 1183 22086 1239 22142
rect 1307 22086 1363 22142
rect 1431 22086 1487 22142
rect 1555 22086 1611 22142
rect 1679 22086 1735 22142
rect 1803 22086 1859 22142
rect 1927 22086 1983 22142
rect 2051 22086 2107 22142
rect 315 21962 371 22018
rect 439 21962 495 22018
rect 563 21962 619 22018
rect 687 21962 743 22018
rect 811 21962 867 22018
rect 935 21962 991 22018
rect 1059 21962 1115 22018
rect 1183 21962 1239 22018
rect 1307 21962 1363 22018
rect 1431 21962 1487 22018
rect 1555 21962 1611 22018
rect 1679 21962 1735 22018
rect 1803 21962 1859 22018
rect 1927 21962 1983 22018
rect 2051 21962 2107 22018
rect 315 21838 371 21894
rect 439 21838 495 21894
rect 563 21838 619 21894
rect 687 21838 743 21894
rect 811 21838 867 21894
rect 935 21838 991 21894
rect 1059 21838 1115 21894
rect 1183 21838 1239 21894
rect 1307 21838 1363 21894
rect 1431 21838 1487 21894
rect 1555 21838 1611 21894
rect 1679 21838 1735 21894
rect 1803 21838 1859 21894
rect 1927 21838 1983 21894
rect 2051 21838 2107 21894
rect 315 21714 371 21770
rect 439 21714 495 21770
rect 563 21714 619 21770
rect 687 21714 743 21770
rect 811 21714 867 21770
rect 935 21714 991 21770
rect 1059 21714 1115 21770
rect 1183 21714 1239 21770
rect 1307 21714 1363 21770
rect 1431 21714 1487 21770
rect 1555 21714 1611 21770
rect 1679 21714 1735 21770
rect 1803 21714 1859 21770
rect 1927 21714 1983 21770
rect 2051 21714 2107 21770
rect 315 21590 371 21646
rect 439 21590 495 21646
rect 563 21590 619 21646
rect 687 21590 743 21646
rect 811 21590 867 21646
rect 935 21590 991 21646
rect 1059 21590 1115 21646
rect 1183 21590 1239 21646
rect 1307 21590 1363 21646
rect 1431 21590 1487 21646
rect 1555 21590 1611 21646
rect 1679 21590 1735 21646
rect 1803 21590 1859 21646
rect 1927 21590 1983 21646
rect 2051 21590 2107 21646
rect 315 21466 371 21522
rect 439 21466 495 21522
rect 563 21466 619 21522
rect 687 21466 743 21522
rect 811 21466 867 21522
rect 935 21466 991 21522
rect 1059 21466 1115 21522
rect 1183 21466 1239 21522
rect 1307 21466 1363 21522
rect 1431 21466 1487 21522
rect 1555 21466 1611 21522
rect 1679 21466 1735 21522
rect 1803 21466 1859 21522
rect 1927 21466 1983 21522
rect 2051 21466 2107 21522
rect 315 21342 371 21398
rect 439 21342 495 21398
rect 563 21342 619 21398
rect 687 21342 743 21398
rect 811 21342 867 21398
rect 935 21342 991 21398
rect 1059 21342 1115 21398
rect 1183 21342 1239 21398
rect 1307 21342 1363 21398
rect 1431 21342 1487 21398
rect 1555 21342 1611 21398
rect 1679 21342 1735 21398
rect 1803 21342 1859 21398
rect 1927 21342 1983 21398
rect 2051 21342 2107 21398
rect 315 21218 371 21274
rect 439 21218 495 21274
rect 563 21218 619 21274
rect 687 21218 743 21274
rect 811 21218 867 21274
rect 935 21218 991 21274
rect 1059 21218 1115 21274
rect 1183 21218 1239 21274
rect 1307 21218 1363 21274
rect 1431 21218 1487 21274
rect 1555 21218 1611 21274
rect 1679 21218 1735 21274
rect 1803 21218 1859 21274
rect 1927 21218 1983 21274
rect 2051 21218 2107 21274
rect 315 21094 371 21150
rect 439 21094 495 21150
rect 563 21094 619 21150
rect 687 21094 743 21150
rect 811 21094 867 21150
rect 935 21094 991 21150
rect 1059 21094 1115 21150
rect 1183 21094 1239 21150
rect 1307 21094 1363 21150
rect 1431 21094 1487 21150
rect 1555 21094 1611 21150
rect 1679 21094 1735 21150
rect 1803 21094 1859 21150
rect 1927 21094 1983 21150
rect 2051 21094 2107 21150
rect 315 20970 371 21026
rect 439 20970 495 21026
rect 563 20970 619 21026
rect 687 20970 743 21026
rect 811 20970 867 21026
rect 935 20970 991 21026
rect 1059 20970 1115 21026
rect 1183 20970 1239 21026
rect 1307 20970 1363 21026
rect 1431 20970 1487 21026
rect 1555 20970 1611 21026
rect 1679 20970 1735 21026
rect 1803 20970 1859 21026
rect 1927 20970 1983 21026
rect 2051 20970 2107 21026
rect 315 20846 371 20902
rect 439 20846 495 20902
rect 563 20846 619 20902
rect 687 20846 743 20902
rect 811 20846 867 20902
rect 935 20846 991 20902
rect 1059 20846 1115 20902
rect 1183 20846 1239 20902
rect 1307 20846 1363 20902
rect 1431 20846 1487 20902
rect 1555 20846 1611 20902
rect 1679 20846 1735 20902
rect 1803 20846 1859 20902
rect 1927 20846 1983 20902
rect 2051 20846 2107 20902
rect 2808 23698 2864 23754
rect 2932 23698 2988 23754
rect 3056 23698 3112 23754
rect 3180 23698 3236 23754
rect 3304 23698 3360 23754
rect 3428 23698 3484 23754
rect 3552 23698 3608 23754
rect 3676 23698 3732 23754
rect 3800 23698 3856 23754
rect 3924 23698 3980 23754
rect 4048 23698 4104 23754
rect 4172 23698 4228 23754
rect 4296 23698 4352 23754
rect 4420 23698 4476 23754
rect 4544 23698 4600 23754
rect 4668 23698 4724 23754
rect 2808 23574 2864 23630
rect 2932 23574 2988 23630
rect 3056 23574 3112 23630
rect 3180 23574 3236 23630
rect 3304 23574 3360 23630
rect 3428 23574 3484 23630
rect 3552 23574 3608 23630
rect 3676 23574 3732 23630
rect 3800 23574 3856 23630
rect 3924 23574 3980 23630
rect 4048 23574 4104 23630
rect 4172 23574 4228 23630
rect 4296 23574 4352 23630
rect 4420 23574 4476 23630
rect 4544 23574 4600 23630
rect 4668 23574 4724 23630
rect 2808 23450 2864 23506
rect 2932 23450 2988 23506
rect 3056 23450 3112 23506
rect 3180 23450 3236 23506
rect 3304 23450 3360 23506
rect 3428 23450 3484 23506
rect 3552 23450 3608 23506
rect 3676 23450 3732 23506
rect 3800 23450 3856 23506
rect 3924 23450 3980 23506
rect 4048 23450 4104 23506
rect 4172 23450 4228 23506
rect 4296 23450 4352 23506
rect 4420 23450 4476 23506
rect 4544 23450 4600 23506
rect 4668 23450 4724 23506
rect 2808 23326 2864 23382
rect 2932 23326 2988 23382
rect 3056 23326 3112 23382
rect 3180 23326 3236 23382
rect 3304 23326 3360 23382
rect 3428 23326 3484 23382
rect 3552 23326 3608 23382
rect 3676 23326 3732 23382
rect 3800 23326 3856 23382
rect 3924 23326 3980 23382
rect 4048 23326 4104 23382
rect 4172 23326 4228 23382
rect 4296 23326 4352 23382
rect 4420 23326 4476 23382
rect 4544 23326 4600 23382
rect 4668 23326 4724 23382
rect 2808 23202 2864 23258
rect 2932 23202 2988 23258
rect 3056 23202 3112 23258
rect 3180 23202 3236 23258
rect 3304 23202 3360 23258
rect 3428 23202 3484 23258
rect 3552 23202 3608 23258
rect 3676 23202 3732 23258
rect 3800 23202 3856 23258
rect 3924 23202 3980 23258
rect 4048 23202 4104 23258
rect 4172 23202 4228 23258
rect 4296 23202 4352 23258
rect 4420 23202 4476 23258
rect 4544 23202 4600 23258
rect 4668 23202 4724 23258
rect 2808 23078 2864 23134
rect 2932 23078 2988 23134
rect 3056 23078 3112 23134
rect 3180 23078 3236 23134
rect 3304 23078 3360 23134
rect 3428 23078 3484 23134
rect 3552 23078 3608 23134
rect 3676 23078 3732 23134
rect 3800 23078 3856 23134
rect 3924 23078 3980 23134
rect 4048 23078 4104 23134
rect 4172 23078 4228 23134
rect 4296 23078 4352 23134
rect 4420 23078 4476 23134
rect 4544 23078 4600 23134
rect 4668 23078 4724 23134
rect 2808 22954 2864 23010
rect 2932 22954 2988 23010
rect 3056 22954 3112 23010
rect 3180 22954 3236 23010
rect 3304 22954 3360 23010
rect 3428 22954 3484 23010
rect 3552 22954 3608 23010
rect 3676 22954 3732 23010
rect 3800 22954 3856 23010
rect 3924 22954 3980 23010
rect 4048 22954 4104 23010
rect 4172 22954 4228 23010
rect 4296 22954 4352 23010
rect 4420 22954 4476 23010
rect 4544 22954 4600 23010
rect 4668 22954 4724 23010
rect 2808 22830 2864 22886
rect 2932 22830 2988 22886
rect 3056 22830 3112 22886
rect 3180 22830 3236 22886
rect 3304 22830 3360 22886
rect 3428 22830 3484 22886
rect 3552 22830 3608 22886
rect 3676 22830 3732 22886
rect 3800 22830 3856 22886
rect 3924 22830 3980 22886
rect 4048 22830 4104 22886
rect 4172 22830 4228 22886
rect 4296 22830 4352 22886
rect 4420 22830 4476 22886
rect 4544 22830 4600 22886
rect 4668 22830 4724 22886
rect 2808 22706 2864 22762
rect 2932 22706 2988 22762
rect 3056 22706 3112 22762
rect 3180 22706 3236 22762
rect 3304 22706 3360 22762
rect 3428 22706 3484 22762
rect 3552 22706 3608 22762
rect 3676 22706 3732 22762
rect 3800 22706 3856 22762
rect 3924 22706 3980 22762
rect 4048 22706 4104 22762
rect 4172 22706 4228 22762
rect 4296 22706 4352 22762
rect 4420 22706 4476 22762
rect 4544 22706 4600 22762
rect 4668 22706 4724 22762
rect 2808 22582 2864 22638
rect 2932 22582 2988 22638
rect 3056 22582 3112 22638
rect 3180 22582 3236 22638
rect 3304 22582 3360 22638
rect 3428 22582 3484 22638
rect 3552 22582 3608 22638
rect 3676 22582 3732 22638
rect 3800 22582 3856 22638
rect 3924 22582 3980 22638
rect 4048 22582 4104 22638
rect 4172 22582 4228 22638
rect 4296 22582 4352 22638
rect 4420 22582 4476 22638
rect 4544 22582 4600 22638
rect 4668 22582 4724 22638
rect 2808 22458 2864 22514
rect 2932 22458 2988 22514
rect 3056 22458 3112 22514
rect 3180 22458 3236 22514
rect 3304 22458 3360 22514
rect 3428 22458 3484 22514
rect 3552 22458 3608 22514
rect 3676 22458 3732 22514
rect 3800 22458 3856 22514
rect 3924 22458 3980 22514
rect 4048 22458 4104 22514
rect 4172 22458 4228 22514
rect 4296 22458 4352 22514
rect 4420 22458 4476 22514
rect 4544 22458 4600 22514
rect 4668 22458 4724 22514
rect 2808 22334 2864 22390
rect 2932 22334 2988 22390
rect 3056 22334 3112 22390
rect 3180 22334 3236 22390
rect 3304 22334 3360 22390
rect 3428 22334 3484 22390
rect 3552 22334 3608 22390
rect 3676 22334 3732 22390
rect 3800 22334 3856 22390
rect 3924 22334 3980 22390
rect 4048 22334 4104 22390
rect 4172 22334 4228 22390
rect 4296 22334 4352 22390
rect 4420 22334 4476 22390
rect 4544 22334 4600 22390
rect 4668 22334 4724 22390
rect 2808 22210 2864 22266
rect 2932 22210 2988 22266
rect 3056 22210 3112 22266
rect 3180 22210 3236 22266
rect 3304 22210 3360 22266
rect 3428 22210 3484 22266
rect 3552 22210 3608 22266
rect 3676 22210 3732 22266
rect 3800 22210 3856 22266
rect 3924 22210 3980 22266
rect 4048 22210 4104 22266
rect 4172 22210 4228 22266
rect 4296 22210 4352 22266
rect 4420 22210 4476 22266
rect 4544 22210 4600 22266
rect 4668 22210 4724 22266
rect 2808 22086 2864 22142
rect 2932 22086 2988 22142
rect 3056 22086 3112 22142
rect 3180 22086 3236 22142
rect 3304 22086 3360 22142
rect 3428 22086 3484 22142
rect 3552 22086 3608 22142
rect 3676 22086 3732 22142
rect 3800 22086 3856 22142
rect 3924 22086 3980 22142
rect 4048 22086 4104 22142
rect 4172 22086 4228 22142
rect 4296 22086 4352 22142
rect 4420 22086 4476 22142
rect 4544 22086 4600 22142
rect 4668 22086 4724 22142
rect 2808 21962 2864 22018
rect 2932 21962 2988 22018
rect 3056 21962 3112 22018
rect 3180 21962 3236 22018
rect 3304 21962 3360 22018
rect 3428 21962 3484 22018
rect 3552 21962 3608 22018
rect 3676 21962 3732 22018
rect 3800 21962 3856 22018
rect 3924 21962 3980 22018
rect 4048 21962 4104 22018
rect 4172 21962 4228 22018
rect 4296 21962 4352 22018
rect 4420 21962 4476 22018
rect 4544 21962 4600 22018
rect 4668 21962 4724 22018
rect 2808 21838 2864 21894
rect 2932 21838 2988 21894
rect 3056 21838 3112 21894
rect 3180 21838 3236 21894
rect 3304 21838 3360 21894
rect 3428 21838 3484 21894
rect 3552 21838 3608 21894
rect 3676 21838 3732 21894
rect 3800 21838 3856 21894
rect 3924 21838 3980 21894
rect 4048 21838 4104 21894
rect 4172 21838 4228 21894
rect 4296 21838 4352 21894
rect 4420 21838 4476 21894
rect 4544 21838 4600 21894
rect 4668 21838 4724 21894
rect 2808 21714 2864 21770
rect 2932 21714 2988 21770
rect 3056 21714 3112 21770
rect 3180 21714 3236 21770
rect 3304 21714 3360 21770
rect 3428 21714 3484 21770
rect 3552 21714 3608 21770
rect 3676 21714 3732 21770
rect 3800 21714 3856 21770
rect 3924 21714 3980 21770
rect 4048 21714 4104 21770
rect 4172 21714 4228 21770
rect 4296 21714 4352 21770
rect 4420 21714 4476 21770
rect 4544 21714 4600 21770
rect 4668 21714 4724 21770
rect 2808 21590 2864 21646
rect 2932 21590 2988 21646
rect 3056 21590 3112 21646
rect 3180 21590 3236 21646
rect 3304 21590 3360 21646
rect 3428 21590 3484 21646
rect 3552 21590 3608 21646
rect 3676 21590 3732 21646
rect 3800 21590 3856 21646
rect 3924 21590 3980 21646
rect 4048 21590 4104 21646
rect 4172 21590 4228 21646
rect 4296 21590 4352 21646
rect 4420 21590 4476 21646
rect 4544 21590 4600 21646
rect 4668 21590 4724 21646
rect 2808 21466 2864 21522
rect 2932 21466 2988 21522
rect 3056 21466 3112 21522
rect 3180 21466 3236 21522
rect 3304 21466 3360 21522
rect 3428 21466 3484 21522
rect 3552 21466 3608 21522
rect 3676 21466 3732 21522
rect 3800 21466 3856 21522
rect 3924 21466 3980 21522
rect 4048 21466 4104 21522
rect 4172 21466 4228 21522
rect 4296 21466 4352 21522
rect 4420 21466 4476 21522
rect 4544 21466 4600 21522
rect 4668 21466 4724 21522
rect 2808 21342 2864 21398
rect 2932 21342 2988 21398
rect 3056 21342 3112 21398
rect 3180 21342 3236 21398
rect 3304 21342 3360 21398
rect 3428 21342 3484 21398
rect 3552 21342 3608 21398
rect 3676 21342 3732 21398
rect 3800 21342 3856 21398
rect 3924 21342 3980 21398
rect 4048 21342 4104 21398
rect 4172 21342 4228 21398
rect 4296 21342 4352 21398
rect 4420 21342 4476 21398
rect 4544 21342 4600 21398
rect 4668 21342 4724 21398
rect 2808 21218 2864 21274
rect 2932 21218 2988 21274
rect 3056 21218 3112 21274
rect 3180 21218 3236 21274
rect 3304 21218 3360 21274
rect 3428 21218 3484 21274
rect 3552 21218 3608 21274
rect 3676 21218 3732 21274
rect 3800 21218 3856 21274
rect 3924 21218 3980 21274
rect 4048 21218 4104 21274
rect 4172 21218 4228 21274
rect 4296 21218 4352 21274
rect 4420 21218 4476 21274
rect 4544 21218 4600 21274
rect 4668 21218 4724 21274
rect 2808 21094 2864 21150
rect 2932 21094 2988 21150
rect 3056 21094 3112 21150
rect 3180 21094 3236 21150
rect 3304 21094 3360 21150
rect 3428 21094 3484 21150
rect 3552 21094 3608 21150
rect 3676 21094 3732 21150
rect 3800 21094 3856 21150
rect 3924 21094 3980 21150
rect 4048 21094 4104 21150
rect 4172 21094 4228 21150
rect 4296 21094 4352 21150
rect 4420 21094 4476 21150
rect 4544 21094 4600 21150
rect 4668 21094 4724 21150
rect 2808 20970 2864 21026
rect 2932 20970 2988 21026
rect 3056 20970 3112 21026
rect 3180 20970 3236 21026
rect 3304 20970 3360 21026
rect 3428 20970 3484 21026
rect 3552 20970 3608 21026
rect 3676 20970 3732 21026
rect 3800 20970 3856 21026
rect 3924 20970 3980 21026
rect 4048 20970 4104 21026
rect 4172 20970 4228 21026
rect 4296 20970 4352 21026
rect 4420 20970 4476 21026
rect 4544 20970 4600 21026
rect 4668 20970 4724 21026
rect 2808 20846 2864 20902
rect 2932 20846 2988 20902
rect 3056 20846 3112 20902
rect 3180 20846 3236 20902
rect 3304 20846 3360 20902
rect 3428 20846 3484 20902
rect 3552 20846 3608 20902
rect 3676 20846 3732 20902
rect 3800 20846 3856 20902
rect 3924 20846 3980 20902
rect 4048 20846 4104 20902
rect 4172 20846 4228 20902
rect 4296 20846 4352 20902
rect 4420 20846 4476 20902
rect 4544 20846 4600 20902
rect 4668 20846 4724 20902
rect 5178 23698 5234 23754
rect 5302 23698 5358 23754
rect 5426 23698 5482 23754
rect 5550 23698 5606 23754
rect 5674 23698 5730 23754
rect 5798 23698 5854 23754
rect 5922 23698 5978 23754
rect 6046 23698 6102 23754
rect 6170 23698 6226 23754
rect 6294 23698 6350 23754
rect 6418 23698 6474 23754
rect 6542 23698 6598 23754
rect 6666 23698 6722 23754
rect 6790 23698 6846 23754
rect 6914 23698 6970 23754
rect 7038 23698 7094 23754
rect 5178 23574 5234 23630
rect 5302 23574 5358 23630
rect 5426 23574 5482 23630
rect 5550 23574 5606 23630
rect 5674 23574 5730 23630
rect 5798 23574 5854 23630
rect 5922 23574 5978 23630
rect 6046 23574 6102 23630
rect 6170 23574 6226 23630
rect 6294 23574 6350 23630
rect 6418 23574 6474 23630
rect 6542 23574 6598 23630
rect 6666 23574 6722 23630
rect 6790 23574 6846 23630
rect 6914 23574 6970 23630
rect 7038 23574 7094 23630
rect 5178 23450 5234 23506
rect 5302 23450 5358 23506
rect 5426 23450 5482 23506
rect 5550 23450 5606 23506
rect 5674 23450 5730 23506
rect 5798 23450 5854 23506
rect 5922 23450 5978 23506
rect 6046 23450 6102 23506
rect 6170 23450 6226 23506
rect 6294 23450 6350 23506
rect 6418 23450 6474 23506
rect 6542 23450 6598 23506
rect 6666 23450 6722 23506
rect 6790 23450 6846 23506
rect 6914 23450 6970 23506
rect 7038 23450 7094 23506
rect 5178 23326 5234 23382
rect 5302 23326 5358 23382
rect 5426 23326 5482 23382
rect 5550 23326 5606 23382
rect 5674 23326 5730 23382
rect 5798 23326 5854 23382
rect 5922 23326 5978 23382
rect 6046 23326 6102 23382
rect 6170 23326 6226 23382
rect 6294 23326 6350 23382
rect 6418 23326 6474 23382
rect 6542 23326 6598 23382
rect 6666 23326 6722 23382
rect 6790 23326 6846 23382
rect 6914 23326 6970 23382
rect 7038 23326 7094 23382
rect 5178 23202 5234 23258
rect 5302 23202 5358 23258
rect 5426 23202 5482 23258
rect 5550 23202 5606 23258
rect 5674 23202 5730 23258
rect 5798 23202 5854 23258
rect 5922 23202 5978 23258
rect 6046 23202 6102 23258
rect 6170 23202 6226 23258
rect 6294 23202 6350 23258
rect 6418 23202 6474 23258
rect 6542 23202 6598 23258
rect 6666 23202 6722 23258
rect 6790 23202 6846 23258
rect 6914 23202 6970 23258
rect 7038 23202 7094 23258
rect 5178 23078 5234 23134
rect 5302 23078 5358 23134
rect 5426 23078 5482 23134
rect 5550 23078 5606 23134
rect 5674 23078 5730 23134
rect 5798 23078 5854 23134
rect 5922 23078 5978 23134
rect 6046 23078 6102 23134
rect 6170 23078 6226 23134
rect 6294 23078 6350 23134
rect 6418 23078 6474 23134
rect 6542 23078 6598 23134
rect 6666 23078 6722 23134
rect 6790 23078 6846 23134
rect 6914 23078 6970 23134
rect 7038 23078 7094 23134
rect 5178 22954 5234 23010
rect 5302 22954 5358 23010
rect 5426 22954 5482 23010
rect 5550 22954 5606 23010
rect 5674 22954 5730 23010
rect 5798 22954 5854 23010
rect 5922 22954 5978 23010
rect 6046 22954 6102 23010
rect 6170 22954 6226 23010
rect 6294 22954 6350 23010
rect 6418 22954 6474 23010
rect 6542 22954 6598 23010
rect 6666 22954 6722 23010
rect 6790 22954 6846 23010
rect 6914 22954 6970 23010
rect 7038 22954 7094 23010
rect 5178 22830 5234 22886
rect 5302 22830 5358 22886
rect 5426 22830 5482 22886
rect 5550 22830 5606 22886
rect 5674 22830 5730 22886
rect 5798 22830 5854 22886
rect 5922 22830 5978 22886
rect 6046 22830 6102 22886
rect 6170 22830 6226 22886
rect 6294 22830 6350 22886
rect 6418 22830 6474 22886
rect 6542 22830 6598 22886
rect 6666 22830 6722 22886
rect 6790 22830 6846 22886
rect 6914 22830 6970 22886
rect 7038 22830 7094 22886
rect 5178 22706 5234 22762
rect 5302 22706 5358 22762
rect 5426 22706 5482 22762
rect 5550 22706 5606 22762
rect 5674 22706 5730 22762
rect 5798 22706 5854 22762
rect 5922 22706 5978 22762
rect 6046 22706 6102 22762
rect 6170 22706 6226 22762
rect 6294 22706 6350 22762
rect 6418 22706 6474 22762
rect 6542 22706 6598 22762
rect 6666 22706 6722 22762
rect 6790 22706 6846 22762
rect 6914 22706 6970 22762
rect 7038 22706 7094 22762
rect 5178 22582 5234 22638
rect 5302 22582 5358 22638
rect 5426 22582 5482 22638
rect 5550 22582 5606 22638
rect 5674 22582 5730 22638
rect 5798 22582 5854 22638
rect 5922 22582 5978 22638
rect 6046 22582 6102 22638
rect 6170 22582 6226 22638
rect 6294 22582 6350 22638
rect 6418 22582 6474 22638
rect 6542 22582 6598 22638
rect 6666 22582 6722 22638
rect 6790 22582 6846 22638
rect 6914 22582 6970 22638
rect 7038 22582 7094 22638
rect 5178 22458 5234 22514
rect 5302 22458 5358 22514
rect 5426 22458 5482 22514
rect 5550 22458 5606 22514
rect 5674 22458 5730 22514
rect 5798 22458 5854 22514
rect 5922 22458 5978 22514
rect 6046 22458 6102 22514
rect 6170 22458 6226 22514
rect 6294 22458 6350 22514
rect 6418 22458 6474 22514
rect 6542 22458 6598 22514
rect 6666 22458 6722 22514
rect 6790 22458 6846 22514
rect 6914 22458 6970 22514
rect 7038 22458 7094 22514
rect 5178 22334 5234 22390
rect 5302 22334 5358 22390
rect 5426 22334 5482 22390
rect 5550 22334 5606 22390
rect 5674 22334 5730 22390
rect 5798 22334 5854 22390
rect 5922 22334 5978 22390
rect 6046 22334 6102 22390
rect 6170 22334 6226 22390
rect 6294 22334 6350 22390
rect 6418 22334 6474 22390
rect 6542 22334 6598 22390
rect 6666 22334 6722 22390
rect 6790 22334 6846 22390
rect 6914 22334 6970 22390
rect 7038 22334 7094 22390
rect 5178 22210 5234 22266
rect 5302 22210 5358 22266
rect 5426 22210 5482 22266
rect 5550 22210 5606 22266
rect 5674 22210 5730 22266
rect 5798 22210 5854 22266
rect 5922 22210 5978 22266
rect 6046 22210 6102 22266
rect 6170 22210 6226 22266
rect 6294 22210 6350 22266
rect 6418 22210 6474 22266
rect 6542 22210 6598 22266
rect 6666 22210 6722 22266
rect 6790 22210 6846 22266
rect 6914 22210 6970 22266
rect 7038 22210 7094 22266
rect 5178 22086 5234 22142
rect 5302 22086 5358 22142
rect 5426 22086 5482 22142
rect 5550 22086 5606 22142
rect 5674 22086 5730 22142
rect 5798 22086 5854 22142
rect 5922 22086 5978 22142
rect 6046 22086 6102 22142
rect 6170 22086 6226 22142
rect 6294 22086 6350 22142
rect 6418 22086 6474 22142
rect 6542 22086 6598 22142
rect 6666 22086 6722 22142
rect 6790 22086 6846 22142
rect 6914 22086 6970 22142
rect 7038 22086 7094 22142
rect 5178 21962 5234 22018
rect 5302 21962 5358 22018
rect 5426 21962 5482 22018
rect 5550 21962 5606 22018
rect 5674 21962 5730 22018
rect 5798 21962 5854 22018
rect 5922 21962 5978 22018
rect 6046 21962 6102 22018
rect 6170 21962 6226 22018
rect 6294 21962 6350 22018
rect 6418 21962 6474 22018
rect 6542 21962 6598 22018
rect 6666 21962 6722 22018
rect 6790 21962 6846 22018
rect 6914 21962 6970 22018
rect 7038 21962 7094 22018
rect 5178 21838 5234 21894
rect 5302 21838 5358 21894
rect 5426 21838 5482 21894
rect 5550 21838 5606 21894
rect 5674 21838 5730 21894
rect 5798 21838 5854 21894
rect 5922 21838 5978 21894
rect 6046 21838 6102 21894
rect 6170 21838 6226 21894
rect 6294 21838 6350 21894
rect 6418 21838 6474 21894
rect 6542 21838 6598 21894
rect 6666 21838 6722 21894
rect 6790 21838 6846 21894
rect 6914 21838 6970 21894
rect 7038 21838 7094 21894
rect 5178 21714 5234 21770
rect 5302 21714 5358 21770
rect 5426 21714 5482 21770
rect 5550 21714 5606 21770
rect 5674 21714 5730 21770
rect 5798 21714 5854 21770
rect 5922 21714 5978 21770
rect 6046 21714 6102 21770
rect 6170 21714 6226 21770
rect 6294 21714 6350 21770
rect 6418 21714 6474 21770
rect 6542 21714 6598 21770
rect 6666 21714 6722 21770
rect 6790 21714 6846 21770
rect 6914 21714 6970 21770
rect 7038 21714 7094 21770
rect 5178 21590 5234 21646
rect 5302 21590 5358 21646
rect 5426 21590 5482 21646
rect 5550 21590 5606 21646
rect 5674 21590 5730 21646
rect 5798 21590 5854 21646
rect 5922 21590 5978 21646
rect 6046 21590 6102 21646
rect 6170 21590 6226 21646
rect 6294 21590 6350 21646
rect 6418 21590 6474 21646
rect 6542 21590 6598 21646
rect 6666 21590 6722 21646
rect 6790 21590 6846 21646
rect 6914 21590 6970 21646
rect 7038 21590 7094 21646
rect 5178 21466 5234 21522
rect 5302 21466 5358 21522
rect 5426 21466 5482 21522
rect 5550 21466 5606 21522
rect 5674 21466 5730 21522
rect 5798 21466 5854 21522
rect 5922 21466 5978 21522
rect 6046 21466 6102 21522
rect 6170 21466 6226 21522
rect 6294 21466 6350 21522
rect 6418 21466 6474 21522
rect 6542 21466 6598 21522
rect 6666 21466 6722 21522
rect 6790 21466 6846 21522
rect 6914 21466 6970 21522
rect 7038 21466 7094 21522
rect 5178 21342 5234 21398
rect 5302 21342 5358 21398
rect 5426 21342 5482 21398
rect 5550 21342 5606 21398
rect 5674 21342 5730 21398
rect 5798 21342 5854 21398
rect 5922 21342 5978 21398
rect 6046 21342 6102 21398
rect 6170 21342 6226 21398
rect 6294 21342 6350 21398
rect 6418 21342 6474 21398
rect 6542 21342 6598 21398
rect 6666 21342 6722 21398
rect 6790 21342 6846 21398
rect 6914 21342 6970 21398
rect 7038 21342 7094 21398
rect 5178 21218 5234 21274
rect 5302 21218 5358 21274
rect 5426 21218 5482 21274
rect 5550 21218 5606 21274
rect 5674 21218 5730 21274
rect 5798 21218 5854 21274
rect 5922 21218 5978 21274
rect 6046 21218 6102 21274
rect 6170 21218 6226 21274
rect 6294 21218 6350 21274
rect 6418 21218 6474 21274
rect 6542 21218 6598 21274
rect 6666 21218 6722 21274
rect 6790 21218 6846 21274
rect 6914 21218 6970 21274
rect 7038 21218 7094 21274
rect 5178 21094 5234 21150
rect 5302 21094 5358 21150
rect 5426 21094 5482 21150
rect 5550 21094 5606 21150
rect 5674 21094 5730 21150
rect 5798 21094 5854 21150
rect 5922 21094 5978 21150
rect 6046 21094 6102 21150
rect 6170 21094 6226 21150
rect 6294 21094 6350 21150
rect 6418 21094 6474 21150
rect 6542 21094 6598 21150
rect 6666 21094 6722 21150
rect 6790 21094 6846 21150
rect 6914 21094 6970 21150
rect 7038 21094 7094 21150
rect 5178 20970 5234 21026
rect 5302 20970 5358 21026
rect 5426 20970 5482 21026
rect 5550 20970 5606 21026
rect 5674 20970 5730 21026
rect 5798 20970 5854 21026
rect 5922 20970 5978 21026
rect 6046 20970 6102 21026
rect 6170 20970 6226 21026
rect 6294 20970 6350 21026
rect 6418 20970 6474 21026
rect 6542 20970 6598 21026
rect 6666 20970 6722 21026
rect 6790 20970 6846 21026
rect 6914 20970 6970 21026
rect 7038 20970 7094 21026
rect 5178 20846 5234 20902
rect 5302 20846 5358 20902
rect 5426 20846 5482 20902
rect 5550 20846 5606 20902
rect 5674 20846 5730 20902
rect 5798 20846 5854 20902
rect 5922 20846 5978 20902
rect 6046 20846 6102 20902
rect 6170 20846 6226 20902
rect 6294 20846 6350 20902
rect 6418 20846 6474 20902
rect 6542 20846 6598 20902
rect 6666 20846 6722 20902
rect 6790 20846 6846 20902
rect 6914 20846 6970 20902
rect 7038 20846 7094 20902
rect 7884 23698 7940 23754
rect 8008 23698 8064 23754
rect 8132 23698 8188 23754
rect 8256 23698 8312 23754
rect 8380 23698 8436 23754
rect 8504 23698 8560 23754
rect 8628 23698 8684 23754
rect 8752 23698 8808 23754
rect 8876 23698 8932 23754
rect 9000 23698 9056 23754
rect 9124 23698 9180 23754
rect 9248 23698 9304 23754
rect 9372 23698 9428 23754
rect 9496 23698 9552 23754
rect 9620 23698 9676 23754
rect 9744 23698 9800 23754
rect 7884 23574 7940 23630
rect 8008 23574 8064 23630
rect 8132 23574 8188 23630
rect 8256 23574 8312 23630
rect 8380 23574 8436 23630
rect 8504 23574 8560 23630
rect 8628 23574 8684 23630
rect 8752 23574 8808 23630
rect 8876 23574 8932 23630
rect 9000 23574 9056 23630
rect 9124 23574 9180 23630
rect 9248 23574 9304 23630
rect 9372 23574 9428 23630
rect 9496 23574 9552 23630
rect 9620 23574 9676 23630
rect 9744 23574 9800 23630
rect 7884 23450 7940 23506
rect 8008 23450 8064 23506
rect 8132 23450 8188 23506
rect 8256 23450 8312 23506
rect 8380 23450 8436 23506
rect 8504 23450 8560 23506
rect 8628 23450 8684 23506
rect 8752 23450 8808 23506
rect 8876 23450 8932 23506
rect 9000 23450 9056 23506
rect 9124 23450 9180 23506
rect 9248 23450 9304 23506
rect 9372 23450 9428 23506
rect 9496 23450 9552 23506
rect 9620 23450 9676 23506
rect 9744 23450 9800 23506
rect 7884 23326 7940 23382
rect 8008 23326 8064 23382
rect 8132 23326 8188 23382
rect 8256 23326 8312 23382
rect 8380 23326 8436 23382
rect 8504 23326 8560 23382
rect 8628 23326 8684 23382
rect 8752 23326 8808 23382
rect 8876 23326 8932 23382
rect 9000 23326 9056 23382
rect 9124 23326 9180 23382
rect 9248 23326 9304 23382
rect 9372 23326 9428 23382
rect 9496 23326 9552 23382
rect 9620 23326 9676 23382
rect 9744 23326 9800 23382
rect 7884 23202 7940 23258
rect 8008 23202 8064 23258
rect 8132 23202 8188 23258
rect 8256 23202 8312 23258
rect 8380 23202 8436 23258
rect 8504 23202 8560 23258
rect 8628 23202 8684 23258
rect 8752 23202 8808 23258
rect 8876 23202 8932 23258
rect 9000 23202 9056 23258
rect 9124 23202 9180 23258
rect 9248 23202 9304 23258
rect 9372 23202 9428 23258
rect 9496 23202 9552 23258
rect 9620 23202 9676 23258
rect 9744 23202 9800 23258
rect 7884 23078 7940 23134
rect 8008 23078 8064 23134
rect 8132 23078 8188 23134
rect 8256 23078 8312 23134
rect 8380 23078 8436 23134
rect 8504 23078 8560 23134
rect 8628 23078 8684 23134
rect 8752 23078 8808 23134
rect 8876 23078 8932 23134
rect 9000 23078 9056 23134
rect 9124 23078 9180 23134
rect 9248 23078 9304 23134
rect 9372 23078 9428 23134
rect 9496 23078 9552 23134
rect 9620 23078 9676 23134
rect 9744 23078 9800 23134
rect 7884 22954 7940 23010
rect 8008 22954 8064 23010
rect 8132 22954 8188 23010
rect 8256 22954 8312 23010
rect 8380 22954 8436 23010
rect 8504 22954 8560 23010
rect 8628 22954 8684 23010
rect 8752 22954 8808 23010
rect 8876 22954 8932 23010
rect 9000 22954 9056 23010
rect 9124 22954 9180 23010
rect 9248 22954 9304 23010
rect 9372 22954 9428 23010
rect 9496 22954 9552 23010
rect 9620 22954 9676 23010
rect 9744 22954 9800 23010
rect 7884 22830 7940 22886
rect 8008 22830 8064 22886
rect 8132 22830 8188 22886
rect 8256 22830 8312 22886
rect 8380 22830 8436 22886
rect 8504 22830 8560 22886
rect 8628 22830 8684 22886
rect 8752 22830 8808 22886
rect 8876 22830 8932 22886
rect 9000 22830 9056 22886
rect 9124 22830 9180 22886
rect 9248 22830 9304 22886
rect 9372 22830 9428 22886
rect 9496 22830 9552 22886
rect 9620 22830 9676 22886
rect 9744 22830 9800 22886
rect 7884 22706 7940 22762
rect 8008 22706 8064 22762
rect 8132 22706 8188 22762
rect 8256 22706 8312 22762
rect 8380 22706 8436 22762
rect 8504 22706 8560 22762
rect 8628 22706 8684 22762
rect 8752 22706 8808 22762
rect 8876 22706 8932 22762
rect 9000 22706 9056 22762
rect 9124 22706 9180 22762
rect 9248 22706 9304 22762
rect 9372 22706 9428 22762
rect 9496 22706 9552 22762
rect 9620 22706 9676 22762
rect 9744 22706 9800 22762
rect 7884 22582 7940 22638
rect 8008 22582 8064 22638
rect 8132 22582 8188 22638
rect 8256 22582 8312 22638
rect 8380 22582 8436 22638
rect 8504 22582 8560 22638
rect 8628 22582 8684 22638
rect 8752 22582 8808 22638
rect 8876 22582 8932 22638
rect 9000 22582 9056 22638
rect 9124 22582 9180 22638
rect 9248 22582 9304 22638
rect 9372 22582 9428 22638
rect 9496 22582 9552 22638
rect 9620 22582 9676 22638
rect 9744 22582 9800 22638
rect 7884 22458 7940 22514
rect 8008 22458 8064 22514
rect 8132 22458 8188 22514
rect 8256 22458 8312 22514
rect 8380 22458 8436 22514
rect 8504 22458 8560 22514
rect 8628 22458 8684 22514
rect 8752 22458 8808 22514
rect 8876 22458 8932 22514
rect 9000 22458 9056 22514
rect 9124 22458 9180 22514
rect 9248 22458 9304 22514
rect 9372 22458 9428 22514
rect 9496 22458 9552 22514
rect 9620 22458 9676 22514
rect 9744 22458 9800 22514
rect 7884 22334 7940 22390
rect 8008 22334 8064 22390
rect 8132 22334 8188 22390
rect 8256 22334 8312 22390
rect 8380 22334 8436 22390
rect 8504 22334 8560 22390
rect 8628 22334 8684 22390
rect 8752 22334 8808 22390
rect 8876 22334 8932 22390
rect 9000 22334 9056 22390
rect 9124 22334 9180 22390
rect 9248 22334 9304 22390
rect 9372 22334 9428 22390
rect 9496 22334 9552 22390
rect 9620 22334 9676 22390
rect 9744 22334 9800 22390
rect 7884 22210 7940 22266
rect 8008 22210 8064 22266
rect 8132 22210 8188 22266
rect 8256 22210 8312 22266
rect 8380 22210 8436 22266
rect 8504 22210 8560 22266
rect 8628 22210 8684 22266
rect 8752 22210 8808 22266
rect 8876 22210 8932 22266
rect 9000 22210 9056 22266
rect 9124 22210 9180 22266
rect 9248 22210 9304 22266
rect 9372 22210 9428 22266
rect 9496 22210 9552 22266
rect 9620 22210 9676 22266
rect 9744 22210 9800 22266
rect 7884 22086 7940 22142
rect 8008 22086 8064 22142
rect 8132 22086 8188 22142
rect 8256 22086 8312 22142
rect 8380 22086 8436 22142
rect 8504 22086 8560 22142
rect 8628 22086 8684 22142
rect 8752 22086 8808 22142
rect 8876 22086 8932 22142
rect 9000 22086 9056 22142
rect 9124 22086 9180 22142
rect 9248 22086 9304 22142
rect 9372 22086 9428 22142
rect 9496 22086 9552 22142
rect 9620 22086 9676 22142
rect 9744 22086 9800 22142
rect 7884 21962 7940 22018
rect 8008 21962 8064 22018
rect 8132 21962 8188 22018
rect 8256 21962 8312 22018
rect 8380 21962 8436 22018
rect 8504 21962 8560 22018
rect 8628 21962 8684 22018
rect 8752 21962 8808 22018
rect 8876 21962 8932 22018
rect 9000 21962 9056 22018
rect 9124 21962 9180 22018
rect 9248 21962 9304 22018
rect 9372 21962 9428 22018
rect 9496 21962 9552 22018
rect 9620 21962 9676 22018
rect 9744 21962 9800 22018
rect 7884 21838 7940 21894
rect 8008 21838 8064 21894
rect 8132 21838 8188 21894
rect 8256 21838 8312 21894
rect 8380 21838 8436 21894
rect 8504 21838 8560 21894
rect 8628 21838 8684 21894
rect 8752 21838 8808 21894
rect 8876 21838 8932 21894
rect 9000 21838 9056 21894
rect 9124 21838 9180 21894
rect 9248 21838 9304 21894
rect 9372 21838 9428 21894
rect 9496 21838 9552 21894
rect 9620 21838 9676 21894
rect 9744 21838 9800 21894
rect 7884 21714 7940 21770
rect 8008 21714 8064 21770
rect 8132 21714 8188 21770
rect 8256 21714 8312 21770
rect 8380 21714 8436 21770
rect 8504 21714 8560 21770
rect 8628 21714 8684 21770
rect 8752 21714 8808 21770
rect 8876 21714 8932 21770
rect 9000 21714 9056 21770
rect 9124 21714 9180 21770
rect 9248 21714 9304 21770
rect 9372 21714 9428 21770
rect 9496 21714 9552 21770
rect 9620 21714 9676 21770
rect 9744 21714 9800 21770
rect 7884 21590 7940 21646
rect 8008 21590 8064 21646
rect 8132 21590 8188 21646
rect 8256 21590 8312 21646
rect 8380 21590 8436 21646
rect 8504 21590 8560 21646
rect 8628 21590 8684 21646
rect 8752 21590 8808 21646
rect 8876 21590 8932 21646
rect 9000 21590 9056 21646
rect 9124 21590 9180 21646
rect 9248 21590 9304 21646
rect 9372 21590 9428 21646
rect 9496 21590 9552 21646
rect 9620 21590 9676 21646
rect 9744 21590 9800 21646
rect 7884 21466 7940 21522
rect 8008 21466 8064 21522
rect 8132 21466 8188 21522
rect 8256 21466 8312 21522
rect 8380 21466 8436 21522
rect 8504 21466 8560 21522
rect 8628 21466 8684 21522
rect 8752 21466 8808 21522
rect 8876 21466 8932 21522
rect 9000 21466 9056 21522
rect 9124 21466 9180 21522
rect 9248 21466 9304 21522
rect 9372 21466 9428 21522
rect 9496 21466 9552 21522
rect 9620 21466 9676 21522
rect 9744 21466 9800 21522
rect 7884 21342 7940 21398
rect 8008 21342 8064 21398
rect 8132 21342 8188 21398
rect 8256 21342 8312 21398
rect 8380 21342 8436 21398
rect 8504 21342 8560 21398
rect 8628 21342 8684 21398
rect 8752 21342 8808 21398
rect 8876 21342 8932 21398
rect 9000 21342 9056 21398
rect 9124 21342 9180 21398
rect 9248 21342 9304 21398
rect 9372 21342 9428 21398
rect 9496 21342 9552 21398
rect 9620 21342 9676 21398
rect 9744 21342 9800 21398
rect 7884 21218 7940 21274
rect 8008 21218 8064 21274
rect 8132 21218 8188 21274
rect 8256 21218 8312 21274
rect 8380 21218 8436 21274
rect 8504 21218 8560 21274
rect 8628 21218 8684 21274
rect 8752 21218 8808 21274
rect 8876 21218 8932 21274
rect 9000 21218 9056 21274
rect 9124 21218 9180 21274
rect 9248 21218 9304 21274
rect 9372 21218 9428 21274
rect 9496 21218 9552 21274
rect 9620 21218 9676 21274
rect 9744 21218 9800 21274
rect 7884 21094 7940 21150
rect 8008 21094 8064 21150
rect 8132 21094 8188 21150
rect 8256 21094 8312 21150
rect 8380 21094 8436 21150
rect 8504 21094 8560 21150
rect 8628 21094 8684 21150
rect 8752 21094 8808 21150
rect 8876 21094 8932 21150
rect 9000 21094 9056 21150
rect 9124 21094 9180 21150
rect 9248 21094 9304 21150
rect 9372 21094 9428 21150
rect 9496 21094 9552 21150
rect 9620 21094 9676 21150
rect 9744 21094 9800 21150
rect 7884 20970 7940 21026
rect 8008 20970 8064 21026
rect 8132 20970 8188 21026
rect 8256 20970 8312 21026
rect 8380 20970 8436 21026
rect 8504 20970 8560 21026
rect 8628 20970 8684 21026
rect 8752 20970 8808 21026
rect 8876 20970 8932 21026
rect 9000 20970 9056 21026
rect 9124 20970 9180 21026
rect 9248 20970 9304 21026
rect 9372 20970 9428 21026
rect 9496 20970 9552 21026
rect 9620 20970 9676 21026
rect 9744 20970 9800 21026
rect 7884 20846 7940 20902
rect 8008 20846 8064 20902
rect 8132 20846 8188 20902
rect 8256 20846 8312 20902
rect 8380 20846 8436 20902
rect 8504 20846 8560 20902
rect 8628 20846 8684 20902
rect 8752 20846 8808 20902
rect 8876 20846 8932 20902
rect 9000 20846 9056 20902
rect 9124 20846 9180 20902
rect 9248 20846 9304 20902
rect 9372 20846 9428 20902
rect 9496 20846 9552 20902
rect 9620 20846 9676 20902
rect 9744 20846 9800 20902
rect 10254 23698 10310 23754
rect 10378 23698 10434 23754
rect 10502 23698 10558 23754
rect 10626 23698 10682 23754
rect 10750 23698 10806 23754
rect 10874 23698 10930 23754
rect 10998 23698 11054 23754
rect 11122 23698 11178 23754
rect 11246 23698 11302 23754
rect 11370 23698 11426 23754
rect 11494 23698 11550 23754
rect 11618 23698 11674 23754
rect 11742 23698 11798 23754
rect 11866 23698 11922 23754
rect 11990 23698 12046 23754
rect 12114 23698 12170 23754
rect 10254 23574 10310 23630
rect 10378 23574 10434 23630
rect 10502 23574 10558 23630
rect 10626 23574 10682 23630
rect 10750 23574 10806 23630
rect 10874 23574 10930 23630
rect 10998 23574 11054 23630
rect 11122 23574 11178 23630
rect 11246 23574 11302 23630
rect 11370 23574 11426 23630
rect 11494 23574 11550 23630
rect 11618 23574 11674 23630
rect 11742 23574 11798 23630
rect 11866 23574 11922 23630
rect 11990 23574 12046 23630
rect 12114 23574 12170 23630
rect 10254 23450 10310 23506
rect 10378 23450 10434 23506
rect 10502 23450 10558 23506
rect 10626 23450 10682 23506
rect 10750 23450 10806 23506
rect 10874 23450 10930 23506
rect 10998 23450 11054 23506
rect 11122 23450 11178 23506
rect 11246 23450 11302 23506
rect 11370 23450 11426 23506
rect 11494 23450 11550 23506
rect 11618 23450 11674 23506
rect 11742 23450 11798 23506
rect 11866 23450 11922 23506
rect 11990 23450 12046 23506
rect 12114 23450 12170 23506
rect 10254 23326 10310 23382
rect 10378 23326 10434 23382
rect 10502 23326 10558 23382
rect 10626 23326 10682 23382
rect 10750 23326 10806 23382
rect 10874 23326 10930 23382
rect 10998 23326 11054 23382
rect 11122 23326 11178 23382
rect 11246 23326 11302 23382
rect 11370 23326 11426 23382
rect 11494 23326 11550 23382
rect 11618 23326 11674 23382
rect 11742 23326 11798 23382
rect 11866 23326 11922 23382
rect 11990 23326 12046 23382
rect 12114 23326 12170 23382
rect 10254 23202 10310 23258
rect 10378 23202 10434 23258
rect 10502 23202 10558 23258
rect 10626 23202 10682 23258
rect 10750 23202 10806 23258
rect 10874 23202 10930 23258
rect 10998 23202 11054 23258
rect 11122 23202 11178 23258
rect 11246 23202 11302 23258
rect 11370 23202 11426 23258
rect 11494 23202 11550 23258
rect 11618 23202 11674 23258
rect 11742 23202 11798 23258
rect 11866 23202 11922 23258
rect 11990 23202 12046 23258
rect 12114 23202 12170 23258
rect 10254 23078 10310 23134
rect 10378 23078 10434 23134
rect 10502 23078 10558 23134
rect 10626 23078 10682 23134
rect 10750 23078 10806 23134
rect 10874 23078 10930 23134
rect 10998 23078 11054 23134
rect 11122 23078 11178 23134
rect 11246 23078 11302 23134
rect 11370 23078 11426 23134
rect 11494 23078 11550 23134
rect 11618 23078 11674 23134
rect 11742 23078 11798 23134
rect 11866 23078 11922 23134
rect 11990 23078 12046 23134
rect 12114 23078 12170 23134
rect 10254 22954 10310 23010
rect 10378 22954 10434 23010
rect 10502 22954 10558 23010
rect 10626 22954 10682 23010
rect 10750 22954 10806 23010
rect 10874 22954 10930 23010
rect 10998 22954 11054 23010
rect 11122 22954 11178 23010
rect 11246 22954 11302 23010
rect 11370 22954 11426 23010
rect 11494 22954 11550 23010
rect 11618 22954 11674 23010
rect 11742 22954 11798 23010
rect 11866 22954 11922 23010
rect 11990 22954 12046 23010
rect 12114 22954 12170 23010
rect 10254 22830 10310 22886
rect 10378 22830 10434 22886
rect 10502 22830 10558 22886
rect 10626 22830 10682 22886
rect 10750 22830 10806 22886
rect 10874 22830 10930 22886
rect 10998 22830 11054 22886
rect 11122 22830 11178 22886
rect 11246 22830 11302 22886
rect 11370 22830 11426 22886
rect 11494 22830 11550 22886
rect 11618 22830 11674 22886
rect 11742 22830 11798 22886
rect 11866 22830 11922 22886
rect 11990 22830 12046 22886
rect 12114 22830 12170 22886
rect 10254 22706 10310 22762
rect 10378 22706 10434 22762
rect 10502 22706 10558 22762
rect 10626 22706 10682 22762
rect 10750 22706 10806 22762
rect 10874 22706 10930 22762
rect 10998 22706 11054 22762
rect 11122 22706 11178 22762
rect 11246 22706 11302 22762
rect 11370 22706 11426 22762
rect 11494 22706 11550 22762
rect 11618 22706 11674 22762
rect 11742 22706 11798 22762
rect 11866 22706 11922 22762
rect 11990 22706 12046 22762
rect 12114 22706 12170 22762
rect 10254 22582 10310 22638
rect 10378 22582 10434 22638
rect 10502 22582 10558 22638
rect 10626 22582 10682 22638
rect 10750 22582 10806 22638
rect 10874 22582 10930 22638
rect 10998 22582 11054 22638
rect 11122 22582 11178 22638
rect 11246 22582 11302 22638
rect 11370 22582 11426 22638
rect 11494 22582 11550 22638
rect 11618 22582 11674 22638
rect 11742 22582 11798 22638
rect 11866 22582 11922 22638
rect 11990 22582 12046 22638
rect 12114 22582 12170 22638
rect 10254 22458 10310 22514
rect 10378 22458 10434 22514
rect 10502 22458 10558 22514
rect 10626 22458 10682 22514
rect 10750 22458 10806 22514
rect 10874 22458 10930 22514
rect 10998 22458 11054 22514
rect 11122 22458 11178 22514
rect 11246 22458 11302 22514
rect 11370 22458 11426 22514
rect 11494 22458 11550 22514
rect 11618 22458 11674 22514
rect 11742 22458 11798 22514
rect 11866 22458 11922 22514
rect 11990 22458 12046 22514
rect 12114 22458 12170 22514
rect 10254 22334 10310 22390
rect 10378 22334 10434 22390
rect 10502 22334 10558 22390
rect 10626 22334 10682 22390
rect 10750 22334 10806 22390
rect 10874 22334 10930 22390
rect 10998 22334 11054 22390
rect 11122 22334 11178 22390
rect 11246 22334 11302 22390
rect 11370 22334 11426 22390
rect 11494 22334 11550 22390
rect 11618 22334 11674 22390
rect 11742 22334 11798 22390
rect 11866 22334 11922 22390
rect 11990 22334 12046 22390
rect 12114 22334 12170 22390
rect 10254 22210 10310 22266
rect 10378 22210 10434 22266
rect 10502 22210 10558 22266
rect 10626 22210 10682 22266
rect 10750 22210 10806 22266
rect 10874 22210 10930 22266
rect 10998 22210 11054 22266
rect 11122 22210 11178 22266
rect 11246 22210 11302 22266
rect 11370 22210 11426 22266
rect 11494 22210 11550 22266
rect 11618 22210 11674 22266
rect 11742 22210 11798 22266
rect 11866 22210 11922 22266
rect 11990 22210 12046 22266
rect 12114 22210 12170 22266
rect 10254 22086 10310 22142
rect 10378 22086 10434 22142
rect 10502 22086 10558 22142
rect 10626 22086 10682 22142
rect 10750 22086 10806 22142
rect 10874 22086 10930 22142
rect 10998 22086 11054 22142
rect 11122 22086 11178 22142
rect 11246 22086 11302 22142
rect 11370 22086 11426 22142
rect 11494 22086 11550 22142
rect 11618 22086 11674 22142
rect 11742 22086 11798 22142
rect 11866 22086 11922 22142
rect 11990 22086 12046 22142
rect 12114 22086 12170 22142
rect 10254 21962 10310 22018
rect 10378 21962 10434 22018
rect 10502 21962 10558 22018
rect 10626 21962 10682 22018
rect 10750 21962 10806 22018
rect 10874 21962 10930 22018
rect 10998 21962 11054 22018
rect 11122 21962 11178 22018
rect 11246 21962 11302 22018
rect 11370 21962 11426 22018
rect 11494 21962 11550 22018
rect 11618 21962 11674 22018
rect 11742 21962 11798 22018
rect 11866 21962 11922 22018
rect 11990 21962 12046 22018
rect 12114 21962 12170 22018
rect 10254 21838 10310 21894
rect 10378 21838 10434 21894
rect 10502 21838 10558 21894
rect 10626 21838 10682 21894
rect 10750 21838 10806 21894
rect 10874 21838 10930 21894
rect 10998 21838 11054 21894
rect 11122 21838 11178 21894
rect 11246 21838 11302 21894
rect 11370 21838 11426 21894
rect 11494 21838 11550 21894
rect 11618 21838 11674 21894
rect 11742 21838 11798 21894
rect 11866 21838 11922 21894
rect 11990 21838 12046 21894
rect 12114 21838 12170 21894
rect 10254 21714 10310 21770
rect 10378 21714 10434 21770
rect 10502 21714 10558 21770
rect 10626 21714 10682 21770
rect 10750 21714 10806 21770
rect 10874 21714 10930 21770
rect 10998 21714 11054 21770
rect 11122 21714 11178 21770
rect 11246 21714 11302 21770
rect 11370 21714 11426 21770
rect 11494 21714 11550 21770
rect 11618 21714 11674 21770
rect 11742 21714 11798 21770
rect 11866 21714 11922 21770
rect 11990 21714 12046 21770
rect 12114 21714 12170 21770
rect 10254 21590 10310 21646
rect 10378 21590 10434 21646
rect 10502 21590 10558 21646
rect 10626 21590 10682 21646
rect 10750 21590 10806 21646
rect 10874 21590 10930 21646
rect 10998 21590 11054 21646
rect 11122 21590 11178 21646
rect 11246 21590 11302 21646
rect 11370 21590 11426 21646
rect 11494 21590 11550 21646
rect 11618 21590 11674 21646
rect 11742 21590 11798 21646
rect 11866 21590 11922 21646
rect 11990 21590 12046 21646
rect 12114 21590 12170 21646
rect 10254 21466 10310 21522
rect 10378 21466 10434 21522
rect 10502 21466 10558 21522
rect 10626 21466 10682 21522
rect 10750 21466 10806 21522
rect 10874 21466 10930 21522
rect 10998 21466 11054 21522
rect 11122 21466 11178 21522
rect 11246 21466 11302 21522
rect 11370 21466 11426 21522
rect 11494 21466 11550 21522
rect 11618 21466 11674 21522
rect 11742 21466 11798 21522
rect 11866 21466 11922 21522
rect 11990 21466 12046 21522
rect 12114 21466 12170 21522
rect 10254 21342 10310 21398
rect 10378 21342 10434 21398
rect 10502 21342 10558 21398
rect 10626 21342 10682 21398
rect 10750 21342 10806 21398
rect 10874 21342 10930 21398
rect 10998 21342 11054 21398
rect 11122 21342 11178 21398
rect 11246 21342 11302 21398
rect 11370 21342 11426 21398
rect 11494 21342 11550 21398
rect 11618 21342 11674 21398
rect 11742 21342 11798 21398
rect 11866 21342 11922 21398
rect 11990 21342 12046 21398
rect 12114 21342 12170 21398
rect 10254 21218 10310 21274
rect 10378 21218 10434 21274
rect 10502 21218 10558 21274
rect 10626 21218 10682 21274
rect 10750 21218 10806 21274
rect 10874 21218 10930 21274
rect 10998 21218 11054 21274
rect 11122 21218 11178 21274
rect 11246 21218 11302 21274
rect 11370 21218 11426 21274
rect 11494 21218 11550 21274
rect 11618 21218 11674 21274
rect 11742 21218 11798 21274
rect 11866 21218 11922 21274
rect 11990 21218 12046 21274
rect 12114 21218 12170 21274
rect 10254 21094 10310 21150
rect 10378 21094 10434 21150
rect 10502 21094 10558 21150
rect 10626 21094 10682 21150
rect 10750 21094 10806 21150
rect 10874 21094 10930 21150
rect 10998 21094 11054 21150
rect 11122 21094 11178 21150
rect 11246 21094 11302 21150
rect 11370 21094 11426 21150
rect 11494 21094 11550 21150
rect 11618 21094 11674 21150
rect 11742 21094 11798 21150
rect 11866 21094 11922 21150
rect 11990 21094 12046 21150
rect 12114 21094 12170 21150
rect 10254 20970 10310 21026
rect 10378 20970 10434 21026
rect 10502 20970 10558 21026
rect 10626 20970 10682 21026
rect 10750 20970 10806 21026
rect 10874 20970 10930 21026
rect 10998 20970 11054 21026
rect 11122 20970 11178 21026
rect 11246 20970 11302 21026
rect 11370 20970 11426 21026
rect 11494 20970 11550 21026
rect 11618 20970 11674 21026
rect 11742 20970 11798 21026
rect 11866 20970 11922 21026
rect 11990 20970 12046 21026
rect 12114 20970 12170 21026
rect 10254 20846 10310 20902
rect 10378 20846 10434 20902
rect 10502 20846 10558 20902
rect 10626 20846 10682 20902
rect 10750 20846 10806 20902
rect 10874 20846 10930 20902
rect 10998 20846 11054 20902
rect 11122 20846 11178 20902
rect 11246 20846 11302 20902
rect 11370 20846 11426 20902
rect 11494 20846 11550 20902
rect 11618 20846 11674 20902
rect 11742 20846 11798 20902
rect 11866 20846 11922 20902
rect 11990 20846 12046 20902
rect 12114 20846 12170 20902
rect 12871 23698 12927 23754
rect 12995 23698 13051 23754
rect 13119 23698 13175 23754
rect 13243 23698 13299 23754
rect 13367 23698 13423 23754
rect 13491 23698 13547 23754
rect 13615 23698 13671 23754
rect 13739 23698 13795 23754
rect 13863 23698 13919 23754
rect 13987 23698 14043 23754
rect 14111 23698 14167 23754
rect 14235 23698 14291 23754
rect 14359 23698 14415 23754
rect 14483 23698 14539 23754
rect 14607 23698 14663 23754
rect 12871 23574 12927 23630
rect 12995 23574 13051 23630
rect 13119 23574 13175 23630
rect 13243 23574 13299 23630
rect 13367 23574 13423 23630
rect 13491 23574 13547 23630
rect 13615 23574 13671 23630
rect 13739 23574 13795 23630
rect 13863 23574 13919 23630
rect 13987 23574 14043 23630
rect 14111 23574 14167 23630
rect 14235 23574 14291 23630
rect 14359 23574 14415 23630
rect 14483 23574 14539 23630
rect 14607 23574 14663 23630
rect 12871 23450 12927 23506
rect 12995 23450 13051 23506
rect 13119 23450 13175 23506
rect 13243 23450 13299 23506
rect 13367 23450 13423 23506
rect 13491 23450 13547 23506
rect 13615 23450 13671 23506
rect 13739 23450 13795 23506
rect 13863 23450 13919 23506
rect 13987 23450 14043 23506
rect 14111 23450 14167 23506
rect 14235 23450 14291 23506
rect 14359 23450 14415 23506
rect 14483 23450 14539 23506
rect 14607 23450 14663 23506
rect 12871 23326 12927 23382
rect 12995 23326 13051 23382
rect 13119 23326 13175 23382
rect 13243 23326 13299 23382
rect 13367 23326 13423 23382
rect 13491 23326 13547 23382
rect 13615 23326 13671 23382
rect 13739 23326 13795 23382
rect 13863 23326 13919 23382
rect 13987 23326 14043 23382
rect 14111 23326 14167 23382
rect 14235 23326 14291 23382
rect 14359 23326 14415 23382
rect 14483 23326 14539 23382
rect 14607 23326 14663 23382
rect 12871 23202 12927 23258
rect 12995 23202 13051 23258
rect 13119 23202 13175 23258
rect 13243 23202 13299 23258
rect 13367 23202 13423 23258
rect 13491 23202 13547 23258
rect 13615 23202 13671 23258
rect 13739 23202 13795 23258
rect 13863 23202 13919 23258
rect 13987 23202 14043 23258
rect 14111 23202 14167 23258
rect 14235 23202 14291 23258
rect 14359 23202 14415 23258
rect 14483 23202 14539 23258
rect 14607 23202 14663 23258
rect 12871 23078 12927 23134
rect 12995 23078 13051 23134
rect 13119 23078 13175 23134
rect 13243 23078 13299 23134
rect 13367 23078 13423 23134
rect 13491 23078 13547 23134
rect 13615 23078 13671 23134
rect 13739 23078 13795 23134
rect 13863 23078 13919 23134
rect 13987 23078 14043 23134
rect 14111 23078 14167 23134
rect 14235 23078 14291 23134
rect 14359 23078 14415 23134
rect 14483 23078 14539 23134
rect 14607 23078 14663 23134
rect 12871 22954 12927 23010
rect 12995 22954 13051 23010
rect 13119 22954 13175 23010
rect 13243 22954 13299 23010
rect 13367 22954 13423 23010
rect 13491 22954 13547 23010
rect 13615 22954 13671 23010
rect 13739 22954 13795 23010
rect 13863 22954 13919 23010
rect 13987 22954 14043 23010
rect 14111 22954 14167 23010
rect 14235 22954 14291 23010
rect 14359 22954 14415 23010
rect 14483 22954 14539 23010
rect 14607 22954 14663 23010
rect 12871 22830 12927 22886
rect 12995 22830 13051 22886
rect 13119 22830 13175 22886
rect 13243 22830 13299 22886
rect 13367 22830 13423 22886
rect 13491 22830 13547 22886
rect 13615 22830 13671 22886
rect 13739 22830 13795 22886
rect 13863 22830 13919 22886
rect 13987 22830 14043 22886
rect 14111 22830 14167 22886
rect 14235 22830 14291 22886
rect 14359 22830 14415 22886
rect 14483 22830 14539 22886
rect 14607 22830 14663 22886
rect 12871 22706 12927 22762
rect 12995 22706 13051 22762
rect 13119 22706 13175 22762
rect 13243 22706 13299 22762
rect 13367 22706 13423 22762
rect 13491 22706 13547 22762
rect 13615 22706 13671 22762
rect 13739 22706 13795 22762
rect 13863 22706 13919 22762
rect 13987 22706 14043 22762
rect 14111 22706 14167 22762
rect 14235 22706 14291 22762
rect 14359 22706 14415 22762
rect 14483 22706 14539 22762
rect 14607 22706 14663 22762
rect 12871 22582 12927 22638
rect 12995 22582 13051 22638
rect 13119 22582 13175 22638
rect 13243 22582 13299 22638
rect 13367 22582 13423 22638
rect 13491 22582 13547 22638
rect 13615 22582 13671 22638
rect 13739 22582 13795 22638
rect 13863 22582 13919 22638
rect 13987 22582 14043 22638
rect 14111 22582 14167 22638
rect 14235 22582 14291 22638
rect 14359 22582 14415 22638
rect 14483 22582 14539 22638
rect 14607 22582 14663 22638
rect 12871 22458 12927 22514
rect 12995 22458 13051 22514
rect 13119 22458 13175 22514
rect 13243 22458 13299 22514
rect 13367 22458 13423 22514
rect 13491 22458 13547 22514
rect 13615 22458 13671 22514
rect 13739 22458 13795 22514
rect 13863 22458 13919 22514
rect 13987 22458 14043 22514
rect 14111 22458 14167 22514
rect 14235 22458 14291 22514
rect 14359 22458 14415 22514
rect 14483 22458 14539 22514
rect 14607 22458 14663 22514
rect 12871 22334 12927 22390
rect 12995 22334 13051 22390
rect 13119 22334 13175 22390
rect 13243 22334 13299 22390
rect 13367 22334 13423 22390
rect 13491 22334 13547 22390
rect 13615 22334 13671 22390
rect 13739 22334 13795 22390
rect 13863 22334 13919 22390
rect 13987 22334 14043 22390
rect 14111 22334 14167 22390
rect 14235 22334 14291 22390
rect 14359 22334 14415 22390
rect 14483 22334 14539 22390
rect 14607 22334 14663 22390
rect 12871 22210 12927 22266
rect 12995 22210 13051 22266
rect 13119 22210 13175 22266
rect 13243 22210 13299 22266
rect 13367 22210 13423 22266
rect 13491 22210 13547 22266
rect 13615 22210 13671 22266
rect 13739 22210 13795 22266
rect 13863 22210 13919 22266
rect 13987 22210 14043 22266
rect 14111 22210 14167 22266
rect 14235 22210 14291 22266
rect 14359 22210 14415 22266
rect 14483 22210 14539 22266
rect 14607 22210 14663 22266
rect 12871 22086 12927 22142
rect 12995 22086 13051 22142
rect 13119 22086 13175 22142
rect 13243 22086 13299 22142
rect 13367 22086 13423 22142
rect 13491 22086 13547 22142
rect 13615 22086 13671 22142
rect 13739 22086 13795 22142
rect 13863 22086 13919 22142
rect 13987 22086 14043 22142
rect 14111 22086 14167 22142
rect 14235 22086 14291 22142
rect 14359 22086 14415 22142
rect 14483 22086 14539 22142
rect 14607 22086 14663 22142
rect 12871 21962 12927 22018
rect 12995 21962 13051 22018
rect 13119 21962 13175 22018
rect 13243 21962 13299 22018
rect 13367 21962 13423 22018
rect 13491 21962 13547 22018
rect 13615 21962 13671 22018
rect 13739 21962 13795 22018
rect 13863 21962 13919 22018
rect 13987 21962 14043 22018
rect 14111 21962 14167 22018
rect 14235 21962 14291 22018
rect 14359 21962 14415 22018
rect 14483 21962 14539 22018
rect 14607 21962 14663 22018
rect 12871 21838 12927 21894
rect 12995 21838 13051 21894
rect 13119 21838 13175 21894
rect 13243 21838 13299 21894
rect 13367 21838 13423 21894
rect 13491 21838 13547 21894
rect 13615 21838 13671 21894
rect 13739 21838 13795 21894
rect 13863 21838 13919 21894
rect 13987 21838 14043 21894
rect 14111 21838 14167 21894
rect 14235 21838 14291 21894
rect 14359 21838 14415 21894
rect 14483 21838 14539 21894
rect 14607 21838 14663 21894
rect 12871 21714 12927 21770
rect 12995 21714 13051 21770
rect 13119 21714 13175 21770
rect 13243 21714 13299 21770
rect 13367 21714 13423 21770
rect 13491 21714 13547 21770
rect 13615 21714 13671 21770
rect 13739 21714 13795 21770
rect 13863 21714 13919 21770
rect 13987 21714 14043 21770
rect 14111 21714 14167 21770
rect 14235 21714 14291 21770
rect 14359 21714 14415 21770
rect 14483 21714 14539 21770
rect 14607 21714 14663 21770
rect 12871 21590 12927 21646
rect 12995 21590 13051 21646
rect 13119 21590 13175 21646
rect 13243 21590 13299 21646
rect 13367 21590 13423 21646
rect 13491 21590 13547 21646
rect 13615 21590 13671 21646
rect 13739 21590 13795 21646
rect 13863 21590 13919 21646
rect 13987 21590 14043 21646
rect 14111 21590 14167 21646
rect 14235 21590 14291 21646
rect 14359 21590 14415 21646
rect 14483 21590 14539 21646
rect 14607 21590 14663 21646
rect 12871 21466 12927 21522
rect 12995 21466 13051 21522
rect 13119 21466 13175 21522
rect 13243 21466 13299 21522
rect 13367 21466 13423 21522
rect 13491 21466 13547 21522
rect 13615 21466 13671 21522
rect 13739 21466 13795 21522
rect 13863 21466 13919 21522
rect 13987 21466 14043 21522
rect 14111 21466 14167 21522
rect 14235 21466 14291 21522
rect 14359 21466 14415 21522
rect 14483 21466 14539 21522
rect 14607 21466 14663 21522
rect 12871 21342 12927 21398
rect 12995 21342 13051 21398
rect 13119 21342 13175 21398
rect 13243 21342 13299 21398
rect 13367 21342 13423 21398
rect 13491 21342 13547 21398
rect 13615 21342 13671 21398
rect 13739 21342 13795 21398
rect 13863 21342 13919 21398
rect 13987 21342 14043 21398
rect 14111 21342 14167 21398
rect 14235 21342 14291 21398
rect 14359 21342 14415 21398
rect 14483 21342 14539 21398
rect 14607 21342 14663 21398
rect 12871 21218 12927 21274
rect 12995 21218 13051 21274
rect 13119 21218 13175 21274
rect 13243 21218 13299 21274
rect 13367 21218 13423 21274
rect 13491 21218 13547 21274
rect 13615 21218 13671 21274
rect 13739 21218 13795 21274
rect 13863 21218 13919 21274
rect 13987 21218 14043 21274
rect 14111 21218 14167 21274
rect 14235 21218 14291 21274
rect 14359 21218 14415 21274
rect 14483 21218 14539 21274
rect 14607 21218 14663 21274
rect 12871 21094 12927 21150
rect 12995 21094 13051 21150
rect 13119 21094 13175 21150
rect 13243 21094 13299 21150
rect 13367 21094 13423 21150
rect 13491 21094 13547 21150
rect 13615 21094 13671 21150
rect 13739 21094 13795 21150
rect 13863 21094 13919 21150
rect 13987 21094 14043 21150
rect 14111 21094 14167 21150
rect 14235 21094 14291 21150
rect 14359 21094 14415 21150
rect 14483 21094 14539 21150
rect 14607 21094 14663 21150
rect 12871 20970 12927 21026
rect 12995 20970 13051 21026
rect 13119 20970 13175 21026
rect 13243 20970 13299 21026
rect 13367 20970 13423 21026
rect 13491 20970 13547 21026
rect 13615 20970 13671 21026
rect 13739 20970 13795 21026
rect 13863 20970 13919 21026
rect 13987 20970 14043 21026
rect 14111 20970 14167 21026
rect 14235 20970 14291 21026
rect 14359 20970 14415 21026
rect 14483 20970 14539 21026
rect 14607 20970 14663 21026
rect 12871 20846 12927 20902
rect 12995 20846 13051 20902
rect 13119 20846 13175 20902
rect 13243 20846 13299 20902
rect 13367 20846 13423 20902
rect 13491 20846 13547 20902
rect 13615 20846 13671 20902
rect 13739 20846 13795 20902
rect 13863 20846 13919 20902
rect 13987 20846 14043 20902
rect 14111 20846 14167 20902
rect 14235 20846 14291 20902
rect 14359 20846 14415 20902
rect 14483 20846 14539 20902
rect 14607 20846 14663 20902
rect 315 20498 371 20554
rect 439 20498 495 20554
rect 563 20498 619 20554
rect 687 20498 743 20554
rect 811 20498 867 20554
rect 935 20498 991 20554
rect 1059 20498 1115 20554
rect 1183 20498 1239 20554
rect 1307 20498 1363 20554
rect 1431 20498 1487 20554
rect 1555 20498 1611 20554
rect 1679 20498 1735 20554
rect 1803 20498 1859 20554
rect 1927 20498 1983 20554
rect 2051 20498 2107 20554
rect 315 20374 371 20430
rect 439 20374 495 20430
rect 563 20374 619 20430
rect 687 20374 743 20430
rect 811 20374 867 20430
rect 935 20374 991 20430
rect 1059 20374 1115 20430
rect 1183 20374 1239 20430
rect 1307 20374 1363 20430
rect 1431 20374 1487 20430
rect 1555 20374 1611 20430
rect 1679 20374 1735 20430
rect 1803 20374 1859 20430
rect 1927 20374 1983 20430
rect 2051 20374 2107 20430
rect 315 20250 371 20306
rect 439 20250 495 20306
rect 563 20250 619 20306
rect 687 20250 743 20306
rect 811 20250 867 20306
rect 935 20250 991 20306
rect 1059 20250 1115 20306
rect 1183 20250 1239 20306
rect 1307 20250 1363 20306
rect 1431 20250 1487 20306
rect 1555 20250 1611 20306
rect 1679 20250 1735 20306
rect 1803 20250 1859 20306
rect 1927 20250 1983 20306
rect 2051 20250 2107 20306
rect 315 20126 371 20182
rect 439 20126 495 20182
rect 563 20126 619 20182
rect 687 20126 743 20182
rect 811 20126 867 20182
rect 935 20126 991 20182
rect 1059 20126 1115 20182
rect 1183 20126 1239 20182
rect 1307 20126 1363 20182
rect 1431 20126 1487 20182
rect 1555 20126 1611 20182
rect 1679 20126 1735 20182
rect 1803 20126 1859 20182
rect 1927 20126 1983 20182
rect 2051 20126 2107 20182
rect 315 20002 371 20058
rect 439 20002 495 20058
rect 563 20002 619 20058
rect 687 20002 743 20058
rect 811 20002 867 20058
rect 935 20002 991 20058
rect 1059 20002 1115 20058
rect 1183 20002 1239 20058
rect 1307 20002 1363 20058
rect 1431 20002 1487 20058
rect 1555 20002 1611 20058
rect 1679 20002 1735 20058
rect 1803 20002 1859 20058
rect 1927 20002 1983 20058
rect 2051 20002 2107 20058
rect 315 19878 371 19934
rect 439 19878 495 19934
rect 563 19878 619 19934
rect 687 19878 743 19934
rect 811 19878 867 19934
rect 935 19878 991 19934
rect 1059 19878 1115 19934
rect 1183 19878 1239 19934
rect 1307 19878 1363 19934
rect 1431 19878 1487 19934
rect 1555 19878 1611 19934
rect 1679 19878 1735 19934
rect 1803 19878 1859 19934
rect 1927 19878 1983 19934
rect 2051 19878 2107 19934
rect 315 19754 371 19810
rect 439 19754 495 19810
rect 563 19754 619 19810
rect 687 19754 743 19810
rect 811 19754 867 19810
rect 935 19754 991 19810
rect 1059 19754 1115 19810
rect 1183 19754 1239 19810
rect 1307 19754 1363 19810
rect 1431 19754 1487 19810
rect 1555 19754 1611 19810
rect 1679 19754 1735 19810
rect 1803 19754 1859 19810
rect 1927 19754 1983 19810
rect 2051 19754 2107 19810
rect 315 19630 371 19686
rect 439 19630 495 19686
rect 563 19630 619 19686
rect 687 19630 743 19686
rect 811 19630 867 19686
rect 935 19630 991 19686
rect 1059 19630 1115 19686
rect 1183 19630 1239 19686
rect 1307 19630 1363 19686
rect 1431 19630 1487 19686
rect 1555 19630 1611 19686
rect 1679 19630 1735 19686
rect 1803 19630 1859 19686
rect 1927 19630 1983 19686
rect 2051 19630 2107 19686
rect 315 19506 371 19562
rect 439 19506 495 19562
rect 563 19506 619 19562
rect 687 19506 743 19562
rect 811 19506 867 19562
rect 935 19506 991 19562
rect 1059 19506 1115 19562
rect 1183 19506 1239 19562
rect 1307 19506 1363 19562
rect 1431 19506 1487 19562
rect 1555 19506 1611 19562
rect 1679 19506 1735 19562
rect 1803 19506 1859 19562
rect 1927 19506 1983 19562
rect 2051 19506 2107 19562
rect 315 19382 371 19438
rect 439 19382 495 19438
rect 563 19382 619 19438
rect 687 19382 743 19438
rect 811 19382 867 19438
rect 935 19382 991 19438
rect 1059 19382 1115 19438
rect 1183 19382 1239 19438
rect 1307 19382 1363 19438
rect 1431 19382 1487 19438
rect 1555 19382 1611 19438
rect 1679 19382 1735 19438
rect 1803 19382 1859 19438
rect 1927 19382 1983 19438
rect 2051 19382 2107 19438
rect 315 19258 371 19314
rect 439 19258 495 19314
rect 563 19258 619 19314
rect 687 19258 743 19314
rect 811 19258 867 19314
rect 935 19258 991 19314
rect 1059 19258 1115 19314
rect 1183 19258 1239 19314
rect 1307 19258 1363 19314
rect 1431 19258 1487 19314
rect 1555 19258 1611 19314
rect 1679 19258 1735 19314
rect 1803 19258 1859 19314
rect 1927 19258 1983 19314
rect 2051 19258 2107 19314
rect 315 19134 371 19190
rect 439 19134 495 19190
rect 563 19134 619 19190
rect 687 19134 743 19190
rect 811 19134 867 19190
rect 935 19134 991 19190
rect 1059 19134 1115 19190
rect 1183 19134 1239 19190
rect 1307 19134 1363 19190
rect 1431 19134 1487 19190
rect 1555 19134 1611 19190
rect 1679 19134 1735 19190
rect 1803 19134 1859 19190
rect 1927 19134 1983 19190
rect 2051 19134 2107 19190
rect 315 19010 371 19066
rect 439 19010 495 19066
rect 563 19010 619 19066
rect 687 19010 743 19066
rect 811 19010 867 19066
rect 935 19010 991 19066
rect 1059 19010 1115 19066
rect 1183 19010 1239 19066
rect 1307 19010 1363 19066
rect 1431 19010 1487 19066
rect 1555 19010 1611 19066
rect 1679 19010 1735 19066
rect 1803 19010 1859 19066
rect 1927 19010 1983 19066
rect 2051 19010 2107 19066
rect 315 18886 371 18942
rect 439 18886 495 18942
rect 563 18886 619 18942
rect 687 18886 743 18942
rect 811 18886 867 18942
rect 935 18886 991 18942
rect 1059 18886 1115 18942
rect 1183 18886 1239 18942
rect 1307 18886 1363 18942
rect 1431 18886 1487 18942
rect 1555 18886 1611 18942
rect 1679 18886 1735 18942
rect 1803 18886 1859 18942
rect 1927 18886 1983 18942
rect 2051 18886 2107 18942
rect 315 18762 371 18818
rect 439 18762 495 18818
rect 563 18762 619 18818
rect 687 18762 743 18818
rect 811 18762 867 18818
rect 935 18762 991 18818
rect 1059 18762 1115 18818
rect 1183 18762 1239 18818
rect 1307 18762 1363 18818
rect 1431 18762 1487 18818
rect 1555 18762 1611 18818
rect 1679 18762 1735 18818
rect 1803 18762 1859 18818
rect 1927 18762 1983 18818
rect 2051 18762 2107 18818
rect 315 18638 371 18694
rect 439 18638 495 18694
rect 563 18638 619 18694
rect 687 18638 743 18694
rect 811 18638 867 18694
rect 935 18638 991 18694
rect 1059 18638 1115 18694
rect 1183 18638 1239 18694
rect 1307 18638 1363 18694
rect 1431 18638 1487 18694
rect 1555 18638 1611 18694
rect 1679 18638 1735 18694
rect 1803 18638 1859 18694
rect 1927 18638 1983 18694
rect 2051 18638 2107 18694
rect 315 18514 371 18570
rect 439 18514 495 18570
rect 563 18514 619 18570
rect 687 18514 743 18570
rect 811 18514 867 18570
rect 935 18514 991 18570
rect 1059 18514 1115 18570
rect 1183 18514 1239 18570
rect 1307 18514 1363 18570
rect 1431 18514 1487 18570
rect 1555 18514 1611 18570
rect 1679 18514 1735 18570
rect 1803 18514 1859 18570
rect 1927 18514 1983 18570
rect 2051 18514 2107 18570
rect 315 18390 371 18446
rect 439 18390 495 18446
rect 563 18390 619 18446
rect 687 18390 743 18446
rect 811 18390 867 18446
rect 935 18390 991 18446
rect 1059 18390 1115 18446
rect 1183 18390 1239 18446
rect 1307 18390 1363 18446
rect 1431 18390 1487 18446
rect 1555 18390 1611 18446
rect 1679 18390 1735 18446
rect 1803 18390 1859 18446
rect 1927 18390 1983 18446
rect 2051 18390 2107 18446
rect 315 18266 371 18322
rect 439 18266 495 18322
rect 563 18266 619 18322
rect 687 18266 743 18322
rect 811 18266 867 18322
rect 935 18266 991 18322
rect 1059 18266 1115 18322
rect 1183 18266 1239 18322
rect 1307 18266 1363 18322
rect 1431 18266 1487 18322
rect 1555 18266 1611 18322
rect 1679 18266 1735 18322
rect 1803 18266 1859 18322
rect 1927 18266 1983 18322
rect 2051 18266 2107 18322
rect 315 18142 371 18198
rect 439 18142 495 18198
rect 563 18142 619 18198
rect 687 18142 743 18198
rect 811 18142 867 18198
rect 935 18142 991 18198
rect 1059 18142 1115 18198
rect 1183 18142 1239 18198
rect 1307 18142 1363 18198
rect 1431 18142 1487 18198
rect 1555 18142 1611 18198
rect 1679 18142 1735 18198
rect 1803 18142 1859 18198
rect 1927 18142 1983 18198
rect 2051 18142 2107 18198
rect 315 18018 371 18074
rect 439 18018 495 18074
rect 563 18018 619 18074
rect 687 18018 743 18074
rect 811 18018 867 18074
rect 935 18018 991 18074
rect 1059 18018 1115 18074
rect 1183 18018 1239 18074
rect 1307 18018 1363 18074
rect 1431 18018 1487 18074
rect 1555 18018 1611 18074
rect 1679 18018 1735 18074
rect 1803 18018 1859 18074
rect 1927 18018 1983 18074
rect 2051 18018 2107 18074
rect 315 17894 371 17950
rect 439 17894 495 17950
rect 563 17894 619 17950
rect 687 17894 743 17950
rect 811 17894 867 17950
rect 935 17894 991 17950
rect 1059 17894 1115 17950
rect 1183 17894 1239 17950
rect 1307 17894 1363 17950
rect 1431 17894 1487 17950
rect 1555 17894 1611 17950
rect 1679 17894 1735 17950
rect 1803 17894 1859 17950
rect 1927 17894 1983 17950
rect 2051 17894 2107 17950
rect 315 17770 371 17826
rect 439 17770 495 17826
rect 563 17770 619 17826
rect 687 17770 743 17826
rect 811 17770 867 17826
rect 935 17770 991 17826
rect 1059 17770 1115 17826
rect 1183 17770 1239 17826
rect 1307 17770 1363 17826
rect 1431 17770 1487 17826
rect 1555 17770 1611 17826
rect 1679 17770 1735 17826
rect 1803 17770 1859 17826
rect 1927 17770 1983 17826
rect 2051 17770 2107 17826
rect 315 17646 371 17702
rect 439 17646 495 17702
rect 563 17646 619 17702
rect 687 17646 743 17702
rect 811 17646 867 17702
rect 935 17646 991 17702
rect 1059 17646 1115 17702
rect 1183 17646 1239 17702
rect 1307 17646 1363 17702
rect 1431 17646 1487 17702
rect 1555 17646 1611 17702
rect 1679 17646 1735 17702
rect 1803 17646 1859 17702
rect 1927 17646 1983 17702
rect 2051 17646 2107 17702
rect 2808 20498 2864 20554
rect 2932 20498 2988 20554
rect 3056 20498 3112 20554
rect 3180 20498 3236 20554
rect 3304 20498 3360 20554
rect 3428 20498 3484 20554
rect 3552 20498 3608 20554
rect 3676 20498 3732 20554
rect 3800 20498 3856 20554
rect 3924 20498 3980 20554
rect 4048 20498 4104 20554
rect 4172 20498 4228 20554
rect 4296 20498 4352 20554
rect 4420 20498 4476 20554
rect 4544 20498 4600 20554
rect 4668 20498 4724 20554
rect 2808 20374 2864 20430
rect 2932 20374 2988 20430
rect 3056 20374 3112 20430
rect 3180 20374 3236 20430
rect 3304 20374 3360 20430
rect 3428 20374 3484 20430
rect 3552 20374 3608 20430
rect 3676 20374 3732 20430
rect 3800 20374 3856 20430
rect 3924 20374 3980 20430
rect 4048 20374 4104 20430
rect 4172 20374 4228 20430
rect 4296 20374 4352 20430
rect 4420 20374 4476 20430
rect 4544 20374 4600 20430
rect 4668 20374 4724 20430
rect 2808 20250 2864 20306
rect 2932 20250 2988 20306
rect 3056 20250 3112 20306
rect 3180 20250 3236 20306
rect 3304 20250 3360 20306
rect 3428 20250 3484 20306
rect 3552 20250 3608 20306
rect 3676 20250 3732 20306
rect 3800 20250 3856 20306
rect 3924 20250 3980 20306
rect 4048 20250 4104 20306
rect 4172 20250 4228 20306
rect 4296 20250 4352 20306
rect 4420 20250 4476 20306
rect 4544 20250 4600 20306
rect 4668 20250 4724 20306
rect 2808 20126 2864 20182
rect 2932 20126 2988 20182
rect 3056 20126 3112 20182
rect 3180 20126 3236 20182
rect 3304 20126 3360 20182
rect 3428 20126 3484 20182
rect 3552 20126 3608 20182
rect 3676 20126 3732 20182
rect 3800 20126 3856 20182
rect 3924 20126 3980 20182
rect 4048 20126 4104 20182
rect 4172 20126 4228 20182
rect 4296 20126 4352 20182
rect 4420 20126 4476 20182
rect 4544 20126 4600 20182
rect 4668 20126 4724 20182
rect 2808 20002 2864 20058
rect 2932 20002 2988 20058
rect 3056 20002 3112 20058
rect 3180 20002 3236 20058
rect 3304 20002 3360 20058
rect 3428 20002 3484 20058
rect 3552 20002 3608 20058
rect 3676 20002 3732 20058
rect 3800 20002 3856 20058
rect 3924 20002 3980 20058
rect 4048 20002 4104 20058
rect 4172 20002 4228 20058
rect 4296 20002 4352 20058
rect 4420 20002 4476 20058
rect 4544 20002 4600 20058
rect 4668 20002 4724 20058
rect 2808 19878 2864 19934
rect 2932 19878 2988 19934
rect 3056 19878 3112 19934
rect 3180 19878 3236 19934
rect 3304 19878 3360 19934
rect 3428 19878 3484 19934
rect 3552 19878 3608 19934
rect 3676 19878 3732 19934
rect 3800 19878 3856 19934
rect 3924 19878 3980 19934
rect 4048 19878 4104 19934
rect 4172 19878 4228 19934
rect 4296 19878 4352 19934
rect 4420 19878 4476 19934
rect 4544 19878 4600 19934
rect 4668 19878 4724 19934
rect 2808 19754 2864 19810
rect 2932 19754 2988 19810
rect 3056 19754 3112 19810
rect 3180 19754 3236 19810
rect 3304 19754 3360 19810
rect 3428 19754 3484 19810
rect 3552 19754 3608 19810
rect 3676 19754 3732 19810
rect 3800 19754 3856 19810
rect 3924 19754 3980 19810
rect 4048 19754 4104 19810
rect 4172 19754 4228 19810
rect 4296 19754 4352 19810
rect 4420 19754 4476 19810
rect 4544 19754 4600 19810
rect 4668 19754 4724 19810
rect 2808 19630 2864 19686
rect 2932 19630 2988 19686
rect 3056 19630 3112 19686
rect 3180 19630 3236 19686
rect 3304 19630 3360 19686
rect 3428 19630 3484 19686
rect 3552 19630 3608 19686
rect 3676 19630 3732 19686
rect 3800 19630 3856 19686
rect 3924 19630 3980 19686
rect 4048 19630 4104 19686
rect 4172 19630 4228 19686
rect 4296 19630 4352 19686
rect 4420 19630 4476 19686
rect 4544 19630 4600 19686
rect 4668 19630 4724 19686
rect 2808 19506 2864 19562
rect 2932 19506 2988 19562
rect 3056 19506 3112 19562
rect 3180 19506 3236 19562
rect 3304 19506 3360 19562
rect 3428 19506 3484 19562
rect 3552 19506 3608 19562
rect 3676 19506 3732 19562
rect 3800 19506 3856 19562
rect 3924 19506 3980 19562
rect 4048 19506 4104 19562
rect 4172 19506 4228 19562
rect 4296 19506 4352 19562
rect 4420 19506 4476 19562
rect 4544 19506 4600 19562
rect 4668 19506 4724 19562
rect 2808 19382 2864 19438
rect 2932 19382 2988 19438
rect 3056 19382 3112 19438
rect 3180 19382 3236 19438
rect 3304 19382 3360 19438
rect 3428 19382 3484 19438
rect 3552 19382 3608 19438
rect 3676 19382 3732 19438
rect 3800 19382 3856 19438
rect 3924 19382 3980 19438
rect 4048 19382 4104 19438
rect 4172 19382 4228 19438
rect 4296 19382 4352 19438
rect 4420 19382 4476 19438
rect 4544 19382 4600 19438
rect 4668 19382 4724 19438
rect 2808 19258 2864 19314
rect 2932 19258 2988 19314
rect 3056 19258 3112 19314
rect 3180 19258 3236 19314
rect 3304 19258 3360 19314
rect 3428 19258 3484 19314
rect 3552 19258 3608 19314
rect 3676 19258 3732 19314
rect 3800 19258 3856 19314
rect 3924 19258 3980 19314
rect 4048 19258 4104 19314
rect 4172 19258 4228 19314
rect 4296 19258 4352 19314
rect 4420 19258 4476 19314
rect 4544 19258 4600 19314
rect 4668 19258 4724 19314
rect 2808 19134 2864 19190
rect 2932 19134 2988 19190
rect 3056 19134 3112 19190
rect 3180 19134 3236 19190
rect 3304 19134 3360 19190
rect 3428 19134 3484 19190
rect 3552 19134 3608 19190
rect 3676 19134 3732 19190
rect 3800 19134 3856 19190
rect 3924 19134 3980 19190
rect 4048 19134 4104 19190
rect 4172 19134 4228 19190
rect 4296 19134 4352 19190
rect 4420 19134 4476 19190
rect 4544 19134 4600 19190
rect 4668 19134 4724 19190
rect 2808 19010 2864 19066
rect 2932 19010 2988 19066
rect 3056 19010 3112 19066
rect 3180 19010 3236 19066
rect 3304 19010 3360 19066
rect 3428 19010 3484 19066
rect 3552 19010 3608 19066
rect 3676 19010 3732 19066
rect 3800 19010 3856 19066
rect 3924 19010 3980 19066
rect 4048 19010 4104 19066
rect 4172 19010 4228 19066
rect 4296 19010 4352 19066
rect 4420 19010 4476 19066
rect 4544 19010 4600 19066
rect 4668 19010 4724 19066
rect 2808 18886 2864 18942
rect 2932 18886 2988 18942
rect 3056 18886 3112 18942
rect 3180 18886 3236 18942
rect 3304 18886 3360 18942
rect 3428 18886 3484 18942
rect 3552 18886 3608 18942
rect 3676 18886 3732 18942
rect 3800 18886 3856 18942
rect 3924 18886 3980 18942
rect 4048 18886 4104 18942
rect 4172 18886 4228 18942
rect 4296 18886 4352 18942
rect 4420 18886 4476 18942
rect 4544 18886 4600 18942
rect 4668 18886 4724 18942
rect 2808 18762 2864 18818
rect 2932 18762 2988 18818
rect 3056 18762 3112 18818
rect 3180 18762 3236 18818
rect 3304 18762 3360 18818
rect 3428 18762 3484 18818
rect 3552 18762 3608 18818
rect 3676 18762 3732 18818
rect 3800 18762 3856 18818
rect 3924 18762 3980 18818
rect 4048 18762 4104 18818
rect 4172 18762 4228 18818
rect 4296 18762 4352 18818
rect 4420 18762 4476 18818
rect 4544 18762 4600 18818
rect 4668 18762 4724 18818
rect 2808 18638 2864 18694
rect 2932 18638 2988 18694
rect 3056 18638 3112 18694
rect 3180 18638 3236 18694
rect 3304 18638 3360 18694
rect 3428 18638 3484 18694
rect 3552 18638 3608 18694
rect 3676 18638 3732 18694
rect 3800 18638 3856 18694
rect 3924 18638 3980 18694
rect 4048 18638 4104 18694
rect 4172 18638 4228 18694
rect 4296 18638 4352 18694
rect 4420 18638 4476 18694
rect 4544 18638 4600 18694
rect 4668 18638 4724 18694
rect 2808 18514 2864 18570
rect 2932 18514 2988 18570
rect 3056 18514 3112 18570
rect 3180 18514 3236 18570
rect 3304 18514 3360 18570
rect 3428 18514 3484 18570
rect 3552 18514 3608 18570
rect 3676 18514 3732 18570
rect 3800 18514 3856 18570
rect 3924 18514 3980 18570
rect 4048 18514 4104 18570
rect 4172 18514 4228 18570
rect 4296 18514 4352 18570
rect 4420 18514 4476 18570
rect 4544 18514 4600 18570
rect 4668 18514 4724 18570
rect 2808 18390 2864 18446
rect 2932 18390 2988 18446
rect 3056 18390 3112 18446
rect 3180 18390 3236 18446
rect 3304 18390 3360 18446
rect 3428 18390 3484 18446
rect 3552 18390 3608 18446
rect 3676 18390 3732 18446
rect 3800 18390 3856 18446
rect 3924 18390 3980 18446
rect 4048 18390 4104 18446
rect 4172 18390 4228 18446
rect 4296 18390 4352 18446
rect 4420 18390 4476 18446
rect 4544 18390 4600 18446
rect 4668 18390 4724 18446
rect 2808 18266 2864 18322
rect 2932 18266 2988 18322
rect 3056 18266 3112 18322
rect 3180 18266 3236 18322
rect 3304 18266 3360 18322
rect 3428 18266 3484 18322
rect 3552 18266 3608 18322
rect 3676 18266 3732 18322
rect 3800 18266 3856 18322
rect 3924 18266 3980 18322
rect 4048 18266 4104 18322
rect 4172 18266 4228 18322
rect 4296 18266 4352 18322
rect 4420 18266 4476 18322
rect 4544 18266 4600 18322
rect 4668 18266 4724 18322
rect 2808 18142 2864 18198
rect 2932 18142 2988 18198
rect 3056 18142 3112 18198
rect 3180 18142 3236 18198
rect 3304 18142 3360 18198
rect 3428 18142 3484 18198
rect 3552 18142 3608 18198
rect 3676 18142 3732 18198
rect 3800 18142 3856 18198
rect 3924 18142 3980 18198
rect 4048 18142 4104 18198
rect 4172 18142 4228 18198
rect 4296 18142 4352 18198
rect 4420 18142 4476 18198
rect 4544 18142 4600 18198
rect 4668 18142 4724 18198
rect 2808 18018 2864 18074
rect 2932 18018 2988 18074
rect 3056 18018 3112 18074
rect 3180 18018 3236 18074
rect 3304 18018 3360 18074
rect 3428 18018 3484 18074
rect 3552 18018 3608 18074
rect 3676 18018 3732 18074
rect 3800 18018 3856 18074
rect 3924 18018 3980 18074
rect 4048 18018 4104 18074
rect 4172 18018 4228 18074
rect 4296 18018 4352 18074
rect 4420 18018 4476 18074
rect 4544 18018 4600 18074
rect 4668 18018 4724 18074
rect 2808 17894 2864 17950
rect 2932 17894 2988 17950
rect 3056 17894 3112 17950
rect 3180 17894 3236 17950
rect 3304 17894 3360 17950
rect 3428 17894 3484 17950
rect 3552 17894 3608 17950
rect 3676 17894 3732 17950
rect 3800 17894 3856 17950
rect 3924 17894 3980 17950
rect 4048 17894 4104 17950
rect 4172 17894 4228 17950
rect 4296 17894 4352 17950
rect 4420 17894 4476 17950
rect 4544 17894 4600 17950
rect 4668 17894 4724 17950
rect 2808 17770 2864 17826
rect 2932 17770 2988 17826
rect 3056 17770 3112 17826
rect 3180 17770 3236 17826
rect 3304 17770 3360 17826
rect 3428 17770 3484 17826
rect 3552 17770 3608 17826
rect 3676 17770 3732 17826
rect 3800 17770 3856 17826
rect 3924 17770 3980 17826
rect 4048 17770 4104 17826
rect 4172 17770 4228 17826
rect 4296 17770 4352 17826
rect 4420 17770 4476 17826
rect 4544 17770 4600 17826
rect 4668 17770 4724 17826
rect 2808 17646 2864 17702
rect 2932 17646 2988 17702
rect 3056 17646 3112 17702
rect 3180 17646 3236 17702
rect 3304 17646 3360 17702
rect 3428 17646 3484 17702
rect 3552 17646 3608 17702
rect 3676 17646 3732 17702
rect 3800 17646 3856 17702
rect 3924 17646 3980 17702
rect 4048 17646 4104 17702
rect 4172 17646 4228 17702
rect 4296 17646 4352 17702
rect 4420 17646 4476 17702
rect 4544 17646 4600 17702
rect 4668 17646 4724 17702
rect 5178 20498 5234 20554
rect 5302 20498 5358 20554
rect 5426 20498 5482 20554
rect 5550 20498 5606 20554
rect 5674 20498 5730 20554
rect 5798 20498 5854 20554
rect 5922 20498 5978 20554
rect 6046 20498 6102 20554
rect 6170 20498 6226 20554
rect 6294 20498 6350 20554
rect 6418 20498 6474 20554
rect 6542 20498 6598 20554
rect 6666 20498 6722 20554
rect 6790 20498 6846 20554
rect 6914 20498 6970 20554
rect 7038 20498 7094 20554
rect 5178 20374 5234 20430
rect 5302 20374 5358 20430
rect 5426 20374 5482 20430
rect 5550 20374 5606 20430
rect 5674 20374 5730 20430
rect 5798 20374 5854 20430
rect 5922 20374 5978 20430
rect 6046 20374 6102 20430
rect 6170 20374 6226 20430
rect 6294 20374 6350 20430
rect 6418 20374 6474 20430
rect 6542 20374 6598 20430
rect 6666 20374 6722 20430
rect 6790 20374 6846 20430
rect 6914 20374 6970 20430
rect 7038 20374 7094 20430
rect 5178 20250 5234 20306
rect 5302 20250 5358 20306
rect 5426 20250 5482 20306
rect 5550 20250 5606 20306
rect 5674 20250 5730 20306
rect 5798 20250 5854 20306
rect 5922 20250 5978 20306
rect 6046 20250 6102 20306
rect 6170 20250 6226 20306
rect 6294 20250 6350 20306
rect 6418 20250 6474 20306
rect 6542 20250 6598 20306
rect 6666 20250 6722 20306
rect 6790 20250 6846 20306
rect 6914 20250 6970 20306
rect 7038 20250 7094 20306
rect 5178 20126 5234 20182
rect 5302 20126 5358 20182
rect 5426 20126 5482 20182
rect 5550 20126 5606 20182
rect 5674 20126 5730 20182
rect 5798 20126 5854 20182
rect 5922 20126 5978 20182
rect 6046 20126 6102 20182
rect 6170 20126 6226 20182
rect 6294 20126 6350 20182
rect 6418 20126 6474 20182
rect 6542 20126 6598 20182
rect 6666 20126 6722 20182
rect 6790 20126 6846 20182
rect 6914 20126 6970 20182
rect 7038 20126 7094 20182
rect 5178 20002 5234 20058
rect 5302 20002 5358 20058
rect 5426 20002 5482 20058
rect 5550 20002 5606 20058
rect 5674 20002 5730 20058
rect 5798 20002 5854 20058
rect 5922 20002 5978 20058
rect 6046 20002 6102 20058
rect 6170 20002 6226 20058
rect 6294 20002 6350 20058
rect 6418 20002 6474 20058
rect 6542 20002 6598 20058
rect 6666 20002 6722 20058
rect 6790 20002 6846 20058
rect 6914 20002 6970 20058
rect 7038 20002 7094 20058
rect 5178 19878 5234 19934
rect 5302 19878 5358 19934
rect 5426 19878 5482 19934
rect 5550 19878 5606 19934
rect 5674 19878 5730 19934
rect 5798 19878 5854 19934
rect 5922 19878 5978 19934
rect 6046 19878 6102 19934
rect 6170 19878 6226 19934
rect 6294 19878 6350 19934
rect 6418 19878 6474 19934
rect 6542 19878 6598 19934
rect 6666 19878 6722 19934
rect 6790 19878 6846 19934
rect 6914 19878 6970 19934
rect 7038 19878 7094 19934
rect 5178 19754 5234 19810
rect 5302 19754 5358 19810
rect 5426 19754 5482 19810
rect 5550 19754 5606 19810
rect 5674 19754 5730 19810
rect 5798 19754 5854 19810
rect 5922 19754 5978 19810
rect 6046 19754 6102 19810
rect 6170 19754 6226 19810
rect 6294 19754 6350 19810
rect 6418 19754 6474 19810
rect 6542 19754 6598 19810
rect 6666 19754 6722 19810
rect 6790 19754 6846 19810
rect 6914 19754 6970 19810
rect 7038 19754 7094 19810
rect 5178 19630 5234 19686
rect 5302 19630 5358 19686
rect 5426 19630 5482 19686
rect 5550 19630 5606 19686
rect 5674 19630 5730 19686
rect 5798 19630 5854 19686
rect 5922 19630 5978 19686
rect 6046 19630 6102 19686
rect 6170 19630 6226 19686
rect 6294 19630 6350 19686
rect 6418 19630 6474 19686
rect 6542 19630 6598 19686
rect 6666 19630 6722 19686
rect 6790 19630 6846 19686
rect 6914 19630 6970 19686
rect 7038 19630 7094 19686
rect 5178 19506 5234 19562
rect 5302 19506 5358 19562
rect 5426 19506 5482 19562
rect 5550 19506 5606 19562
rect 5674 19506 5730 19562
rect 5798 19506 5854 19562
rect 5922 19506 5978 19562
rect 6046 19506 6102 19562
rect 6170 19506 6226 19562
rect 6294 19506 6350 19562
rect 6418 19506 6474 19562
rect 6542 19506 6598 19562
rect 6666 19506 6722 19562
rect 6790 19506 6846 19562
rect 6914 19506 6970 19562
rect 7038 19506 7094 19562
rect 5178 19382 5234 19438
rect 5302 19382 5358 19438
rect 5426 19382 5482 19438
rect 5550 19382 5606 19438
rect 5674 19382 5730 19438
rect 5798 19382 5854 19438
rect 5922 19382 5978 19438
rect 6046 19382 6102 19438
rect 6170 19382 6226 19438
rect 6294 19382 6350 19438
rect 6418 19382 6474 19438
rect 6542 19382 6598 19438
rect 6666 19382 6722 19438
rect 6790 19382 6846 19438
rect 6914 19382 6970 19438
rect 7038 19382 7094 19438
rect 5178 19258 5234 19314
rect 5302 19258 5358 19314
rect 5426 19258 5482 19314
rect 5550 19258 5606 19314
rect 5674 19258 5730 19314
rect 5798 19258 5854 19314
rect 5922 19258 5978 19314
rect 6046 19258 6102 19314
rect 6170 19258 6226 19314
rect 6294 19258 6350 19314
rect 6418 19258 6474 19314
rect 6542 19258 6598 19314
rect 6666 19258 6722 19314
rect 6790 19258 6846 19314
rect 6914 19258 6970 19314
rect 7038 19258 7094 19314
rect 5178 19134 5234 19190
rect 5302 19134 5358 19190
rect 5426 19134 5482 19190
rect 5550 19134 5606 19190
rect 5674 19134 5730 19190
rect 5798 19134 5854 19190
rect 5922 19134 5978 19190
rect 6046 19134 6102 19190
rect 6170 19134 6226 19190
rect 6294 19134 6350 19190
rect 6418 19134 6474 19190
rect 6542 19134 6598 19190
rect 6666 19134 6722 19190
rect 6790 19134 6846 19190
rect 6914 19134 6970 19190
rect 7038 19134 7094 19190
rect 5178 19010 5234 19066
rect 5302 19010 5358 19066
rect 5426 19010 5482 19066
rect 5550 19010 5606 19066
rect 5674 19010 5730 19066
rect 5798 19010 5854 19066
rect 5922 19010 5978 19066
rect 6046 19010 6102 19066
rect 6170 19010 6226 19066
rect 6294 19010 6350 19066
rect 6418 19010 6474 19066
rect 6542 19010 6598 19066
rect 6666 19010 6722 19066
rect 6790 19010 6846 19066
rect 6914 19010 6970 19066
rect 7038 19010 7094 19066
rect 5178 18886 5234 18942
rect 5302 18886 5358 18942
rect 5426 18886 5482 18942
rect 5550 18886 5606 18942
rect 5674 18886 5730 18942
rect 5798 18886 5854 18942
rect 5922 18886 5978 18942
rect 6046 18886 6102 18942
rect 6170 18886 6226 18942
rect 6294 18886 6350 18942
rect 6418 18886 6474 18942
rect 6542 18886 6598 18942
rect 6666 18886 6722 18942
rect 6790 18886 6846 18942
rect 6914 18886 6970 18942
rect 7038 18886 7094 18942
rect 5178 18762 5234 18818
rect 5302 18762 5358 18818
rect 5426 18762 5482 18818
rect 5550 18762 5606 18818
rect 5674 18762 5730 18818
rect 5798 18762 5854 18818
rect 5922 18762 5978 18818
rect 6046 18762 6102 18818
rect 6170 18762 6226 18818
rect 6294 18762 6350 18818
rect 6418 18762 6474 18818
rect 6542 18762 6598 18818
rect 6666 18762 6722 18818
rect 6790 18762 6846 18818
rect 6914 18762 6970 18818
rect 7038 18762 7094 18818
rect 5178 18638 5234 18694
rect 5302 18638 5358 18694
rect 5426 18638 5482 18694
rect 5550 18638 5606 18694
rect 5674 18638 5730 18694
rect 5798 18638 5854 18694
rect 5922 18638 5978 18694
rect 6046 18638 6102 18694
rect 6170 18638 6226 18694
rect 6294 18638 6350 18694
rect 6418 18638 6474 18694
rect 6542 18638 6598 18694
rect 6666 18638 6722 18694
rect 6790 18638 6846 18694
rect 6914 18638 6970 18694
rect 7038 18638 7094 18694
rect 5178 18514 5234 18570
rect 5302 18514 5358 18570
rect 5426 18514 5482 18570
rect 5550 18514 5606 18570
rect 5674 18514 5730 18570
rect 5798 18514 5854 18570
rect 5922 18514 5978 18570
rect 6046 18514 6102 18570
rect 6170 18514 6226 18570
rect 6294 18514 6350 18570
rect 6418 18514 6474 18570
rect 6542 18514 6598 18570
rect 6666 18514 6722 18570
rect 6790 18514 6846 18570
rect 6914 18514 6970 18570
rect 7038 18514 7094 18570
rect 5178 18390 5234 18446
rect 5302 18390 5358 18446
rect 5426 18390 5482 18446
rect 5550 18390 5606 18446
rect 5674 18390 5730 18446
rect 5798 18390 5854 18446
rect 5922 18390 5978 18446
rect 6046 18390 6102 18446
rect 6170 18390 6226 18446
rect 6294 18390 6350 18446
rect 6418 18390 6474 18446
rect 6542 18390 6598 18446
rect 6666 18390 6722 18446
rect 6790 18390 6846 18446
rect 6914 18390 6970 18446
rect 7038 18390 7094 18446
rect 5178 18266 5234 18322
rect 5302 18266 5358 18322
rect 5426 18266 5482 18322
rect 5550 18266 5606 18322
rect 5674 18266 5730 18322
rect 5798 18266 5854 18322
rect 5922 18266 5978 18322
rect 6046 18266 6102 18322
rect 6170 18266 6226 18322
rect 6294 18266 6350 18322
rect 6418 18266 6474 18322
rect 6542 18266 6598 18322
rect 6666 18266 6722 18322
rect 6790 18266 6846 18322
rect 6914 18266 6970 18322
rect 7038 18266 7094 18322
rect 5178 18142 5234 18198
rect 5302 18142 5358 18198
rect 5426 18142 5482 18198
rect 5550 18142 5606 18198
rect 5674 18142 5730 18198
rect 5798 18142 5854 18198
rect 5922 18142 5978 18198
rect 6046 18142 6102 18198
rect 6170 18142 6226 18198
rect 6294 18142 6350 18198
rect 6418 18142 6474 18198
rect 6542 18142 6598 18198
rect 6666 18142 6722 18198
rect 6790 18142 6846 18198
rect 6914 18142 6970 18198
rect 7038 18142 7094 18198
rect 5178 18018 5234 18074
rect 5302 18018 5358 18074
rect 5426 18018 5482 18074
rect 5550 18018 5606 18074
rect 5674 18018 5730 18074
rect 5798 18018 5854 18074
rect 5922 18018 5978 18074
rect 6046 18018 6102 18074
rect 6170 18018 6226 18074
rect 6294 18018 6350 18074
rect 6418 18018 6474 18074
rect 6542 18018 6598 18074
rect 6666 18018 6722 18074
rect 6790 18018 6846 18074
rect 6914 18018 6970 18074
rect 7038 18018 7094 18074
rect 5178 17894 5234 17950
rect 5302 17894 5358 17950
rect 5426 17894 5482 17950
rect 5550 17894 5606 17950
rect 5674 17894 5730 17950
rect 5798 17894 5854 17950
rect 5922 17894 5978 17950
rect 6046 17894 6102 17950
rect 6170 17894 6226 17950
rect 6294 17894 6350 17950
rect 6418 17894 6474 17950
rect 6542 17894 6598 17950
rect 6666 17894 6722 17950
rect 6790 17894 6846 17950
rect 6914 17894 6970 17950
rect 7038 17894 7094 17950
rect 5178 17770 5234 17826
rect 5302 17770 5358 17826
rect 5426 17770 5482 17826
rect 5550 17770 5606 17826
rect 5674 17770 5730 17826
rect 5798 17770 5854 17826
rect 5922 17770 5978 17826
rect 6046 17770 6102 17826
rect 6170 17770 6226 17826
rect 6294 17770 6350 17826
rect 6418 17770 6474 17826
rect 6542 17770 6598 17826
rect 6666 17770 6722 17826
rect 6790 17770 6846 17826
rect 6914 17770 6970 17826
rect 7038 17770 7094 17826
rect 5178 17646 5234 17702
rect 5302 17646 5358 17702
rect 5426 17646 5482 17702
rect 5550 17646 5606 17702
rect 5674 17646 5730 17702
rect 5798 17646 5854 17702
rect 5922 17646 5978 17702
rect 6046 17646 6102 17702
rect 6170 17646 6226 17702
rect 6294 17646 6350 17702
rect 6418 17646 6474 17702
rect 6542 17646 6598 17702
rect 6666 17646 6722 17702
rect 6790 17646 6846 17702
rect 6914 17646 6970 17702
rect 7038 17646 7094 17702
rect 7884 20498 7940 20554
rect 8008 20498 8064 20554
rect 8132 20498 8188 20554
rect 8256 20498 8312 20554
rect 8380 20498 8436 20554
rect 8504 20498 8560 20554
rect 8628 20498 8684 20554
rect 8752 20498 8808 20554
rect 8876 20498 8932 20554
rect 9000 20498 9056 20554
rect 9124 20498 9180 20554
rect 9248 20498 9304 20554
rect 9372 20498 9428 20554
rect 9496 20498 9552 20554
rect 9620 20498 9676 20554
rect 9744 20498 9800 20554
rect 7884 20374 7940 20430
rect 8008 20374 8064 20430
rect 8132 20374 8188 20430
rect 8256 20374 8312 20430
rect 8380 20374 8436 20430
rect 8504 20374 8560 20430
rect 8628 20374 8684 20430
rect 8752 20374 8808 20430
rect 8876 20374 8932 20430
rect 9000 20374 9056 20430
rect 9124 20374 9180 20430
rect 9248 20374 9304 20430
rect 9372 20374 9428 20430
rect 9496 20374 9552 20430
rect 9620 20374 9676 20430
rect 9744 20374 9800 20430
rect 7884 20250 7940 20306
rect 8008 20250 8064 20306
rect 8132 20250 8188 20306
rect 8256 20250 8312 20306
rect 8380 20250 8436 20306
rect 8504 20250 8560 20306
rect 8628 20250 8684 20306
rect 8752 20250 8808 20306
rect 8876 20250 8932 20306
rect 9000 20250 9056 20306
rect 9124 20250 9180 20306
rect 9248 20250 9304 20306
rect 9372 20250 9428 20306
rect 9496 20250 9552 20306
rect 9620 20250 9676 20306
rect 9744 20250 9800 20306
rect 7884 20126 7940 20182
rect 8008 20126 8064 20182
rect 8132 20126 8188 20182
rect 8256 20126 8312 20182
rect 8380 20126 8436 20182
rect 8504 20126 8560 20182
rect 8628 20126 8684 20182
rect 8752 20126 8808 20182
rect 8876 20126 8932 20182
rect 9000 20126 9056 20182
rect 9124 20126 9180 20182
rect 9248 20126 9304 20182
rect 9372 20126 9428 20182
rect 9496 20126 9552 20182
rect 9620 20126 9676 20182
rect 9744 20126 9800 20182
rect 7884 20002 7940 20058
rect 8008 20002 8064 20058
rect 8132 20002 8188 20058
rect 8256 20002 8312 20058
rect 8380 20002 8436 20058
rect 8504 20002 8560 20058
rect 8628 20002 8684 20058
rect 8752 20002 8808 20058
rect 8876 20002 8932 20058
rect 9000 20002 9056 20058
rect 9124 20002 9180 20058
rect 9248 20002 9304 20058
rect 9372 20002 9428 20058
rect 9496 20002 9552 20058
rect 9620 20002 9676 20058
rect 9744 20002 9800 20058
rect 7884 19878 7940 19934
rect 8008 19878 8064 19934
rect 8132 19878 8188 19934
rect 8256 19878 8312 19934
rect 8380 19878 8436 19934
rect 8504 19878 8560 19934
rect 8628 19878 8684 19934
rect 8752 19878 8808 19934
rect 8876 19878 8932 19934
rect 9000 19878 9056 19934
rect 9124 19878 9180 19934
rect 9248 19878 9304 19934
rect 9372 19878 9428 19934
rect 9496 19878 9552 19934
rect 9620 19878 9676 19934
rect 9744 19878 9800 19934
rect 7884 19754 7940 19810
rect 8008 19754 8064 19810
rect 8132 19754 8188 19810
rect 8256 19754 8312 19810
rect 8380 19754 8436 19810
rect 8504 19754 8560 19810
rect 8628 19754 8684 19810
rect 8752 19754 8808 19810
rect 8876 19754 8932 19810
rect 9000 19754 9056 19810
rect 9124 19754 9180 19810
rect 9248 19754 9304 19810
rect 9372 19754 9428 19810
rect 9496 19754 9552 19810
rect 9620 19754 9676 19810
rect 9744 19754 9800 19810
rect 7884 19630 7940 19686
rect 8008 19630 8064 19686
rect 8132 19630 8188 19686
rect 8256 19630 8312 19686
rect 8380 19630 8436 19686
rect 8504 19630 8560 19686
rect 8628 19630 8684 19686
rect 8752 19630 8808 19686
rect 8876 19630 8932 19686
rect 9000 19630 9056 19686
rect 9124 19630 9180 19686
rect 9248 19630 9304 19686
rect 9372 19630 9428 19686
rect 9496 19630 9552 19686
rect 9620 19630 9676 19686
rect 9744 19630 9800 19686
rect 7884 19506 7940 19562
rect 8008 19506 8064 19562
rect 8132 19506 8188 19562
rect 8256 19506 8312 19562
rect 8380 19506 8436 19562
rect 8504 19506 8560 19562
rect 8628 19506 8684 19562
rect 8752 19506 8808 19562
rect 8876 19506 8932 19562
rect 9000 19506 9056 19562
rect 9124 19506 9180 19562
rect 9248 19506 9304 19562
rect 9372 19506 9428 19562
rect 9496 19506 9552 19562
rect 9620 19506 9676 19562
rect 9744 19506 9800 19562
rect 7884 19382 7940 19438
rect 8008 19382 8064 19438
rect 8132 19382 8188 19438
rect 8256 19382 8312 19438
rect 8380 19382 8436 19438
rect 8504 19382 8560 19438
rect 8628 19382 8684 19438
rect 8752 19382 8808 19438
rect 8876 19382 8932 19438
rect 9000 19382 9056 19438
rect 9124 19382 9180 19438
rect 9248 19382 9304 19438
rect 9372 19382 9428 19438
rect 9496 19382 9552 19438
rect 9620 19382 9676 19438
rect 9744 19382 9800 19438
rect 7884 19258 7940 19314
rect 8008 19258 8064 19314
rect 8132 19258 8188 19314
rect 8256 19258 8312 19314
rect 8380 19258 8436 19314
rect 8504 19258 8560 19314
rect 8628 19258 8684 19314
rect 8752 19258 8808 19314
rect 8876 19258 8932 19314
rect 9000 19258 9056 19314
rect 9124 19258 9180 19314
rect 9248 19258 9304 19314
rect 9372 19258 9428 19314
rect 9496 19258 9552 19314
rect 9620 19258 9676 19314
rect 9744 19258 9800 19314
rect 7884 19134 7940 19190
rect 8008 19134 8064 19190
rect 8132 19134 8188 19190
rect 8256 19134 8312 19190
rect 8380 19134 8436 19190
rect 8504 19134 8560 19190
rect 8628 19134 8684 19190
rect 8752 19134 8808 19190
rect 8876 19134 8932 19190
rect 9000 19134 9056 19190
rect 9124 19134 9180 19190
rect 9248 19134 9304 19190
rect 9372 19134 9428 19190
rect 9496 19134 9552 19190
rect 9620 19134 9676 19190
rect 9744 19134 9800 19190
rect 7884 19010 7940 19066
rect 8008 19010 8064 19066
rect 8132 19010 8188 19066
rect 8256 19010 8312 19066
rect 8380 19010 8436 19066
rect 8504 19010 8560 19066
rect 8628 19010 8684 19066
rect 8752 19010 8808 19066
rect 8876 19010 8932 19066
rect 9000 19010 9056 19066
rect 9124 19010 9180 19066
rect 9248 19010 9304 19066
rect 9372 19010 9428 19066
rect 9496 19010 9552 19066
rect 9620 19010 9676 19066
rect 9744 19010 9800 19066
rect 7884 18886 7940 18942
rect 8008 18886 8064 18942
rect 8132 18886 8188 18942
rect 8256 18886 8312 18942
rect 8380 18886 8436 18942
rect 8504 18886 8560 18942
rect 8628 18886 8684 18942
rect 8752 18886 8808 18942
rect 8876 18886 8932 18942
rect 9000 18886 9056 18942
rect 9124 18886 9180 18942
rect 9248 18886 9304 18942
rect 9372 18886 9428 18942
rect 9496 18886 9552 18942
rect 9620 18886 9676 18942
rect 9744 18886 9800 18942
rect 7884 18762 7940 18818
rect 8008 18762 8064 18818
rect 8132 18762 8188 18818
rect 8256 18762 8312 18818
rect 8380 18762 8436 18818
rect 8504 18762 8560 18818
rect 8628 18762 8684 18818
rect 8752 18762 8808 18818
rect 8876 18762 8932 18818
rect 9000 18762 9056 18818
rect 9124 18762 9180 18818
rect 9248 18762 9304 18818
rect 9372 18762 9428 18818
rect 9496 18762 9552 18818
rect 9620 18762 9676 18818
rect 9744 18762 9800 18818
rect 7884 18638 7940 18694
rect 8008 18638 8064 18694
rect 8132 18638 8188 18694
rect 8256 18638 8312 18694
rect 8380 18638 8436 18694
rect 8504 18638 8560 18694
rect 8628 18638 8684 18694
rect 8752 18638 8808 18694
rect 8876 18638 8932 18694
rect 9000 18638 9056 18694
rect 9124 18638 9180 18694
rect 9248 18638 9304 18694
rect 9372 18638 9428 18694
rect 9496 18638 9552 18694
rect 9620 18638 9676 18694
rect 9744 18638 9800 18694
rect 7884 18514 7940 18570
rect 8008 18514 8064 18570
rect 8132 18514 8188 18570
rect 8256 18514 8312 18570
rect 8380 18514 8436 18570
rect 8504 18514 8560 18570
rect 8628 18514 8684 18570
rect 8752 18514 8808 18570
rect 8876 18514 8932 18570
rect 9000 18514 9056 18570
rect 9124 18514 9180 18570
rect 9248 18514 9304 18570
rect 9372 18514 9428 18570
rect 9496 18514 9552 18570
rect 9620 18514 9676 18570
rect 9744 18514 9800 18570
rect 7884 18390 7940 18446
rect 8008 18390 8064 18446
rect 8132 18390 8188 18446
rect 8256 18390 8312 18446
rect 8380 18390 8436 18446
rect 8504 18390 8560 18446
rect 8628 18390 8684 18446
rect 8752 18390 8808 18446
rect 8876 18390 8932 18446
rect 9000 18390 9056 18446
rect 9124 18390 9180 18446
rect 9248 18390 9304 18446
rect 9372 18390 9428 18446
rect 9496 18390 9552 18446
rect 9620 18390 9676 18446
rect 9744 18390 9800 18446
rect 7884 18266 7940 18322
rect 8008 18266 8064 18322
rect 8132 18266 8188 18322
rect 8256 18266 8312 18322
rect 8380 18266 8436 18322
rect 8504 18266 8560 18322
rect 8628 18266 8684 18322
rect 8752 18266 8808 18322
rect 8876 18266 8932 18322
rect 9000 18266 9056 18322
rect 9124 18266 9180 18322
rect 9248 18266 9304 18322
rect 9372 18266 9428 18322
rect 9496 18266 9552 18322
rect 9620 18266 9676 18322
rect 9744 18266 9800 18322
rect 7884 18142 7940 18198
rect 8008 18142 8064 18198
rect 8132 18142 8188 18198
rect 8256 18142 8312 18198
rect 8380 18142 8436 18198
rect 8504 18142 8560 18198
rect 8628 18142 8684 18198
rect 8752 18142 8808 18198
rect 8876 18142 8932 18198
rect 9000 18142 9056 18198
rect 9124 18142 9180 18198
rect 9248 18142 9304 18198
rect 9372 18142 9428 18198
rect 9496 18142 9552 18198
rect 9620 18142 9676 18198
rect 9744 18142 9800 18198
rect 7884 18018 7940 18074
rect 8008 18018 8064 18074
rect 8132 18018 8188 18074
rect 8256 18018 8312 18074
rect 8380 18018 8436 18074
rect 8504 18018 8560 18074
rect 8628 18018 8684 18074
rect 8752 18018 8808 18074
rect 8876 18018 8932 18074
rect 9000 18018 9056 18074
rect 9124 18018 9180 18074
rect 9248 18018 9304 18074
rect 9372 18018 9428 18074
rect 9496 18018 9552 18074
rect 9620 18018 9676 18074
rect 9744 18018 9800 18074
rect 7884 17894 7940 17950
rect 8008 17894 8064 17950
rect 8132 17894 8188 17950
rect 8256 17894 8312 17950
rect 8380 17894 8436 17950
rect 8504 17894 8560 17950
rect 8628 17894 8684 17950
rect 8752 17894 8808 17950
rect 8876 17894 8932 17950
rect 9000 17894 9056 17950
rect 9124 17894 9180 17950
rect 9248 17894 9304 17950
rect 9372 17894 9428 17950
rect 9496 17894 9552 17950
rect 9620 17894 9676 17950
rect 9744 17894 9800 17950
rect 7884 17770 7940 17826
rect 8008 17770 8064 17826
rect 8132 17770 8188 17826
rect 8256 17770 8312 17826
rect 8380 17770 8436 17826
rect 8504 17770 8560 17826
rect 8628 17770 8684 17826
rect 8752 17770 8808 17826
rect 8876 17770 8932 17826
rect 9000 17770 9056 17826
rect 9124 17770 9180 17826
rect 9248 17770 9304 17826
rect 9372 17770 9428 17826
rect 9496 17770 9552 17826
rect 9620 17770 9676 17826
rect 9744 17770 9800 17826
rect 7884 17646 7940 17702
rect 8008 17646 8064 17702
rect 8132 17646 8188 17702
rect 8256 17646 8312 17702
rect 8380 17646 8436 17702
rect 8504 17646 8560 17702
rect 8628 17646 8684 17702
rect 8752 17646 8808 17702
rect 8876 17646 8932 17702
rect 9000 17646 9056 17702
rect 9124 17646 9180 17702
rect 9248 17646 9304 17702
rect 9372 17646 9428 17702
rect 9496 17646 9552 17702
rect 9620 17646 9676 17702
rect 9744 17646 9800 17702
rect 10254 20498 10310 20554
rect 10378 20498 10434 20554
rect 10502 20498 10558 20554
rect 10626 20498 10682 20554
rect 10750 20498 10806 20554
rect 10874 20498 10930 20554
rect 10998 20498 11054 20554
rect 11122 20498 11178 20554
rect 11246 20498 11302 20554
rect 11370 20498 11426 20554
rect 11494 20498 11550 20554
rect 11618 20498 11674 20554
rect 11742 20498 11798 20554
rect 11866 20498 11922 20554
rect 11990 20498 12046 20554
rect 12114 20498 12170 20554
rect 10254 20374 10310 20430
rect 10378 20374 10434 20430
rect 10502 20374 10558 20430
rect 10626 20374 10682 20430
rect 10750 20374 10806 20430
rect 10874 20374 10930 20430
rect 10998 20374 11054 20430
rect 11122 20374 11178 20430
rect 11246 20374 11302 20430
rect 11370 20374 11426 20430
rect 11494 20374 11550 20430
rect 11618 20374 11674 20430
rect 11742 20374 11798 20430
rect 11866 20374 11922 20430
rect 11990 20374 12046 20430
rect 12114 20374 12170 20430
rect 10254 20250 10310 20306
rect 10378 20250 10434 20306
rect 10502 20250 10558 20306
rect 10626 20250 10682 20306
rect 10750 20250 10806 20306
rect 10874 20250 10930 20306
rect 10998 20250 11054 20306
rect 11122 20250 11178 20306
rect 11246 20250 11302 20306
rect 11370 20250 11426 20306
rect 11494 20250 11550 20306
rect 11618 20250 11674 20306
rect 11742 20250 11798 20306
rect 11866 20250 11922 20306
rect 11990 20250 12046 20306
rect 12114 20250 12170 20306
rect 10254 20126 10310 20182
rect 10378 20126 10434 20182
rect 10502 20126 10558 20182
rect 10626 20126 10682 20182
rect 10750 20126 10806 20182
rect 10874 20126 10930 20182
rect 10998 20126 11054 20182
rect 11122 20126 11178 20182
rect 11246 20126 11302 20182
rect 11370 20126 11426 20182
rect 11494 20126 11550 20182
rect 11618 20126 11674 20182
rect 11742 20126 11798 20182
rect 11866 20126 11922 20182
rect 11990 20126 12046 20182
rect 12114 20126 12170 20182
rect 10254 20002 10310 20058
rect 10378 20002 10434 20058
rect 10502 20002 10558 20058
rect 10626 20002 10682 20058
rect 10750 20002 10806 20058
rect 10874 20002 10930 20058
rect 10998 20002 11054 20058
rect 11122 20002 11178 20058
rect 11246 20002 11302 20058
rect 11370 20002 11426 20058
rect 11494 20002 11550 20058
rect 11618 20002 11674 20058
rect 11742 20002 11798 20058
rect 11866 20002 11922 20058
rect 11990 20002 12046 20058
rect 12114 20002 12170 20058
rect 10254 19878 10310 19934
rect 10378 19878 10434 19934
rect 10502 19878 10558 19934
rect 10626 19878 10682 19934
rect 10750 19878 10806 19934
rect 10874 19878 10930 19934
rect 10998 19878 11054 19934
rect 11122 19878 11178 19934
rect 11246 19878 11302 19934
rect 11370 19878 11426 19934
rect 11494 19878 11550 19934
rect 11618 19878 11674 19934
rect 11742 19878 11798 19934
rect 11866 19878 11922 19934
rect 11990 19878 12046 19934
rect 12114 19878 12170 19934
rect 10254 19754 10310 19810
rect 10378 19754 10434 19810
rect 10502 19754 10558 19810
rect 10626 19754 10682 19810
rect 10750 19754 10806 19810
rect 10874 19754 10930 19810
rect 10998 19754 11054 19810
rect 11122 19754 11178 19810
rect 11246 19754 11302 19810
rect 11370 19754 11426 19810
rect 11494 19754 11550 19810
rect 11618 19754 11674 19810
rect 11742 19754 11798 19810
rect 11866 19754 11922 19810
rect 11990 19754 12046 19810
rect 12114 19754 12170 19810
rect 10254 19630 10310 19686
rect 10378 19630 10434 19686
rect 10502 19630 10558 19686
rect 10626 19630 10682 19686
rect 10750 19630 10806 19686
rect 10874 19630 10930 19686
rect 10998 19630 11054 19686
rect 11122 19630 11178 19686
rect 11246 19630 11302 19686
rect 11370 19630 11426 19686
rect 11494 19630 11550 19686
rect 11618 19630 11674 19686
rect 11742 19630 11798 19686
rect 11866 19630 11922 19686
rect 11990 19630 12046 19686
rect 12114 19630 12170 19686
rect 10254 19506 10310 19562
rect 10378 19506 10434 19562
rect 10502 19506 10558 19562
rect 10626 19506 10682 19562
rect 10750 19506 10806 19562
rect 10874 19506 10930 19562
rect 10998 19506 11054 19562
rect 11122 19506 11178 19562
rect 11246 19506 11302 19562
rect 11370 19506 11426 19562
rect 11494 19506 11550 19562
rect 11618 19506 11674 19562
rect 11742 19506 11798 19562
rect 11866 19506 11922 19562
rect 11990 19506 12046 19562
rect 12114 19506 12170 19562
rect 10254 19382 10310 19438
rect 10378 19382 10434 19438
rect 10502 19382 10558 19438
rect 10626 19382 10682 19438
rect 10750 19382 10806 19438
rect 10874 19382 10930 19438
rect 10998 19382 11054 19438
rect 11122 19382 11178 19438
rect 11246 19382 11302 19438
rect 11370 19382 11426 19438
rect 11494 19382 11550 19438
rect 11618 19382 11674 19438
rect 11742 19382 11798 19438
rect 11866 19382 11922 19438
rect 11990 19382 12046 19438
rect 12114 19382 12170 19438
rect 10254 19258 10310 19314
rect 10378 19258 10434 19314
rect 10502 19258 10558 19314
rect 10626 19258 10682 19314
rect 10750 19258 10806 19314
rect 10874 19258 10930 19314
rect 10998 19258 11054 19314
rect 11122 19258 11178 19314
rect 11246 19258 11302 19314
rect 11370 19258 11426 19314
rect 11494 19258 11550 19314
rect 11618 19258 11674 19314
rect 11742 19258 11798 19314
rect 11866 19258 11922 19314
rect 11990 19258 12046 19314
rect 12114 19258 12170 19314
rect 10254 19134 10310 19190
rect 10378 19134 10434 19190
rect 10502 19134 10558 19190
rect 10626 19134 10682 19190
rect 10750 19134 10806 19190
rect 10874 19134 10930 19190
rect 10998 19134 11054 19190
rect 11122 19134 11178 19190
rect 11246 19134 11302 19190
rect 11370 19134 11426 19190
rect 11494 19134 11550 19190
rect 11618 19134 11674 19190
rect 11742 19134 11798 19190
rect 11866 19134 11922 19190
rect 11990 19134 12046 19190
rect 12114 19134 12170 19190
rect 10254 19010 10310 19066
rect 10378 19010 10434 19066
rect 10502 19010 10558 19066
rect 10626 19010 10682 19066
rect 10750 19010 10806 19066
rect 10874 19010 10930 19066
rect 10998 19010 11054 19066
rect 11122 19010 11178 19066
rect 11246 19010 11302 19066
rect 11370 19010 11426 19066
rect 11494 19010 11550 19066
rect 11618 19010 11674 19066
rect 11742 19010 11798 19066
rect 11866 19010 11922 19066
rect 11990 19010 12046 19066
rect 12114 19010 12170 19066
rect 10254 18886 10310 18942
rect 10378 18886 10434 18942
rect 10502 18886 10558 18942
rect 10626 18886 10682 18942
rect 10750 18886 10806 18942
rect 10874 18886 10930 18942
rect 10998 18886 11054 18942
rect 11122 18886 11178 18942
rect 11246 18886 11302 18942
rect 11370 18886 11426 18942
rect 11494 18886 11550 18942
rect 11618 18886 11674 18942
rect 11742 18886 11798 18942
rect 11866 18886 11922 18942
rect 11990 18886 12046 18942
rect 12114 18886 12170 18942
rect 10254 18762 10310 18818
rect 10378 18762 10434 18818
rect 10502 18762 10558 18818
rect 10626 18762 10682 18818
rect 10750 18762 10806 18818
rect 10874 18762 10930 18818
rect 10998 18762 11054 18818
rect 11122 18762 11178 18818
rect 11246 18762 11302 18818
rect 11370 18762 11426 18818
rect 11494 18762 11550 18818
rect 11618 18762 11674 18818
rect 11742 18762 11798 18818
rect 11866 18762 11922 18818
rect 11990 18762 12046 18818
rect 12114 18762 12170 18818
rect 10254 18638 10310 18694
rect 10378 18638 10434 18694
rect 10502 18638 10558 18694
rect 10626 18638 10682 18694
rect 10750 18638 10806 18694
rect 10874 18638 10930 18694
rect 10998 18638 11054 18694
rect 11122 18638 11178 18694
rect 11246 18638 11302 18694
rect 11370 18638 11426 18694
rect 11494 18638 11550 18694
rect 11618 18638 11674 18694
rect 11742 18638 11798 18694
rect 11866 18638 11922 18694
rect 11990 18638 12046 18694
rect 12114 18638 12170 18694
rect 10254 18514 10310 18570
rect 10378 18514 10434 18570
rect 10502 18514 10558 18570
rect 10626 18514 10682 18570
rect 10750 18514 10806 18570
rect 10874 18514 10930 18570
rect 10998 18514 11054 18570
rect 11122 18514 11178 18570
rect 11246 18514 11302 18570
rect 11370 18514 11426 18570
rect 11494 18514 11550 18570
rect 11618 18514 11674 18570
rect 11742 18514 11798 18570
rect 11866 18514 11922 18570
rect 11990 18514 12046 18570
rect 12114 18514 12170 18570
rect 10254 18390 10310 18446
rect 10378 18390 10434 18446
rect 10502 18390 10558 18446
rect 10626 18390 10682 18446
rect 10750 18390 10806 18446
rect 10874 18390 10930 18446
rect 10998 18390 11054 18446
rect 11122 18390 11178 18446
rect 11246 18390 11302 18446
rect 11370 18390 11426 18446
rect 11494 18390 11550 18446
rect 11618 18390 11674 18446
rect 11742 18390 11798 18446
rect 11866 18390 11922 18446
rect 11990 18390 12046 18446
rect 12114 18390 12170 18446
rect 10254 18266 10310 18322
rect 10378 18266 10434 18322
rect 10502 18266 10558 18322
rect 10626 18266 10682 18322
rect 10750 18266 10806 18322
rect 10874 18266 10930 18322
rect 10998 18266 11054 18322
rect 11122 18266 11178 18322
rect 11246 18266 11302 18322
rect 11370 18266 11426 18322
rect 11494 18266 11550 18322
rect 11618 18266 11674 18322
rect 11742 18266 11798 18322
rect 11866 18266 11922 18322
rect 11990 18266 12046 18322
rect 12114 18266 12170 18322
rect 10254 18142 10310 18198
rect 10378 18142 10434 18198
rect 10502 18142 10558 18198
rect 10626 18142 10682 18198
rect 10750 18142 10806 18198
rect 10874 18142 10930 18198
rect 10998 18142 11054 18198
rect 11122 18142 11178 18198
rect 11246 18142 11302 18198
rect 11370 18142 11426 18198
rect 11494 18142 11550 18198
rect 11618 18142 11674 18198
rect 11742 18142 11798 18198
rect 11866 18142 11922 18198
rect 11990 18142 12046 18198
rect 12114 18142 12170 18198
rect 10254 18018 10310 18074
rect 10378 18018 10434 18074
rect 10502 18018 10558 18074
rect 10626 18018 10682 18074
rect 10750 18018 10806 18074
rect 10874 18018 10930 18074
rect 10998 18018 11054 18074
rect 11122 18018 11178 18074
rect 11246 18018 11302 18074
rect 11370 18018 11426 18074
rect 11494 18018 11550 18074
rect 11618 18018 11674 18074
rect 11742 18018 11798 18074
rect 11866 18018 11922 18074
rect 11990 18018 12046 18074
rect 12114 18018 12170 18074
rect 10254 17894 10310 17950
rect 10378 17894 10434 17950
rect 10502 17894 10558 17950
rect 10626 17894 10682 17950
rect 10750 17894 10806 17950
rect 10874 17894 10930 17950
rect 10998 17894 11054 17950
rect 11122 17894 11178 17950
rect 11246 17894 11302 17950
rect 11370 17894 11426 17950
rect 11494 17894 11550 17950
rect 11618 17894 11674 17950
rect 11742 17894 11798 17950
rect 11866 17894 11922 17950
rect 11990 17894 12046 17950
rect 12114 17894 12170 17950
rect 10254 17770 10310 17826
rect 10378 17770 10434 17826
rect 10502 17770 10558 17826
rect 10626 17770 10682 17826
rect 10750 17770 10806 17826
rect 10874 17770 10930 17826
rect 10998 17770 11054 17826
rect 11122 17770 11178 17826
rect 11246 17770 11302 17826
rect 11370 17770 11426 17826
rect 11494 17770 11550 17826
rect 11618 17770 11674 17826
rect 11742 17770 11798 17826
rect 11866 17770 11922 17826
rect 11990 17770 12046 17826
rect 12114 17770 12170 17826
rect 10254 17646 10310 17702
rect 10378 17646 10434 17702
rect 10502 17646 10558 17702
rect 10626 17646 10682 17702
rect 10750 17646 10806 17702
rect 10874 17646 10930 17702
rect 10998 17646 11054 17702
rect 11122 17646 11178 17702
rect 11246 17646 11302 17702
rect 11370 17646 11426 17702
rect 11494 17646 11550 17702
rect 11618 17646 11674 17702
rect 11742 17646 11798 17702
rect 11866 17646 11922 17702
rect 11990 17646 12046 17702
rect 12114 17646 12170 17702
rect 12871 20498 12927 20554
rect 12995 20498 13051 20554
rect 13119 20498 13175 20554
rect 13243 20498 13299 20554
rect 13367 20498 13423 20554
rect 13491 20498 13547 20554
rect 13615 20498 13671 20554
rect 13739 20498 13795 20554
rect 13863 20498 13919 20554
rect 13987 20498 14043 20554
rect 14111 20498 14167 20554
rect 14235 20498 14291 20554
rect 14359 20498 14415 20554
rect 14483 20498 14539 20554
rect 14607 20498 14663 20554
rect 12871 20374 12927 20430
rect 12995 20374 13051 20430
rect 13119 20374 13175 20430
rect 13243 20374 13299 20430
rect 13367 20374 13423 20430
rect 13491 20374 13547 20430
rect 13615 20374 13671 20430
rect 13739 20374 13795 20430
rect 13863 20374 13919 20430
rect 13987 20374 14043 20430
rect 14111 20374 14167 20430
rect 14235 20374 14291 20430
rect 14359 20374 14415 20430
rect 14483 20374 14539 20430
rect 14607 20374 14663 20430
rect 12871 20250 12927 20306
rect 12995 20250 13051 20306
rect 13119 20250 13175 20306
rect 13243 20250 13299 20306
rect 13367 20250 13423 20306
rect 13491 20250 13547 20306
rect 13615 20250 13671 20306
rect 13739 20250 13795 20306
rect 13863 20250 13919 20306
rect 13987 20250 14043 20306
rect 14111 20250 14167 20306
rect 14235 20250 14291 20306
rect 14359 20250 14415 20306
rect 14483 20250 14539 20306
rect 14607 20250 14663 20306
rect 12871 20126 12927 20182
rect 12995 20126 13051 20182
rect 13119 20126 13175 20182
rect 13243 20126 13299 20182
rect 13367 20126 13423 20182
rect 13491 20126 13547 20182
rect 13615 20126 13671 20182
rect 13739 20126 13795 20182
rect 13863 20126 13919 20182
rect 13987 20126 14043 20182
rect 14111 20126 14167 20182
rect 14235 20126 14291 20182
rect 14359 20126 14415 20182
rect 14483 20126 14539 20182
rect 14607 20126 14663 20182
rect 12871 20002 12927 20058
rect 12995 20002 13051 20058
rect 13119 20002 13175 20058
rect 13243 20002 13299 20058
rect 13367 20002 13423 20058
rect 13491 20002 13547 20058
rect 13615 20002 13671 20058
rect 13739 20002 13795 20058
rect 13863 20002 13919 20058
rect 13987 20002 14043 20058
rect 14111 20002 14167 20058
rect 14235 20002 14291 20058
rect 14359 20002 14415 20058
rect 14483 20002 14539 20058
rect 14607 20002 14663 20058
rect 12871 19878 12927 19934
rect 12995 19878 13051 19934
rect 13119 19878 13175 19934
rect 13243 19878 13299 19934
rect 13367 19878 13423 19934
rect 13491 19878 13547 19934
rect 13615 19878 13671 19934
rect 13739 19878 13795 19934
rect 13863 19878 13919 19934
rect 13987 19878 14043 19934
rect 14111 19878 14167 19934
rect 14235 19878 14291 19934
rect 14359 19878 14415 19934
rect 14483 19878 14539 19934
rect 14607 19878 14663 19934
rect 12871 19754 12927 19810
rect 12995 19754 13051 19810
rect 13119 19754 13175 19810
rect 13243 19754 13299 19810
rect 13367 19754 13423 19810
rect 13491 19754 13547 19810
rect 13615 19754 13671 19810
rect 13739 19754 13795 19810
rect 13863 19754 13919 19810
rect 13987 19754 14043 19810
rect 14111 19754 14167 19810
rect 14235 19754 14291 19810
rect 14359 19754 14415 19810
rect 14483 19754 14539 19810
rect 14607 19754 14663 19810
rect 12871 19630 12927 19686
rect 12995 19630 13051 19686
rect 13119 19630 13175 19686
rect 13243 19630 13299 19686
rect 13367 19630 13423 19686
rect 13491 19630 13547 19686
rect 13615 19630 13671 19686
rect 13739 19630 13795 19686
rect 13863 19630 13919 19686
rect 13987 19630 14043 19686
rect 14111 19630 14167 19686
rect 14235 19630 14291 19686
rect 14359 19630 14415 19686
rect 14483 19630 14539 19686
rect 14607 19630 14663 19686
rect 12871 19506 12927 19562
rect 12995 19506 13051 19562
rect 13119 19506 13175 19562
rect 13243 19506 13299 19562
rect 13367 19506 13423 19562
rect 13491 19506 13547 19562
rect 13615 19506 13671 19562
rect 13739 19506 13795 19562
rect 13863 19506 13919 19562
rect 13987 19506 14043 19562
rect 14111 19506 14167 19562
rect 14235 19506 14291 19562
rect 14359 19506 14415 19562
rect 14483 19506 14539 19562
rect 14607 19506 14663 19562
rect 12871 19382 12927 19438
rect 12995 19382 13051 19438
rect 13119 19382 13175 19438
rect 13243 19382 13299 19438
rect 13367 19382 13423 19438
rect 13491 19382 13547 19438
rect 13615 19382 13671 19438
rect 13739 19382 13795 19438
rect 13863 19382 13919 19438
rect 13987 19382 14043 19438
rect 14111 19382 14167 19438
rect 14235 19382 14291 19438
rect 14359 19382 14415 19438
rect 14483 19382 14539 19438
rect 14607 19382 14663 19438
rect 12871 19258 12927 19314
rect 12995 19258 13051 19314
rect 13119 19258 13175 19314
rect 13243 19258 13299 19314
rect 13367 19258 13423 19314
rect 13491 19258 13547 19314
rect 13615 19258 13671 19314
rect 13739 19258 13795 19314
rect 13863 19258 13919 19314
rect 13987 19258 14043 19314
rect 14111 19258 14167 19314
rect 14235 19258 14291 19314
rect 14359 19258 14415 19314
rect 14483 19258 14539 19314
rect 14607 19258 14663 19314
rect 12871 19134 12927 19190
rect 12995 19134 13051 19190
rect 13119 19134 13175 19190
rect 13243 19134 13299 19190
rect 13367 19134 13423 19190
rect 13491 19134 13547 19190
rect 13615 19134 13671 19190
rect 13739 19134 13795 19190
rect 13863 19134 13919 19190
rect 13987 19134 14043 19190
rect 14111 19134 14167 19190
rect 14235 19134 14291 19190
rect 14359 19134 14415 19190
rect 14483 19134 14539 19190
rect 14607 19134 14663 19190
rect 12871 19010 12927 19066
rect 12995 19010 13051 19066
rect 13119 19010 13175 19066
rect 13243 19010 13299 19066
rect 13367 19010 13423 19066
rect 13491 19010 13547 19066
rect 13615 19010 13671 19066
rect 13739 19010 13795 19066
rect 13863 19010 13919 19066
rect 13987 19010 14043 19066
rect 14111 19010 14167 19066
rect 14235 19010 14291 19066
rect 14359 19010 14415 19066
rect 14483 19010 14539 19066
rect 14607 19010 14663 19066
rect 12871 18886 12927 18942
rect 12995 18886 13051 18942
rect 13119 18886 13175 18942
rect 13243 18886 13299 18942
rect 13367 18886 13423 18942
rect 13491 18886 13547 18942
rect 13615 18886 13671 18942
rect 13739 18886 13795 18942
rect 13863 18886 13919 18942
rect 13987 18886 14043 18942
rect 14111 18886 14167 18942
rect 14235 18886 14291 18942
rect 14359 18886 14415 18942
rect 14483 18886 14539 18942
rect 14607 18886 14663 18942
rect 12871 18762 12927 18818
rect 12995 18762 13051 18818
rect 13119 18762 13175 18818
rect 13243 18762 13299 18818
rect 13367 18762 13423 18818
rect 13491 18762 13547 18818
rect 13615 18762 13671 18818
rect 13739 18762 13795 18818
rect 13863 18762 13919 18818
rect 13987 18762 14043 18818
rect 14111 18762 14167 18818
rect 14235 18762 14291 18818
rect 14359 18762 14415 18818
rect 14483 18762 14539 18818
rect 14607 18762 14663 18818
rect 12871 18638 12927 18694
rect 12995 18638 13051 18694
rect 13119 18638 13175 18694
rect 13243 18638 13299 18694
rect 13367 18638 13423 18694
rect 13491 18638 13547 18694
rect 13615 18638 13671 18694
rect 13739 18638 13795 18694
rect 13863 18638 13919 18694
rect 13987 18638 14043 18694
rect 14111 18638 14167 18694
rect 14235 18638 14291 18694
rect 14359 18638 14415 18694
rect 14483 18638 14539 18694
rect 14607 18638 14663 18694
rect 12871 18514 12927 18570
rect 12995 18514 13051 18570
rect 13119 18514 13175 18570
rect 13243 18514 13299 18570
rect 13367 18514 13423 18570
rect 13491 18514 13547 18570
rect 13615 18514 13671 18570
rect 13739 18514 13795 18570
rect 13863 18514 13919 18570
rect 13987 18514 14043 18570
rect 14111 18514 14167 18570
rect 14235 18514 14291 18570
rect 14359 18514 14415 18570
rect 14483 18514 14539 18570
rect 14607 18514 14663 18570
rect 12871 18390 12927 18446
rect 12995 18390 13051 18446
rect 13119 18390 13175 18446
rect 13243 18390 13299 18446
rect 13367 18390 13423 18446
rect 13491 18390 13547 18446
rect 13615 18390 13671 18446
rect 13739 18390 13795 18446
rect 13863 18390 13919 18446
rect 13987 18390 14043 18446
rect 14111 18390 14167 18446
rect 14235 18390 14291 18446
rect 14359 18390 14415 18446
rect 14483 18390 14539 18446
rect 14607 18390 14663 18446
rect 12871 18266 12927 18322
rect 12995 18266 13051 18322
rect 13119 18266 13175 18322
rect 13243 18266 13299 18322
rect 13367 18266 13423 18322
rect 13491 18266 13547 18322
rect 13615 18266 13671 18322
rect 13739 18266 13795 18322
rect 13863 18266 13919 18322
rect 13987 18266 14043 18322
rect 14111 18266 14167 18322
rect 14235 18266 14291 18322
rect 14359 18266 14415 18322
rect 14483 18266 14539 18322
rect 14607 18266 14663 18322
rect 12871 18142 12927 18198
rect 12995 18142 13051 18198
rect 13119 18142 13175 18198
rect 13243 18142 13299 18198
rect 13367 18142 13423 18198
rect 13491 18142 13547 18198
rect 13615 18142 13671 18198
rect 13739 18142 13795 18198
rect 13863 18142 13919 18198
rect 13987 18142 14043 18198
rect 14111 18142 14167 18198
rect 14235 18142 14291 18198
rect 14359 18142 14415 18198
rect 14483 18142 14539 18198
rect 14607 18142 14663 18198
rect 12871 18018 12927 18074
rect 12995 18018 13051 18074
rect 13119 18018 13175 18074
rect 13243 18018 13299 18074
rect 13367 18018 13423 18074
rect 13491 18018 13547 18074
rect 13615 18018 13671 18074
rect 13739 18018 13795 18074
rect 13863 18018 13919 18074
rect 13987 18018 14043 18074
rect 14111 18018 14167 18074
rect 14235 18018 14291 18074
rect 14359 18018 14415 18074
rect 14483 18018 14539 18074
rect 14607 18018 14663 18074
rect 12871 17894 12927 17950
rect 12995 17894 13051 17950
rect 13119 17894 13175 17950
rect 13243 17894 13299 17950
rect 13367 17894 13423 17950
rect 13491 17894 13547 17950
rect 13615 17894 13671 17950
rect 13739 17894 13795 17950
rect 13863 17894 13919 17950
rect 13987 17894 14043 17950
rect 14111 17894 14167 17950
rect 14235 17894 14291 17950
rect 14359 17894 14415 17950
rect 14483 17894 14539 17950
rect 14607 17894 14663 17950
rect 12871 17770 12927 17826
rect 12995 17770 13051 17826
rect 13119 17770 13175 17826
rect 13243 17770 13299 17826
rect 13367 17770 13423 17826
rect 13491 17770 13547 17826
rect 13615 17770 13671 17826
rect 13739 17770 13795 17826
rect 13863 17770 13919 17826
rect 13987 17770 14043 17826
rect 14111 17770 14167 17826
rect 14235 17770 14291 17826
rect 14359 17770 14415 17826
rect 14483 17770 14539 17826
rect 14607 17770 14663 17826
rect 12871 17646 12927 17702
rect 12995 17646 13051 17702
rect 13119 17646 13175 17702
rect 13243 17646 13299 17702
rect 13367 17646 13423 17702
rect 13491 17646 13547 17702
rect 13615 17646 13671 17702
rect 13739 17646 13795 17702
rect 13863 17646 13919 17702
rect 13987 17646 14043 17702
rect 14111 17646 14167 17702
rect 14235 17646 14291 17702
rect 14359 17646 14415 17702
rect 14483 17646 14539 17702
rect 14607 17646 14663 17702
rect 315 17298 371 17354
rect 439 17298 495 17354
rect 563 17298 619 17354
rect 687 17298 743 17354
rect 811 17298 867 17354
rect 935 17298 991 17354
rect 1059 17298 1115 17354
rect 1183 17298 1239 17354
rect 1307 17298 1363 17354
rect 1431 17298 1487 17354
rect 1555 17298 1611 17354
rect 1679 17298 1735 17354
rect 1803 17298 1859 17354
rect 1927 17298 1983 17354
rect 2051 17298 2107 17354
rect 315 17174 371 17230
rect 439 17174 495 17230
rect 563 17174 619 17230
rect 687 17174 743 17230
rect 811 17174 867 17230
rect 935 17174 991 17230
rect 1059 17174 1115 17230
rect 1183 17174 1239 17230
rect 1307 17174 1363 17230
rect 1431 17174 1487 17230
rect 1555 17174 1611 17230
rect 1679 17174 1735 17230
rect 1803 17174 1859 17230
rect 1927 17174 1983 17230
rect 2051 17174 2107 17230
rect 315 17050 371 17106
rect 439 17050 495 17106
rect 563 17050 619 17106
rect 687 17050 743 17106
rect 811 17050 867 17106
rect 935 17050 991 17106
rect 1059 17050 1115 17106
rect 1183 17050 1239 17106
rect 1307 17050 1363 17106
rect 1431 17050 1487 17106
rect 1555 17050 1611 17106
rect 1679 17050 1735 17106
rect 1803 17050 1859 17106
rect 1927 17050 1983 17106
rect 2051 17050 2107 17106
rect 315 16926 371 16982
rect 439 16926 495 16982
rect 563 16926 619 16982
rect 687 16926 743 16982
rect 811 16926 867 16982
rect 935 16926 991 16982
rect 1059 16926 1115 16982
rect 1183 16926 1239 16982
rect 1307 16926 1363 16982
rect 1431 16926 1487 16982
rect 1555 16926 1611 16982
rect 1679 16926 1735 16982
rect 1803 16926 1859 16982
rect 1927 16926 1983 16982
rect 2051 16926 2107 16982
rect 315 16802 371 16858
rect 439 16802 495 16858
rect 563 16802 619 16858
rect 687 16802 743 16858
rect 811 16802 867 16858
rect 935 16802 991 16858
rect 1059 16802 1115 16858
rect 1183 16802 1239 16858
rect 1307 16802 1363 16858
rect 1431 16802 1487 16858
rect 1555 16802 1611 16858
rect 1679 16802 1735 16858
rect 1803 16802 1859 16858
rect 1927 16802 1983 16858
rect 2051 16802 2107 16858
rect 315 16678 371 16734
rect 439 16678 495 16734
rect 563 16678 619 16734
rect 687 16678 743 16734
rect 811 16678 867 16734
rect 935 16678 991 16734
rect 1059 16678 1115 16734
rect 1183 16678 1239 16734
rect 1307 16678 1363 16734
rect 1431 16678 1487 16734
rect 1555 16678 1611 16734
rect 1679 16678 1735 16734
rect 1803 16678 1859 16734
rect 1927 16678 1983 16734
rect 2051 16678 2107 16734
rect 315 16554 371 16610
rect 439 16554 495 16610
rect 563 16554 619 16610
rect 687 16554 743 16610
rect 811 16554 867 16610
rect 935 16554 991 16610
rect 1059 16554 1115 16610
rect 1183 16554 1239 16610
rect 1307 16554 1363 16610
rect 1431 16554 1487 16610
rect 1555 16554 1611 16610
rect 1679 16554 1735 16610
rect 1803 16554 1859 16610
rect 1927 16554 1983 16610
rect 2051 16554 2107 16610
rect 315 16430 371 16486
rect 439 16430 495 16486
rect 563 16430 619 16486
rect 687 16430 743 16486
rect 811 16430 867 16486
rect 935 16430 991 16486
rect 1059 16430 1115 16486
rect 1183 16430 1239 16486
rect 1307 16430 1363 16486
rect 1431 16430 1487 16486
rect 1555 16430 1611 16486
rect 1679 16430 1735 16486
rect 1803 16430 1859 16486
rect 1927 16430 1983 16486
rect 2051 16430 2107 16486
rect 315 16306 371 16362
rect 439 16306 495 16362
rect 563 16306 619 16362
rect 687 16306 743 16362
rect 811 16306 867 16362
rect 935 16306 991 16362
rect 1059 16306 1115 16362
rect 1183 16306 1239 16362
rect 1307 16306 1363 16362
rect 1431 16306 1487 16362
rect 1555 16306 1611 16362
rect 1679 16306 1735 16362
rect 1803 16306 1859 16362
rect 1927 16306 1983 16362
rect 2051 16306 2107 16362
rect 315 16182 371 16238
rect 439 16182 495 16238
rect 563 16182 619 16238
rect 687 16182 743 16238
rect 811 16182 867 16238
rect 935 16182 991 16238
rect 1059 16182 1115 16238
rect 1183 16182 1239 16238
rect 1307 16182 1363 16238
rect 1431 16182 1487 16238
rect 1555 16182 1611 16238
rect 1679 16182 1735 16238
rect 1803 16182 1859 16238
rect 1927 16182 1983 16238
rect 2051 16182 2107 16238
rect 315 16058 371 16114
rect 439 16058 495 16114
rect 563 16058 619 16114
rect 687 16058 743 16114
rect 811 16058 867 16114
rect 935 16058 991 16114
rect 1059 16058 1115 16114
rect 1183 16058 1239 16114
rect 1307 16058 1363 16114
rect 1431 16058 1487 16114
rect 1555 16058 1611 16114
rect 1679 16058 1735 16114
rect 1803 16058 1859 16114
rect 1927 16058 1983 16114
rect 2051 16058 2107 16114
rect 315 15934 371 15990
rect 439 15934 495 15990
rect 563 15934 619 15990
rect 687 15934 743 15990
rect 811 15934 867 15990
rect 935 15934 991 15990
rect 1059 15934 1115 15990
rect 1183 15934 1239 15990
rect 1307 15934 1363 15990
rect 1431 15934 1487 15990
rect 1555 15934 1611 15990
rect 1679 15934 1735 15990
rect 1803 15934 1859 15990
rect 1927 15934 1983 15990
rect 2051 15934 2107 15990
rect 315 15810 371 15866
rect 439 15810 495 15866
rect 563 15810 619 15866
rect 687 15810 743 15866
rect 811 15810 867 15866
rect 935 15810 991 15866
rect 1059 15810 1115 15866
rect 1183 15810 1239 15866
rect 1307 15810 1363 15866
rect 1431 15810 1487 15866
rect 1555 15810 1611 15866
rect 1679 15810 1735 15866
rect 1803 15810 1859 15866
rect 1927 15810 1983 15866
rect 2051 15810 2107 15866
rect 315 15686 371 15742
rect 439 15686 495 15742
rect 563 15686 619 15742
rect 687 15686 743 15742
rect 811 15686 867 15742
rect 935 15686 991 15742
rect 1059 15686 1115 15742
rect 1183 15686 1239 15742
rect 1307 15686 1363 15742
rect 1431 15686 1487 15742
rect 1555 15686 1611 15742
rect 1679 15686 1735 15742
rect 1803 15686 1859 15742
rect 1927 15686 1983 15742
rect 2051 15686 2107 15742
rect 315 15562 371 15618
rect 439 15562 495 15618
rect 563 15562 619 15618
rect 687 15562 743 15618
rect 811 15562 867 15618
rect 935 15562 991 15618
rect 1059 15562 1115 15618
rect 1183 15562 1239 15618
rect 1307 15562 1363 15618
rect 1431 15562 1487 15618
rect 1555 15562 1611 15618
rect 1679 15562 1735 15618
rect 1803 15562 1859 15618
rect 1927 15562 1983 15618
rect 2051 15562 2107 15618
rect 315 15438 371 15494
rect 439 15438 495 15494
rect 563 15438 619 15494
rect 687 15438 743 15494
rect 811 15438 867 15494
rect 935 15438 991 15494
rect 1059 15438 1115 15494
rect 1183 15438 1239 15494
rect 1307 15438 1363 15494
rect 1431 15438 1487 15494
rect 1555 15438 1611 15494
rect 1679 15438 1735 15494
rect 1803 15438 1859 15494
rect 1927 15438 1983 15494
rect 2051 15438 2107 15494
rect 315 15314 371 15370
rect 439 15314 495 15370
rect 563 15314 619 15370
rect 687 15314 743 15370
rect 811 15314 867 15370
rect 935 15314 991 15370
rect 1059 15314 1115 15370
rect 1183 15314 1239 15370
rect 1307 15314 1363 15370
rect 1431 15314 1487 15370
rect 1555 15314 1611 15370
rect 1679 15314 1735 15370
rect 1803 15314 1859 15370
rect 1927 15314 1983 15370
rect 2051 15314 2107 15370
rect 315 15190 371 15246
rect 439 15190 495 15246
rect 563 15190 619 15246
rect 687 15190 743 15246
rect 811 15190 867 15246
rect 935 15190 991 15246
rect 1059 15190 1115 15246
rect 1183 15190 1239 15246
rect 1307 15190 1363 15246
rect 1431 15190 1487 15246
rect 1555 15190 1611 15246
rect 1679 15190 1735 15246
rect 1803 15190 1859 15246
rect 1927 15190 1983 15246
rect 2051 15190 2107 15246
rect 315 15066 371 15122
rect 439 15066 495 15122
rect 563 15066 619 15122
rect 687 15066 743 15122
rect 811 15066 867 15122
rect 935 15066 991 15122
rect 1059 15066 1115 15122
rect 1183 15066 1239 15122
rect 1307 15066 1363 15122
rect 1431 15066 1487 15122
rect 1555 15066 1611 15122
rect 1679 15066 1735 15122
rect 1803 15066 1859 15122
rect 1927 15066 1983 15122
rect 2051 15066 2107 15122
rect 315 14942 371 14998
rect 439 14942 495 14998
rect 563 14942 619 14998
rect 687 14942 743 14998
rect 811 14942 867 14998
rect 935 14942 991 14998
rect 1059 14942 1115 14998
rect 1183 14942 1239 14998
rect 1307 14942 1363 14998
rect 1431 14942 1487 14998
rect 1555 14942 1611 14998
rect 1679 14942 1735 14998
rect 1803 14942 1859 14998
rect 1927 14942 1983 14998
rect 2051 14942 2107 14998
rect 315 14818 371 14874
rect 439 14818 495 14874
rect 563 14818 619 14874
rect 687 14818 743 14874
rect 811 14818 867 14874
rect 935 14818 991 14874
rect 1059 14818 1115 14874
rect 1183 14818 1239 14874
rect 1307 14818 1363 14874
rect 1431 14818 1487 14874
rect 1555 14818 1611 14874
rect 1679 14818 1735 14874
rect 1803 14818 1859 14874
rect 1927 14818 1983 14874
rect 2051 14818 2107 14874
rect 315 14694 371 14750
rect 439 14694 495 14750
rect 563 14694 619 14750
rect 687 14694 743 14750
rect 811 14694 867 14750
rect 935 14694 991 14750
rect 1059 14694 1115 14750
rect 1183 14694 1239 14750
rect 1307 14694 1363 14750
rect 1431 14694 1487 14750
rect 1555 14694 1611 14750
rect 1679 14694 1735 14750
rect 1803 14694 1859 14750
rect 1927 14694 1983 14750
rect 2051 14694 2107 14750
rect 315 14570 371 14626
rect 439 14570 495 14626
rect 563 14570 619 14626
rect 687 14570 743 14626
rect 811 14570 867 14626
rect 935 14570 991 14626
rect 1059 14570 1115 14626
rect 1183 14570 1239 14626
rect 1307 14570 1363 14626
rect 1431 14570 1487 14626
rect 1555 14570 1611 14626
rect 1679 14570 1735 14626
rect 1803 14570 1859 14626
rect 1927 14570 1983 14626
rect 2051 14570 2107 14626
rect 315 14446 371 14502
rect 439 14446 495 14502
rect 563 14446 619 14502
rect 687 14446 743 14502
rect 811 14446 867 14502
rect 935 14446 991 14502
rect 1059 14446 1115 14502
rect 1183 14446 1239 14502
rect 1307 14446 1363 14502
rect 1431 14446 1487 14502
rect 1555 14446 1611 14502
rect 1679 14446 1735 14502
rect 1803 14446 1859 14502
rect 1927 14446 1983 14502
rect 2051 14446 2107 14502
rect 2808 17298 2864 17354
rect 2932 17298 2988 17354
rect 3056 17298 3112 17354
rect 3180 17298 3236 17354
rect 3304 17298 3360 17354
rect 3428 17298 3484 17354
rect 3552 17298 3608 17354
rect 3676 17298 3732 17354
rect 3800 17298 3856 17354
rect 3924 17298 3980 17354
rect 4048 17298 4104 17354
rect 4172 17298 4228 17354
rect 4296 17298 4352 17354
rect 4420 17298 4476 17354
rect 4544 17298 4600 17354
rect 4668 17298 4724 17354
rect 2808 17174 2864 17230
rect 2932 17174 2988 17230
rect 3056 17174 3112 17230
rect 3180 17174 3236 17230
rect 3304 17174 3360 17230
rect 3428 17174 3484 17230
rect 3552 17174 3608 17230
rect 3676 17174 3732 17230
rect 3800 17174 3856 17230
rect 3924 17174 3980 17230
rect 4048 17174 4104 17230
rect 4172 17174 4228 17230
rect 4296 17174 4352 17230
rect 4420 17174 4476 17230
rect 4544 17174 4600 17230
rect 4668 17174 4724 17230
rect 2808 17050 2864 17106
rect 2932 17050 2988 17106
rect 3056 17050 3112 17106
rect 3180 17050 3236 17106
rect 3304 17050 3360 17106
rect 3428 17050 3484 17106
rect 3552 17050 3608 17106
rect 3676 17050 3732 17106
rect 3800 17050 3856 17106
rect 3924 17050 3980 17106
rect 4048 17050 4104 17106
rect 4172 17050 4228 17106
rect 4296 17050 4352 17106
rect 4420 17050 4476 17106
rect 4544 17050 4600 17106
rect 4668 17050 4724 17106
rect 2808 16926 2864 16982
rect 2932 16926 2988 16982
rect 3056 16926 3112 16982
rect 3180 16926 3236 16982
rect 3304 16926 3360 16982
rect 3428 16926 3484 16982
rect 3552 16926 3608 16982
rect 3676 16926 3732 16982
rect 3800 16926 3856 16982
rect 3924 16926 3980 16982
rect 4048 16926 4104 16982
rect 4172 16926 4228 16982
rect 4296 16926 4352 16982
rect 4420 16926 4476 16982
rect 4544 16926 4600 16982
rect 4668 16926 4724 16982
rect 2808 16802 2864 16858
rect 2932 16802 2988 16858
rect 3056 16802 3112 16858
rect 3180 16802 3236 16858
rect 3304 16802 3360 16858
rect 3428 16802 3484 16858
rect 3552 16802 3608 16858
rect 3676 16802 3732 16858
rect 3800 16802 3856 16858
rect 3924 16802 3980 16858
rect 4048 16802 4104 16858
rect 4172 16802 4228 16858
rect 4296 16802 4352 16858
rect 4420 16802 4476 16858
rect 4544 16802 4600 16858
rect 4668 16802 4724 16858
rect 2808 16678 2864 16734
rect 2932 16678 2988 16734
rect 3056 16678 3112 16734
rect 3180 16678 3236 16734
rect 3304 16678 3360 16734
rect 3428 16678 3484 16734
rect 3552 16678 3608 16734
rect 3676 16678 3732 16734
rect 3800 16678 3856 16734
rect 3924 16678 3980 16734
rect 4048 16678 4104 16734
rect 4172 16678 4228 16734
rect 4296 16678 4352 16734
rect 4420 16678 4476 16734
rect 4544 16678 4600 16734
rect 4668 16678 4724 16734
rect 2808 16554 2864 16610
rect 2932 16554 2988 16610
rect 3056 16554 3112 16610
rect 3180 16554 3236 16610
rect 3304 16554 3360 16610
rect 3428 16554 3484 16610
rect 3552 16554 3608 16610
rect 3676 16554 3732 16610
rect 3800 16554 3856 16610
rect 3924 16554 3980 16610
rect 4048 16554 4104 16610
rect 4172 16554 4228 16610
rect 4296 16554 4352 16610
rect 4420 16554 4476 16610
rect 4544 16554 4600 16610
rect 4668 16554 4724 16610
rect 2808 16430 2864 16486
rect 2932 16430 2988 16486
rect 3056 16430 3112 16486
rect 3180 16430 3236 16486
rect 3304 16430 3360 16486
rect 3428 16430 3484 16486
rect 3552 16430 3608 16486
rect 3676 16430 3732 16486
rect 3800 16430 3856 16486
rect 3924 16430 3980 16486
rect 4048 16430 4104 16486
rect 4172 16430 4228 16486
rect 4296 16430 4352 16486
rect 4420 16430 4476 16486
rect 4544 16430 4600 16486
rect 4668 16430 4724 16486
rect 2808 16306 2864 16362
rect 2932 16306 2988 16362
rect 3056 16306 3112 16362
rect 3180 16306 3236 16362
rect 3304 16306 3360 16362
rect 3428 16306 3484 16362
rect 3552 16306 3608 16362
rect 3676 16306 3732 16362
rect 3800 16306 3856 16362
rect 3924 16306 3980 16362
rect 4048 16306 4104 16362
rect 4172 16306 4228 16362
rect 4296 16306 4352 16362
rect 4420 16306 4476 16362
rect 4544 16306 4600 16362
rect 4668 16306 4724 16362
rect 2808 16182 2864 16238
rect 2932 16182 2988 16238
rect 3056 16182 3112 16238
rect 3180 16182 3236 16238
rect 3304 16182 3360 16238
rect 3428 16182 3484 16238
rect 3552 16182 3608 16238
rect 3676 16182 3732 16238
rect 3800 16182 3856 16238
rect 3924 16182 3980 16238
rect 4048 16182 4104 16238
rect 4172 16182 4228 16238
rect 4296 16182 4352 16238
rect 4420 16182 4476 16238
rect 4544 16182 4600 16238
rect 4668 16182 4724 16238
rect 2808 16058 2864 16114
rect 2932 16058 2988 16114
rect 3056 16058 3112 16114
rect 3180 16058 3236 16114
rect 3304 16058 3360 16114
rect 3428 16058 3484 16114
rect 3552 16058 3608 16114
rect 3676 16058 3732 16114
rect 3800 16058 3856 16114
rect 3924 16058 3980 16114
rect 4048 16058 4104 16114
rect 4172 16058 4228 16114
rect 4296 16058 4352 16114
rect 4420 16058 4476 16114
rect 4544 16058 4600 16114
rect 4668 16058 4724 16114
rect 2808 15934 2864 15990
rect 2932 15934 2988 15990
rect 3056 15934 3112 15990
rect 3180 15934 3236 15990
rect 3304 15934 3360 15990
rect 3428 15934 3484 15990
rect 3552 15934 3608 15990
rect 3676 15934 3732 15990
rect 3800 15934 3856 15990
rect 3924 15934 3980 15990
rect 4048 15934 4104 15990
rect 4172 15934 4228 15990
rect 4296 15934 4352 15990
rect 4420 15934 4476 15990
rect 4544 15934 4600 15990
rect 4668 15934 4724 15990
rect 2808 15810 2864 15866
rect 2932 15810 2988 15866
rect 3056 15810 3112 15866
rect 3180 15810 3236 15866
rect 3304 15810 3360 15866
rect 3428 15810 3484 15866
rect 3552 15810 3608 15866
rect 3676 15810 3732 15866
rect 3800 15810 3856 15866
rect 3924 15810 3980 15866
rect 4048 15810 4104 15866
rect 4172 15810 4228 15866
rect 4296 15810 4352 15866
rect 4420 15810 4476 15866
rect 4544 15810 4600 15866
rect 4668 15810 4724 15866
rect 2808 15686 2864 15742
rect 2932 15686 2988 15742
rect 3056 15686 3112 15742
rect 3180 15686 3236 15742
rect 3304 15686 3360 15742
rect 3428 15686 3484 15742
rect 3552 15686 3608 15742
rect 3676 15686 3732 15742
rect 3800 15686 3856 15742
rect 3924 15686 3980 15742
rect 4048 15686 4104 15742
rect 4172 15686 4228 15742
rect 4296 15686 4352 15742
rect 4420 15686 4476 15742
rect 4544 15686 4600 15742
rect 4668 15686 4724 15742
rect 2808 15562 2864 15618
rect 2932 15562 2988 15618
rect 3056 15562 3112 15618
rect 3180 15562 3236 15618
rect 3304 15562 3360 15618
rect 3428 15562 3484 15618
rect 3552 15562 3608 15618
rect 3676 15562 3732 15618
rect 3800 15562 3856 15618
rect 3924 15562 3980 15618
rect 4048 15562 4104 15618
rect 4172 15562 4228 15618
rect 4296 15562 4352 15618
rect 4420 15562 4476 15618
rect 4544 15562 4600 15618
rect 4668 15562 4724 15618
rect 2808 15438 2864 15494
rect 2932 15438 2988 15494
rect 3056 15438 3112 15494
rect 3180 15438 3236 15494
rect 3304 15438 3360 15494
rect 3428 15438 3484 15494
rect 3552 15438 3608 15494
rect 3676 15438 3732 15494
rect 3800 15438 3856 15494
rect 3924 15438 3980 15494
rect 4048 15438 4104 15494
rect 4172 15438 4228 15494
rect 4296 15438 4352 15494
rect 4420 15438 4476 15494
rect 4544 15438 4600 15494
rect 4668 15438 4724 15494
rect 2808 15314 2864 15370
rect 2932 15314 2988 15370
rect 3056 15314 3112 15370
rect 3180 15314 3236 15370
rect 3304 15314 3360 15370
rect 3428 15314 3484 15370
rect 3552 15314 3608 15370
rect 3676 15314 3732 15370
rect 3800 15314 3856 15370
rect 3924 15314 3980 15370
rect 4048 15314 4104 15370
rect 4172 15314 4228 15370
rect 4296 15314 4352 15370
rect 4420 15314 4476 15370
rect 4544 15314 4600 15370
rect 4668 15314 4724 15370
rect 2808 15190 2864 15246
rect 2932 15190 2988 15246
rect 3056 15190 3112 15246
rect 3180 15190 3236 15246
rect 3304 15190 3360 15246
rect 3428 15190 3484 15246
rect 3552 15190 3608 15246
rect 3676 15190 3732 15246
rect 3800 15190 3856 15246
rect 3924 15190 3980 15246
rect 4048 15190 4104 15246
rect 4172 15190 4228 15246
rect 4296 15190 4352 15246
rect 4420 15190 4476 15246
rect 4544 15190 4600 15246
rect 4668 15190 4724 15246
rect 2808 15066 2864 15122
rect 2932 15066 2988 15122
rect 3056 15066 3112 15122
rect 3180 15066 3236 15122
rect 3304 15066 3360 15122
rect 3428 15066 3484 15122
rect 3552 15066 3608 15122
rect 3676 15066 3732 15122
rect 3800 15066 3856 15122
rect 3924 15066 3980 15122
rect 4048 15066 4104 15122
rect 4172 15066 4228 15122
rect 4296 15066 4352 15122
rect 4420 15066 4476 15122
rect 4544 15066 4600 15122
rect 4668 15066 4724 15122
rect 2808 14942 2864 14998
rect 2932 14942 2988 14998
rect 3056 14942 3112 14998
rect 3180 14942 3236 14998
rect 3304 14942 3360 14998
rect 3428 14942 3484 14998
rect 3552 14942 3608 14998
rect 3676 14942 3732 14998
rect 3800 14942 3856 14998
rect 3924 14942 3980 14998
rect 4048 14942 4104 14998
rect 4172 14942 4228 14998
rect 4296 14942 4352 14998
rect 4420 14942 4476 14998
rect 4544 14942 4600 14998
rect 4668 14942 4724 14998
rect 2808 14818 2864 14874
rect 2932 14818 2988 14874
rect 3056 14818 3112 14874
rect 3180 14818 3236 14874
rect 3304 14818 3360 14874
rect 3428 14818 3484 14874
rect 3552 14818 3608 14874
rect 3676 14818 3732 14874
rect 3800 14818 3856 14874
rect 3924 14818 3980 14874
rect 4048 14818 4104 14874
rect 4172 14818 4228 14874
rect 4296 14818 4352 14874
rect 4420 14818 4476 14874
rect 4544 14818 4600 14874
rect 4668 14818 4724 14874
rect 2808 14694 2864 14750
rect 2932 14694 2988 14750
rect 3056 14694 3112 14750
rect 3180 14694 3236 14750
rect 3304 14694 3360 14750
rect 3428 14694 3484 14750
rect 3552 14694 3608 14750
rect 3676 14694 3732 14750
rect 3800 14694 3856 14750
rect 3924 14694 3980 14750
rect 4048 14694 4104 14750
rect 4172 14694 4228 14750
rect 4296 14694 4352 14750
rect 4420 14694 4476 14750
rect 4544 14694 4600 14750
rect 4668 14694 4724 14750
rect 2808 14570 2864 14626
rect 2932 14570 2988 14626
rect 3056 14570 3112 14626
rect 3180 14570 3236 14626
rect 3304 14570 3360 14626
rect 3428 14570 3484 14626
rect 3552 14570 3608 14626
rect 3676 14570 3732 14626
rect 3800 14570 3856 14626
rect 3924 14570 3980 14626
rect 4048 14570 4104 14626
rect 4172 14570 4228 14626
rect 4296 14570 4352 14626
rect 4420 14570 4476 14626
rect 4544 14570 4600 14626
rect 4668 14570 4724 14626
rect 2808 14446 2864 14502
rect 2932 14446 2988 14502
rect 3056 14446 3112 14502
rect 3180 14446 3236 14502
rect 3304 14446 3360 14502
rect 3428 14446 3484 14502
rect 3552 14446 3608 14502
rect 3676 14446 3732 14502
rect 3800 14446 3856 14502
rect 3924 14446 3980 14502
rect 4048 14446 4104 14502
rect 4172 14446 4228 14502
rect 4296 14446 4352 14502
rect 4420 14446 4476 14502
rect 4544 14446 4600 14502
rect 4668 14446 4724 14502
rect 5178 17298 5234 17354
rect 5302 17298 5358 17354
rect 5426 17298 5482 17354
rect 5550 17298 5606 17354
rect 5674 17298 5730 17354
rect 5798 17298 5854 17354
rect 5922 17298 5978 17354
rect 6046 17298 6102 17354
rect 6170 17298 6226 17354
rect 6294 17298 6350 17354
rect 6418 17298 6474 17354
rect 6542 17298 6598 17354
rect 6666 17298 6722 17354
rect 6790 17298 6846 17354
rect 6914 17298 6970 17354
rect 7038 17298 7094 17354
rect 5178 17174 5234 17230
rect 5302 17174 5358 17230
rect 5426 17174 5482 17230
rect 5550 17174 5606 17230
rect 5674 17174 5730 17230
rect 5798 17174 5854 17230
rect 5922 17174 5978 17230
rect 6046 17174 6102 17230
rect 6170 17174 6226 17230
rect 6294 17174 6350 17230
rect 6418 17174 6474 17230
rect 6542 17174 6598 17230
rect 6666 17174 6722 17230
rect 6790 17174 6846 17230
rect 6914 17174 6970 17230
rect 7038 17174 7094 17230
rect 5178 17050 5234 17106
rect 5302 17050 5358 17106
rect 5426 17050 5482 17106
rect 5550 17050 5606 17106
rect 5674 17050 5730 17106
rect 5798 17050 5854 17106
rect 5922 17050 5978 17106
rect 6046 17050 6102 17106
rect 6170 17050 6226 17106
rect 6294 17050 6350 17106
rect 6418 17050 6474 17106
rect 6542 17050 6598 17106
rect 6666 17050 6722 17106
rect 6790 17050 6846 17106
rect 6914 17050 6970 17106
rect 7038 17050 7094 17106
rect 5178 16926 5234 16982
rect 5302 16926 5358 16982
rect 5426 16926 5482 16982
rect 5550 16926 5606 16982
rect 5674 16926 5730 16982
rect 5798 16926 5854 16982
rect 5922 16926 5978 16982
rect 6046 16926 6102 16982
rect 6170 16926 6226 16982
rect 6294 16926 6350 16982
rect 6418 16926 6474 16982
rect 6542 16926 6598 16982
rect 6666 16926 6722 16982
rect 6790 16926 6846 16982
rect 6914 16926 6970 16982
rect 7038 16926 7094 16982
rect 5178 16802 5234 16858
rect 5302 16802 5358 16858
rect 5426 16802 5482 16858
rect 5550 16802 5606 16858
rect 5674 16802 5730 16858
rect 5798 16802 5854 16858
rect 5922 16802 5978 16858
rect 6046 16802 6102 16858
rect 6170 16802 6226 16858
rect 6294 16802 6350 16858
rect 6418 16802 6474 16858
rect 6542 16802 6598 16858
rect 6666 16802 6722 16858
rect 6790 16802 6846 16858
rect 6914 16802 6970 16858
rect 7038 16802 7094 16858
rect 5178 16678 5234 16734
rect 5302 16678 5358 16734
rect 5426 16678 5482 16734
rect 5550 16678 5606 16734
rect 5674 16678 5730 16734
rect 5798 16678 5854 16734
rect 5922 16678 5978 16734
rect 6046 16678 6102 16734
rect 6170 16678 6226 16734
rect 6294 16678 6350 16734
rect 6418 16678 6474 16734
rect 6542 16678 6598 16734
rect 6666 16678 6722 16734
rect 6790 16678 6846 16734
rect 6914 16678 6970 16734
rect 7038 16678 7094 16734
rect 5178 16554 5234 16610
rect 5302 16554 5358 16610
rect 5426 16554 5482 16610
rect 5550 16554 5606 16610
rect 5674 16554 5730 16610
rect 5798 16554 5854 16610
rect 5922 16554 5978 16610
rect 6046 16554 6102 16610
rect 6170 16554 6226 16610
rect 6294 16554 6350 16610
rect 6418 16554 6474 16610
rect 6542 16554 6598 16610
rect 6666 16554 6722 16610
rect 6790 16554 6846 16610
rect 6914 16554 6970 16610
rect 7038 16554 7094 16610
rect 5178 16430 5234 16486
rect 5302 16430 5358 16486
rect 5426 16430 5482 16486
rect 5550 16430 5606 16486
rect 5674 16430 5730 16486
rect 5798 16430 5854 16486
rect 5922 16430 5978 16486
rect 6046 16430 6102 16486
rect 6170 16430 6226 16486
rect 6294 16430 6350 16486
rect 6418 16430 6474 16486
rect 6542 16430 6598 16486
rect 6666 16430 6722 16486
rect 6790 16430 6846 16486
rect 6914 16430 6970 16486
rect 7038 16430 7094 16486
rect 5178 16306 5234 16362
rect 5302 16306 5358 16362
rect 5426 16306 5482 16362
rect 5550 16306 5606 16362
rect 5674 16306 5730 16362
rect 5798 16306 5854 16362
rect 5922 16306 5978 16362
rect 6046 16306 6102 16362
rect 6170 16306 6226 16362
rect 6294 16306 6350 16362
rect 6418 16306 6474 16362
rect 6542 16306 6598 16362
rect 6666 16306 6722 16362
rect 6790 16306 6846 16362
rect 6914 16306 6970 16362
rect 7038 16306 7094 16362
rect 5178 16182 5234 16238
rect 5302 16182 5358 16238
rect 5426 16182 5482 16238
rect 5550 16182 5606 16238
rect 5674 16182 5730 16238
rect 5798 16182 5854 16238
rect 5922 16182 5978 16238
rect 6046 16182 6102 16238
rect 6170 16182 6226 16238
rect 6294 16182 6350 16238
rect 6418 16182 6474 16238
rect 6542 16182 6598 16238
rect 6666 16182 6722 16238
rect 6790 16182 6846 16238
rect 6914 16182 6970 16238
rect 7038 16182 7094 16238
rect 5178 16058 5234 16114
rect 5302 16058 5358 16114
rect 5426 16058 5482 16114
rect 5550 16058 5606 16114
rect 5674 16058 5730 16114
rect 5798 16058 5854 16114
rect 5922 16058 5978 16114
rect 6046 16058 6102 16114
rect 6170 16058 6226 16114
rect 6294 16058 6350 16114
rect 6418 16058 6474 16114
rect 6542 16058 6598 16114
rect 6666 16058 6722 16114
rect 6790 16058 6846 16114
rect 6914 16058 6970 16114
rect 7038 16058 7094 16114
rect 5178 15934 5234 15990
rect 5302 15934 5358 15990
rect 5426 15934 5482 15990
rect 5550 15934 5606 15990
rect 5674 15934 5730 15990
rect 5798 15934 5854 15990
rect 5922 15934 5978 15990
rect 6046 15934 6102 15990
rect 6170 15934 6226 15990
rect 6294 15934 6350 15990
rect 6418 15934 6474 15990
rect 6542 15934 6598 15990
rect 6666 15934 6722 15990
rect 6790 15934 6846 15990
rect 6914 15934 6970 15990
rect 7038 15934 7094 15990
rect 5178 15810 5234 15866
rect 5302 15810 5358 15866
rect 5426 15810 5482 15866
rect 5550 15810 5606 15866
rect 5674 15810 5730 15866
rect 5798 15810 5854 15866
rect 5922 15810 5978 15866
rect 6046 15810 6102 15866
rect 6170 15810 6226 15866
rect 6294 15810 6350 15866
rect 6418 15810 6474 15866
rect 6542 15810 6598 15866
rect 6666 15810 6722 15866
rect 6790 15810 6846 15866
rect 6914 15810 6970 15866
rect 7038 15810 7094 15866
rect 5178 15686 5234 15742
rect 5302 15686 5358 15742
rect 5426 15686 5482 15742
rect 5550 15686 5606 15742
rect 5674 15686 5730 15742
rect 5798 15686 5854 15742
rect 5922 15686 5978 15742
rect 6046 15686 6102 15742
rect 6170 15686 6226 15742
rect 6294 15686 6350 15742
rect 6418 15686 6474 15742
rect 6542 15686 6598 15742
rect 6666 15686 6722 15742
rect 6790 15686 6846 15742
rect 6914 15686 6970 15742
rect 7038 15686 7094 15742
rect 5178 15562 5234 15618
rect 5302 15562 5358 15618
rect 5426 15562 5482 15618
rect 5550 15562 5606 15618
rect 5674 15562 5730 15618
rect 5798 15562 5854 15618
rect 5922 15562 5978 15618
rect 6046 15562 6102 15618
rect 6170 15562 6226 15618
rect 6294 15562 6350 15618
rect 6418 15562 6474 15618
rect 6542 15562 6598 15618
rect 6666 15562 6722 15618
rect 6790 15562 6846 15618
rect 6914 15562 6970 15618
rect 7038 15562 7094 15618
rect 5178 15438 5234 15494
rect 5302 15438 5358 15494
rect 5426 15438 5482 15494
rect 5550 15438 5606 15494
rect 5674 15438 5730 15494
rect 5798 15438 5854 15494
rect 5922 15438 5978 15494
rect 6046 15438 6102 15494
rect 6170 15438 6226 15494
rect 6294 15438 6350 15494
rect 6418 15438 6474 15494
rect 6542 15438 6598 15494
rect 6666 15438 6722 15494
rect 6790 15438 6846 15494
rect 6914 15438 6970 15494
rect 7038 15438 7094 15494
rect 5178 15314 5234 15370
rect 5302 15314 5358 15370
rect 5426 15314 5482 15370
rect 5550 15314 5606 15370
rect 5674 15314 5730 15370
rect 5798 15314 5854 15370
rect 5922 15314 5978 15370
rect 6046 15314 6102 15370
rect 6170 15314 6226 15370
rect 6294 15314 6350 15370
rect 6418 15314 6474 15370
rect 6542 15314 6598 15370
rect 6666 15314 6722 15370
rect 6790 15314 6846 15370
rect 6914 15314 6970 15370
rect 7038 15314 7094 15370
rect 5178 15190 5234 15246
rect 5302 15190 5358 15246
rect 5426 15190 5482 15246
rect 5550 15190 5606 15246
rect 5674 15190 5730 15246
rect 5798 15190 5854 15246
rect 5922 15190 5978 15246
rect 6046 15190 6102 15246
rect 6170 15190 6226 15246
rect 6294 15190 6350 15246
rect 6418 15190 6474 15246
rect 6542 15190 6598 15246
rect 6666 15190 6722 15246
rect 6790 15190 6846 15246
rect 6914 15190 6970 15246
rect 7038 15190 7094 15246
rect 5178 15066 5234 15122
rect 5302 15066 5358 15122
rect 5426 15066 5482 15122
rect 5550 15066 5606 15122
rect 5674 15066 5730 15122
rect 5798 15066 5854 15122
rect 5922 15066 5978 15122
rect 6046 15066 6102 15122
rect 6170 15066 6226 15122
rect 6294 15066 6350 15122
rect 6418 15066 6474 15122
rect 6542 15066 6598 15122
rect 6666 15066 6722 15122
rect 6790 15066 6846 15122
rect 6914 15066 6970 15122
rect 7038 15066 7094 15122
rect 5178 14942 5234 14998
rect 5302 14942 5358 14998
rect 5426 14942 5482 14998
rect 5550 14942 5606 14998
rect 5674 14942 5730 14998
rect 5798 14942 5854 14998
rect 5922 14942 5978 14998
rect 6046 14942 6102 14998
rect 6170 14942 6226 14998
rect 6294 14942 6350 14998
rect 6418 14942 6474 14998
rect 6542 14942 6598 14998
rect 6666 14942 6722 14998
rect 6790 14942 6846 14998
rect 6914 14942 6970 14998
rect 7038 14942 7094 14998
rect 5178 14818 5234 14874
rect 5302 14818 5358 14874
rect 5426 14818 5482 14874
rect 5550 14818 5606 14874
rect 5674 14818 5730 14874
rect 5798 14818 5854 14874
rect 5922 14818 5978 14874
rect 6046 14818 6102 14874
rect 6170 14818 6226 14874
rect 6294 14818 6350 14874
rect 6418 14818 6474 14874
rect 6542 14818 6598 14874
rect 6666 14818 6722 14874
rect 6790 14818 6846 14874
rect 6914 14818 6970 14874
rect 7038 14818 7094 14874
rect 5178 14694 5234 14750
rect 5302 14694 5358 14750
rect 5426 14694 5482 14750
rect 5550 14694 5606 14750
rect 5674 14694 5730 14750
rect 5798 14694 5854 14750
rect 5922 14694 5978 14750
rect 6046 14694 6102 14750
rect 6170 14694 6226 14750
rect 6294 14694 6350 14750
rect 6418 14694 6474 14750
rect 6542 14694 6598 14750
rect 6666 14694 6722 14750
rect 6790 14694 6846 14750
rect 6914 14694 6970 14750
rect 7038 14694 7094 14750
rect 5178 14570 5234 14626
rect 5302 14570 5358 14626
rect 5426 14570 5482 14626
rect 5550 14570 5606 14626
rect 5674 14570 5730 14626
rect 5798 14570 5854 14626
rect 5922 14570 5978 14626
rect 6046 14570 6102 14626
rect 6170 14570 6226 14626
rect 6294 14570 6350 14626
rect 6418 14570 6474 14626
rect 6542 14570 6598 14626
rect 6666 14570 6722 14626
rect 6790 14570 6846 14626
rect 6914 14570 6970 14626
rect 7038 14570 7094 14626
rect 5178 14446 5234 14502
rect 5302 14446 5358 14502
rect 5426 14446 5482 14502
rect 5550 14446 5606 14502
rect 5674 14446 5730 14502
rect 5798 14446 5854 14502
rect 5922 14446 5978 14502
rect 6046 14446 6102 14502
rect 6170 14446 6226 14502
rect 6294 14446 6350 14502
rect 6418 14446 6474 14502
rect 6542 14446 6598 14502
rect 6666 14446 6722 14502
rect 6790 14446 6846 14502
rect 6914 14446 6970 14502
rect 7038 14446 7094 14502
rect 7884 17298 7940 17354
rect 8008 17298 8064 17354
rect 8132 17298 8188 17354
rect 8256 17298 8312 17354
rect 8380 17298 8436 17354
rect 8504 17298 8560 17354
rect 8628 17298 8684 17354
rect 8752 17298 8808 17354
rect 8876 17298 8932 17354
rect 9000 17298 9056 17354
rect 9124 17298 9180 17354
rect 9248 17298 9304 17354
rect 9372 17298 9428 17354
rect 9496 17298 9552 17354
rect 9620 17298 9676 17354
rect 9744 17298 9800 17354
rect 7884 17174 7940 17230
rect 8008 17174 8064 17230
rect 8132 17174 8188 17230
rect 8256 17174 8312 17230
rect 8380 17174 8436 17230
rect 8504 17174 8560 17230
rect 8628 17174 8684 17230
rect 8752 17174 8808 17230
rect 8876 17174 8932 17230
rect 9000 17174 9056 17230
rect 9124 17174 9180 17230
rect 9248 17174 9304 17230
rect 9372 17174 9428 17230
rect 9496 17174 9552 17230
rect 9620 17174 9676 17230
rect 9744 17174 9800 17230
rect 7884 17050 7940 17106
rect 8008 17050 8064 17106
rect 8132 17050 8188 17106
rect 8256 17050 8312 17106
rect 8380 17050 8436 17106
rect 8504 17050 8560 17106
rect 8628 17050 8684 17106
rect 8752 17050 8808 17106
rect 8876 17050 8932 17106
rect 9000 17050 9056 17106
rect 9124 17050 9180 17106
rect 9248 17050 9304 17106
rect 9372 17050 9428 17106
rect 9496 17050 9552 17106
rect 9620 17050 9676 17106
rect 9744 17050 9800 17106
rect 7884 16926 7940 16982
rect 8008 16926 8064 16982
rect 8132 16926 8188 16982
rect 8256 16926 8312 16982
rect 8380 16926 8436 16982
rect 8504 16926 8560 16982
rect 8628 16926 8684 16982
rect 8752 16926 8808 16982
rect 8876 16926 8932 16982
rect 9000 16926 9056 16982
rect 9124 16926 9180 16982
rect 9248 16926 9304 16982
rect 9372 16926 9428 16982
rect 9496 16926 9552 16982
rect 9620 16926 9676 16982
rect 9744 16926 9800 16982
rect 7884 16802 7940 16858
rect 8008 16802 8064 16858
rect 8132 16802 8188 16858
rect 8256 16802 8312 16858
rect 8380 16802 8436 16858
rect 8504 16802 8560 16858
rect 8628 16802 8684 16858
rect 8752 16802 8808 16858
rect 8876 16802 8932 16858
rect 9000 16802 9056 16858
rect 9124 16802 9180 16858
rect 9248 16802 9304 16858
rect 9372 16802 9428 16858
rect 9496 16802 9552 16858
rect 9620 16802 9676 16858
rect 9744 16802 9800 16858
rect 7884 16678 7940 16734
rect 8008 16678 8064 16734
rect 8132 16678 8188 16734
rect 8256 16678 8312 16734
rect 8380 16678 8436 16734
rect 8504 16678 8560 16734
rect 8628 16678 8684 16734
rect 8752 16678 8808 16734
rect 8876 16678 8932 16734
rect 9000 16678 9056 16734
rect 9124 16678 9180 16734
rect 9248 16678 9304 16734
rect 9372 16678 9428 16734
rect 9496 16678 9552 16734
rect 9620 16678 9676 16734
rect 9744 16678 9800 16734
rect 7884 16554 7940 16610
rect 8008 16554 8064 16610
rect 8132 16554 8188 16610
rect 8256 16554 8312 16610
rect 8380 16554 8436 16610
rect 8504 16554 8560 16610
rect 8628 16554 8684 16610
rect 8752 16554 8808 16610
rect 8876 16554 8932 16610
rect 9000 16554 9056 16610
rect 9124 16554 9180 16610
rect 9248 16554 9304 16610
rect 9372 16554 9428 16610
rect 9496 16554 9552 16610
rect 9620 16554 9676 16610
rect 9744 16554 9800 16610
rect 7884 16430 7940 16486
rect 8008 16430 8064 16486
rect 8132 16430 8188 16486
rect 8256 16430 8312 16486
rect 8380 16430 8436 16486
rect 8504 16430 8560 16486
rect 8628 16430 8684 16486
rect 8752 16430 8808 16486
rect 8876 16430 8932 16486
rect 9000 16430 9056 16486
rect 9124 16430 9180 16486
rect 9248 16430 9304 16486
rect 9372 16430 9428 16486
rect 9496 16430 9552 16486
rect 9620 16430 9676 16486
rect 9744 16430 9800 16486
rect 7884 16306 7940 16362
rect 8008 16306 8064 16362
rect 8132 16306 8188 16362
rect 8256 16306 8312 16362
rect 8380 16306 8436 16362
rect 8504 16306 8560 16362
rect 8628 16306 8684 16362
rect 8752 16306 8808 16362
rect 8876 16306 8932 16362
rect 9000 16306 9056 16362
rect 9124 16306 9180 16362
rect 9248 16306 9304 16362
rect 9372 16306 9428 16362
rect 9496 16306 9552 16362
rect 9620 16306 9676 16362
rect 9744 16306 9800 16362
rect 7884 16182 7940 16238
rect 8008 16182 8064 16238
rect 8132 16182 8188 16238
rect 8256 16182 8312 16238
rect 8380 16182 8436 16238
rect 8504 16182 8560 16238
rect 8628 16182 8684 16238
rect 8752 16182 8808 16238
rect 8876 16182 8932 16238
rect 9000 16182 9056 16238
rect 9124 16182 9180 16238
rect 9248 16182 9304 16238
rect 9372 16182 9428 16238
rect 9496 16182 9552 16238
rect 9620 16182 9676 16238
rect 9744 16182 9800 16238
rect 7884 16058 7940 16114
rect 8008 16058 8064 16114
rect 8132 16058 8188 16114
rect 8256 16058 8312 16114
rect 8380 16058 8436 16114
rect 8504 16058 8560 16114
rect 8628 16058 8684 16114
rect 8752 16058 8808 16114
rect 8876 16058 8932 16114
rect 9000 16058 9056 16114
rect 9124 16058 9180 16114
rect 9248 16058 9304 16114
rect 9372 16058 9428 16114
rect 9496 16058 9552 16114
rect 9620 16058 9676 16114
rect 9744 16058 9800 16114
rect 7884 15934 7940 15990
rect 8008 15934 8064 15990
rect 8132 15934 8188 15990
rect 8256 15934 8312 15990
rect 8380 15934 8436 15990
rect 8504 15934 8560 15990
rect 8628 15934 8684 15990
rect 8752 15934 8808 15990
rect 8876 15934 8932 15990
rect 9000 15934 9056 15990
rect 9124 15934 9180 15990
rect 9248 15934 9304 15990
rect 9372 15934 9428 15990
rect 9496 15934 9552 15990
rect 9620 15934 9676 15990
rect 9744 15934 9800 15990
rect 7884 15810 7940 15866
rect 8008 15810 8064 15866
rect 8132 15810 8188 15866
rect 8256 15810 8312 15866
rect 8380 15810 8436 15866
rect 8504 15810 8560 15866
rect 8628 15810 8684 15866
rect 8752 15810 8808 15866
rect 8876 15810 8932 15866
rect 9000 15810 9056 15866
rect 9124 15810 9180 15866
rect 9248 15810 9304 15866
rect 9372 15810 9428 15866
rect 9496 15810 9552 15866
rect 9620 15810 9676 15866
rect 9744 15810 9800 15866
rect 7884 15686 7940 15742
rect 8008 15686 8064 15742
rect 8132 15686 8188 15742
rect 8256 15686 8312 15742
rect 8380 15686 8436 15742
rect 8504 15686 8560 15742
rect 8628 15686 8684 15742
rect 8752 15686 8808 15742
rect 8876 15686 8932 15742
rect 9000 15686 9056 15742
rect 9124 15686 9180 15742
rect 9248 15686 9304 15742
rect 9372 15686 9428 15742
rect 9496 15686 9552 15742
rect 9620 15686 9676 15742
rect 9744 15686 9800 15742
rect 7884 15562 7940 15618
rect 8008 15562 8064 15618
rect 8132 15562 8188 15618
rect 8256 15562 8312 15618
rect 8380 15562 8436 15618
rect 8504 15562 8560 15618
rect 8628 15562 8684 15618
rect 8752 15562 8808 15618
rect 8876 15562 8932 15618
rect 9000 15562 9056 15618
rect 9124 15562 9180 15618
rect 9248 15562 9304 15618
rect 9372 15562 9428 15618
rect 9496 15562 9552 15618
rect 9620 15562 9676 15618
rect 9744 15562 9800 15618
rect 7884 15438 7940 15494
rect 8008 15438 8064 15494
rect 8132 15438 8188 15494
rect 8256 15438 8312 15494
rect 8380 15438 8436 15494
rect 8504 15438 8560 15494
rect 8628 15438 8684 15494
rect 8752 15438 8808 15494
rect 8876 15438 8932 15494
rect 9000 15438 9056 15494
rect 9124 15438 9180 15494
rect 9248 15438 9304 15494
rect 9372 15438 9428 15494
rect 9496 15438 9552 15494
rect 9620 15438 9676 15494
rect 9744 15438 9800 15494
rect 7884 15314 7940 15370
rect 8008 15314 8064 15370
rect 8132 15314 8188 15370
rect 8256 15314 8312 15370
rect 8380 15314 8436 15370
rect 8504 15314 8560 15370
rect 8628 15314 8684 15370
rect 8752 15314 8808 15370
rect 8876 15314 8932 15370
rect 9000 15314 9056 15370
rect 9124 15314 9180 15370
rect 9248 15314 9304 15370
rect 9372 15314 9428 15370
rect 9496 15314 9552 15370
rect 9620 15314 9676 15370
rect 9744 15314 9800 15370
rect 7884 15190 7940 15246
rect 8008 15190 8064 15246
rect 8132 15190 8188 15246
rect 8256 15190 8312 15246
rect 8380 15190 8436 15246
rect 8504 15190 8560 15246
rect 8628 15190 8684 15246
rect 8752 15190 8808 15246
rect 8876 15190 8932 15246
rect 9000 15190 9056 15246
rect 9124 15190 9180 15246
rect 9248 15190 9304 15246
rect 9372 15190 9428 15246
rect 9496 15190 9552 15246
rect 9620 15190 9676 15246
rect 9744 15190 9800 15246
rect 7884 15066 7940 15122
rect 8008 15066 8064 15122
rect 8132 15066 8188 15122
rect 8256 15066 8312 15122
rect 8380 15066 8436 15122
rect 8504 15066 8560 15122
rect 8628 15066 8684 15122
rect 8752 15066 8808 15122
rect 8876 15066 8932 15122
rect 9000 15066 9056 15122
rect 9124 15066 9180 15122
rect 9248 15066 9304 15122
rect 9372 15066 9428 15122
rect 9496 15066 9552 15122
rect 9620 15066 9676 15122
rect 9744 15066 9800 15122
rect 7884 14942 7940 14998
rect 8008 14942 8064 14998
rect 8132 14942 8188 14998
rect 8256 14942 8312 14998
rect 8380 14942 8436 14998
rect 8504 14942 8560 14998
rect 8628 14942 8684 14998
rect 8752 14942 8808 14998
rect 8876 14942 8932 14998
rect 9000 14942 9056 14998
rect 9124 14942 9180 14998
rect 9248 14942 9304 14998
rect 9372 14942 9428 14998
rect 9496 14942 9552 14998
rect 9620 14942 9676 14998
rect 9744 14942 9800 14998
rect 7884 14818 7940 14874
rect 8008 14818 8064 14874
rect 8132 14818 8188 14874
rect 8256 14818 8312 14874
rect 8380 14818 8436 14874
rect 8504 14818 8560 14874
rect 8628 14818 8684 14874
rect 8752 14818 8808 14874
rect 8876 14818 8932 14874
rect 9000 14818 9056 14874
rect 9124 14818 9180 14874
rect 9248 14818 9304 14874
rect 9372 14818 9428 14874
rect 9496 14818 9552 14874
rect 9620 14818 9676 14874
rect 9744 14818 9800 14874
rect 7884 14694 7940 14750
rect 8008 14694 8064 14750
rect 8132 14694 8188 14750
rect 8256 14694 8312 14750
rect 8380 14694 8436 14750
rect 8504 14694 8560 14750
rect 8628 14694 8684 14750
rect 8752 14694 8808 14750
rect 8876 14694 8932 14750
rect 9000 14694 9056 14750
rect 9124 14694 9180 14750
rect 9248 14694 9304 14750
rect 9372 14694 9428 14750
rect 9496 14694 9552 14750
rect 9620 14694 9676 14750
rect 9744 14694 9800 14750
rect 7884 14570 7940 14626
rect 8008 14570 8064 14626
rect 8132 14570 8188 14626
rect 8256 14570 8312 14626
rect 8380 14570 8436 14626
rect 8504 14570 8560 14626
rect 8628 14570 8684 14626
rect 8752 14570 8808 14626
rect 8876 14570 8932 14626
rect 9000 14570 9056 14626
rect 9124 14570 9180 14626
rect 9248 14570 9304 14626
rect 9372 14570 9428 14626
rect 9496 14570 9552 14626
rect 9620 14570 9676 14626
rect 9744 14570 9800 14626
rect 7884 14446 7940 14502
rect 8008 14446 8064 14502
rect 8132 14446 8188 14502
rect 8256 14446 8312 14502
rect 8380 14446 8436 14502
rect 8504 14446 8560 14502
rect 8628 14446 8684 14502
rect 8752 14446 8808 14502
rect 8876 14446 8932 14502
rect 9000 14446 9056 14502
rect 9124 14446 9180 14502
rect 9248 14446 9304 14502
rect 9372 14446 9428 14502
rect 9496 14446 9552 14502
rect 9620 14446 9676 14502
rect 9744 14446 9800 14502
rect 10254 17298 10310 17354
rect 10378 17298 10434 17354
rect 10502 17298 10558 17354
rect 10626 17298 10682 17354
rect 10750 17298 10806 17354
rect 10874 17298 10930 17354
rect 10998 17298 11054 17354
rect 11122 17298 11178 17354
rect 11246 17298 11302 17354
rect 11370 17298 11426 17354
rect 11494 17298 11550 17354
rect 11618 17298 11674 17354
rect 11742 17298 11798 17354
rect 11866 17298 11922 17354
rect 11990 17298 12046 17354
rect 12114 17298 12170 17354
rect 10254 17174 10310 17230
rect 10378 17174 10434 17230
rect 10502 17174 10558 17230
rect 10626 17174 10682 17230
rect 10750 17174 10806 17230
rect 10874 17174 10930 17230
rect 10998 17174 11054 17230
rect 11122 17174 11178 17230
rect 11246 17174 11302 17230
rect 11370 17174 11426 17230
rect 11494 17174 11550 17230
rect 11618 17174 11674 17230
rect 11742 17174 11798 17230
rect 11866 17174 11922 17230
rect 11990 17174 12046 17230
rect 12114 17174 12170 17230
rect 10254 17050 10310 17106
rect 10378 17050 10434 17106
rect 10502 17050 10558 17106
rect 10626 17050 10682 17106
rect 10750 17050 10806 17106
rect 10874 17050 10930 17106
rect 10998 17050 11054 17106
rect 11122 17050 11178 17106
rect 11246 17050 11302 17106
rect 11370 17050 11426 17106
rect 11494 17050 11550 17106
rect 11618 17050 11674 17106
rect 11742 17050 11798 17106
rect 11866 17050 11922 17106
rect 11990 17050 12046 17106
rect 12114 17050 12170 17106
rect 10254 16926 10310 16982
rect 10378 16926 10434 16982
rect 10502 16926 10558 16982
rect 10626 16926 10682 16982
rect 10750 16926 10806 16982
rect 10874 16926 10930 16982
rect 10998 16926 11054 16982
rect 11122 16926 11178 16982
rect 11246 16926 11302 16982
rect 11370 16926 11426 16982
rect 11494 16926 11550 16982
rect 11618 16926 11674 16982
rect 11742 16926 11798 16982
rect 11866 16926 11922 16982
rect 11990 16926 12046 16982
rect 12114 16926 12170 16982
rect 10254 16802 10310 16858
rect 10378 16802 10434 16858
rect 10502 16802 10558 16858
rect 10626 16802 10682 16858
rect 10750 16802 10806 16858
rect 10874 16802 10930 16858
rect 10998 16802 11054 16858
rect 11122 16802 11178 16858
rect 11246 16802 11302 16858
rect 11370 16802 11426 16858
rect 11494 16802 11550 16858
rect 11618 16802 11674 16858
rect 11742 16802 11798 16858
rect 11866 16802 11922 16858
rect 11990 16802 12046 16858
rect 12114 16802 12170 16858
rect 10254 16678 10310 16734
rect 10378 16678 10434 16734
rect 10502 16678 10558 16734
rect 10626 16678 10682 16734
rect 10750 16678 10806 16734
rect 10874 16678 10930 16734
rect 10998 16678 11054 16734
rect 11122 16678 11178 16734
rect 11246 16678 11302 16734
rect 11370 16678 11426 16734
rect 11494 16678 11550 16734
rect 11618 16678 11674 16734
rect 11742 16678 11798 16734
rect 11866 16678 11922 16734
rect 11990 16678 12046 16734
rect 12114 16678 12170 16734
rect 10254 16554 10310 16610
rect 10378 16554 10434 16610
rect 10502 16554 10558 16610
rect 10626 16554 10682 16610
rect 10750 16554 10806 16610
rect 10874 16554 10930 16610
rect 10998 16554 11054 16610
rect 11122 16554 11178 16610
rect 11246 16554 11302 16610
rect 11370 16554 11426 16610
rect 11494 16554 11550 16610
rect 11618 16554 11674 16610
rect 11742 16554 11798 16610
rect 11866 16554 11922 16610
rect 11990 16554 12046 16610
rect 12114 16554 12170 16610
rect 10254 16430 10310 16486
rect 10378 16430 10434 16486
rect 10502 16430 10558 16486
rect 10626 16430 10682 16486
rect 10750 16430 10806 16486
rect 10874 16430 10930 16486
rect 10998 16430 11054 16486
rect 11122 16430 11178 16486
rect 11246 16430 11302 16486
rect 11370 16430 11426 16486
rect 11494 16430 11550 16486
rect 11618 16430 11674 16486
rect 11742 16430 11798 16486
rect 11866 16430 11922 16486
rect 11990 16430 12046 16486
rect 12114 16430 12170 16486
rect 10254 16306 10310 16362
rect 10378 16306 10434 16362
rect 10502 16306 10558 16362
rect 10626 16306 10682 16362
rect 10750 16306 10806 16362
rect 10874 16306 10930 16362
rect 10998 16306 11054 16362
rect 11122 16306 11178 16362
rect 11246 16306 11302 16362
rect 11370 16306 11426 16362
rect 11494 16306 11550 16362
rect 11618 16306 11674 16362
rect 11742 16306 11798 16362
rect 11866 16306 11922 16362
rect 11990 16306 12046 16362
rect 12114 16306 12170 16362
rect 10254 16182 10310 16238
rect 10378 16182 10434 16238
rect 10502 16182 10558 16238
rect 10626 16182 10682 16238
rect 10750 16182 10806 16238
rect 10874 16182 10930 16238
rect 10998 16182 11054 16238
rect 11122 16182 11178 16238
rect 11246 16182 11302 16238
rect 11370 16182 11426 16238
rect 11494 16182 11550 16238
rect 11618 16182 11674 16238
rect 11742 16182 11798 16238
rect 11866 16182 11922 16238
rect 11990 16182 12046 16238
rect 12114 16182 12170 16238
rect 10254 16058 10310 16114
rect 10378 16058 10434 16114
rect 10502 16058 10558 16114
rect 10626 16058 10682 16114
rect 10750 16058 10806 16114
rect 10874 16058 10930 16114
rect 10998 16058 11054 16114
rect 11122 16058 11178 16114
rect 11246 16058 11302 16114
rect 11370 16058 11426 16114
rect 11494 16058 11550 16114
rect 11618 16058 11674 16114
rect 11742 16058 11798 16114
rect 11866 16058 11922 16114
rect 11990 16058 12046 16114
rect 12114 16058 12170 16114
rect 10254 15934 10310 15990
rect 10378 15934 10434 15990
rect 10502 15934 10558 15990
rect 10626 15934 10682 15990
rect 10750 15934 10806 15990
rect 10874 15934 10930 15990
rect 10998 15934 11054 15990
rect 11122 15934 11178 15990
rect 11246 15934 11302 15990
rect 11370 15934 11426 15990
rect 11494 15934 11550 15990
rect 11618 15934 11674 15990
rect 11742 15934 11798 15990
rect 11866 15934 11922 15990
rect 11990 15934 12046 15990
rect 12114 15934 12170 15990
rect 10254 15810 10310 15866
rect 10378 15810 10434 15866
rect 10502 15810 10558 15866
rect 10626 15810 10682 15866
rect 10750 15810 10806 15866
rect 10874 15810 10930 15866
rect 10998 15810 11054 15866
rect 11122 15810 11178 15866
rect 11246 15810 11302 15866
rect 11370 15810 11426 15866
rect 11494 15810 11550 15866
rect 11618 15810 11674 15866
rect 11742 15810 11798 15866
rect 11866 15810 11922 15866
rect 11990 15810 12046 15866
rect 12114 15810 12170 15866
rect 10254 15686 10310 15742
rect 10378 15686 10434 15742
rect 10502 15686 10558 15742
rect 10626 15686 10682 15742
rect 10750 15686 10806 15742
rect 10874 15686 10930 15742
rect 10998 15686 11054 15742
rect 11122 15686 11178 15742
rect 11246 15686 11302 15742
rect 11370 15686 11426 15742
rect 11494 15686 11550 15742
rect 11618 15686 11674 15742
rect 11742 15686 11798 15742
rect 11866 15686 11922 15742
rect 11990 15686 12046 15742
rect 12114 15686 12170 15742
rect 10254 15562 10310 15618
rect 10378 15562 10434 15618
rect 10502 15562 10558 15618
rect 10626 15562 10682 15618
rect 10750 15562 10806 15618
rect 10874 15562 10930 15618
rect 10998 15562 11054 15618
rect 11122 15562 11178 15618
rect 11246 15562 11302 15618
rect 11370 15562 11426 15618
rect 11494 15562 11550 15618
rect 11618 15562 11674 15618
rect 11742 15562 11798 15618
rect 11866 15562 11922 15618
rect 11990 15562 12046 15618
rect 12114 15562 12170 15618
rect 10254 15438 10310 15494
rect 10378 15438 10434 15494
rect 10502 15438 10558 15494
rect 10626 15438 10682 15494
rect 10750 15438 10806 15494
rect 10874 15438 10930 15494
rect 10998 15438 11054 15494
rect 11122 15438 11178 15494
rect 11246 15438 11302 15494
rect 11370 15438 11426 15494
rect 11494 15438 11550 15494
rect 11618 15438 11674 15494
rect 11742 15438 11798 15494
rect 11866 15438 11922 15494
rect 11990 15438 12046 15494
rect 12114 15438 12170 15494
rect 10254 15314 10310 15370
rect 10378 15314 10434 15370
rect 10502 15314 10558 15370
rect 10626 15314 10682 15370
rect 10750 15314 10806 15370
rect 10874 15314 10930 15370
rect 10998 15314 11054 15370
rect 11122 15314 11178 15370
rect 11246 15314 11302 15370
rect 11370 15314 11426 15370
rect 11494 15314 11550 15370
rect 11618 15314 11674 15370
rect 11742 15314 11798 15370
rect 11866 15314 11922 15370
rect 11990 15314 12046 15370
rect 12114 15314 12170 15370
rect 10254 15190 10310 15246
rect 10378 15190 10434 15246
rect 10502 15190 10558 15246
rect 10626 15190 10682 15246
rect 10750 15190 10806 15246
rect 10874 15190 10930 15246
rect 10998 15190 11054 15246
rect 11122 15190 11178 15246
rect 11246 15190 11302 15246
rect 11370 15190 11426 15246
rect 11494 15190 11550 15246
rect 11618 15190 11674 15246
rect 11742 15190 11798 15246
rect 11866 15190 11922 15246
rect 11990 15190 12046 15246
rect 12114 15190 12170 15246
rect 10254 15066 10310 15122
rect 10378 15066 10434 15122
rect 10502 15066 10558 15122
rect 10626 15066 10682 15122
rect 10750 15066 10806 15122
rect 10874 15066 10930 15122
rect 10998 15066 11054 15122
rect 11122 15066 11178 15122
rect 11246 15066 11302 15122
rect 11370 15066 11426 15122
rect 11494 15066 11550 15122
rect 11618 15066 11674 15122
rect 11742 15066 11798 15122
rect 11866 15066 11922 15122
rect 11990 15066 12046 15122
rect 12114 15066 12170 15122
rect 10254 14942 10310 14998
rect 10378 14942 10434 14998
rect 10502 14942 10558 14998
rect 10626 14942 10682 14998
rect 10750 14942 10806 14998
rect 10874 14942 10930 14998
rect 10998 14942 11054 14998
rect 11122 14942 11178 14998
rect 11246 14942 11302 14998
rect 11370 14942 11426 14998
rect 11494 14942 11550 14998
rect 11618 14942 11674 14998
rect 11742 14942 11798 14998
rect 11866 14942 11922 14998
rect 11990 14942 12046 14998
rect 12114 14942 12170 14998
rect 10254 14818 10310 14874
rect 10378 14818 10434 14874
rect 10502 14818 10558 14874
rect 10626 14818 10682 14874
rect 10750 14818 10806 14874
rect 10874 14818 10930 14874
rect 10998 14818 11054 14874
rect 11122 14818 11178 14874
rect 11246 14818 11302 14874
rect 11370 14818 11426 14874
rect 11494 14818 11550 14874
rect 11618 14818 11674 14874
rect 11742 14818 11798 14874
rect 11866 14818 11922 14874
rect 11990 14818 12046 14874
rect 12114 14818 12170 14874
rect 10254 14694 10310 14750
rect 10378 14694 10434 14750
rect 10502 14694 10558 14750
rect 10626 14694 10682 14750
rect 10750 14694 10806 14750
rect 10874 14694 10930 14750
rect 10998 14694 11054 14750
rect 11122 14694 11178 14750
rect 11246 14694 11302 14750
rect 11370 14694 11426 14750
rect 11494 14694 11550 14750
rect 11618 14694 11674 14750
rect 11742 14694 11798 14750
rect 11866 14694 11922 14750
rect 11990 14694 12046 14750
rect 12114 14694 12170 14750
rect 10254 14570 10310 14626
rect 10378 14570 10434 14626
rect 10502 14570 10558 14626
rect 10626 14570 10682 14626
rect 10750 14570 10806 14626
rect 10874 14570 10930 14626
rect 10998 14570 11054 14626
rect 11122 14570 11178 14626
rect 11246 14570 11302 14626
rect 11370 14570 11426 14626
rect 11494 14570 11550 14626
rect 11618 14570 11674 14626
rect 11742 14570 11798 14626
rect 11866 14570 11922 14626
rect 11990 14570 12046 14626
rect 12114 14570 12170 14626
rect 10254 14446 10310 14502
rect 10378 14446 10434 14502
rect 10502 14446 10558 14502
rect 10626 14446 10682 14502
rect 10750 14446 10806 14502
rect 10874 14446 10930 14502
rect 10998 14446 11054 14502
rect 11122 14446 11178 14502
rect 11246 14446 11302 14502
rect 11370 14446 11426 14502
rect 11494 14446 11550 14502
rect 11618 14446 11674 14502
rect 11742 14446 11798 14502
rect 11866 14446 11922 14502
rect 11990 14446 12046 14502
rect 12114 14446 12170 14502
rect 12871 17298 12927 17354
rect 12995 17298 13051 17354
rect 13119 17298 13175 17354
rect 13243 17298 13299 17354
rect 13367 17298 13423 17354
rect 13491 17298 13547 17354
rect 13615 17298 13671 17354
rect 13739 17298 13795 17354
rect 13863 17298 13919 17354
rect 13987 17298 14043 17354
rect 14111 17298 14167 17354
rect 14235 17298 14291 17354
rect 14359 17298 14415 17354
rect 14483 17298 14539 17354
rect 14607 17298 14663 17354
rect 12871 17174 12927 17230
rect 12995 17174 13051 17230
rect 13119 17174 13175 17230
rect 13243 17174 13299 17230
rect 13367 17174 13423 17230
rect 13491 17174 13547 17230
rect 13615 17174 13671 17230
rect 13739 17174 13795 17230
rect 13863 17174 13919 17230
rect 13987 17174 14043 17230
rect 14111 17174 14167 17230
rect 14235 17174 14291 17230
rect 14359 17174 14415 17230
rect 14483 17174 14539 17230
rect 14607 17174 14663 17230
rect 12871 17050 12927 17106
rect 12995 17050 13051 17106
rect 13119 17050 13175 17106
rect 13243 17050 13299 17106
rect 13367 17050 13423 17106
rect 13491 17050 13547 17106
rect 13615 17050 13671 17106
rect 13739 17050 13795 17106
rect 13863 17050 13919 17106
rect 13987 17050 14043 17106
rect 14111 17050 14167 17106
rect 14235 17050 14291 17106
rect 14359 17050 14415 17106
rect 14483 17050 14539 17106
rect 14607 17050 14663 17106
rect 12871 16926 12927 16982
rect 12995 16926 13051 16982
rect 13119 16926 13175 16982
rect 13243 16926 13299 16982
rect 13367 16926 13423 16982
rect 13491 16926 13547 16982
rect 13615 16926 13671 16982
rect 13739 16926 13795 16982
rect 13863 16926 13919 16982
rect 13987 16926 14043 16982
rect 14111 16926 14167 16982
rect 14235 16926 14291 16982
rect 14359 16926 14415 16982
rect 14483 16926 14539 16982
rect 14607 16926 14663 16982
rect 12871 16802 12927 16858
rect 12995 16802 13051 16858
rect 13119 16802 13175 16858
rect 13243 16802 13299 16858
rect 13367 16802 13423 16858
rect 13491 16802 13547 16858
rect 13615 16802 13671 16858
rect 13739 16802 13795 16858
rect 13863 16802 13919 16858
rect 13987 16802 14043 16858
rect 14111 16802 14167 16858
rect 14235 16802 14291 16858
rect 14359 16802 14415 16858
rect 14483 16802 14539 16858
rect 14607 16802 14663 16858
rect 12871 16678 12927 16734
rect 12995 16678 13051 16734
rect 13119 16678 13175 16734
rect 13243 16678 13299 16734
rect 13367 16678 13423 16734
rect 13491 16678 13547 16734
rect 13615 16678 13671 16734
rect 13739 16678 13795 16734
rect 13863 16678 13919 16734
rect 13987 16678 14043 16734
rect 14111 16678 14167 16734
rect 14235 16678 14291 16734
rect 14359 16678 14415 16734
rect 14483 16678 14539 16734
rect 14607 16678 14663 16734
rect 12871 16554 12927 16610
rect 12995 16554 13051 16610
rect 13119 16554 13175 16610
rect 13243 16554 13299 16610
rect 13367 16554 13423 16610
rect 13491 16554 13547 16610
rect 13615 16554 13671 16610
rect 13739 16554 13795 16610
rect 13863 16554 13919 16610
rect 13987 16554 14043 16610
rect 14111 16554 14167 16610
rect 14235 16554 14291 16610
rect 14359 16554 14415 16610
rect 14483 16554 14539 16610
rect 14607 16554 14663 16610
rect 12871 16430 12927 16486
rect 12995 16430 13051 16486
rect 13119 16430 13175 16486
rect 13243 16430 13299 16486
rect 13367 16430 13423 16486
rect 13491 16430 13547 16486
rect 13615 16430 13671 16486
rect 13739 16430 13795 16486
rect 13863 16430 13919 16486
rect 13987 16430 14043 16486
rect 14111 16430 14167 16486
rect 14235 16430 14291 16486
rect 14359 16430 14415 16486
rect 14483 16430 14539 16486
rect 14607 16430 14663 16486
rect 12871 16306 12927 16362
rect 12995 16306 13051 16362
rect 13119 16306 13175 16362
rect 13243 16306 13299 16362
rect 13367 16306 13423 16362
rect 13491 16306 13547 16362
rect 13615 16306 13671 16362
rect 13739 16306 13795 16362
rect 13863 16306 13919 16362
rect 13987 16306 14043 16362
rect 14111 16306 14167 16362
rect 14235 16306 14291 16362
rect 14359 16306 14415 16362
rect 14483 16306 14539 16362
rect 14607 16306 14663 16362
rect 12871 16182 12927 16238
rect 12995 16182 13051 16238
rect 13119 16182 13175 16238
rect 13243 16182 13299 16238
rect 13367 16182 13423 16238
rect 13491 16182 13547 16238
rect 13615 16182 13671 16238
rect 13739 16182 13795 16238
rect 13863 16182 13919 16238
rect 13987 16182 14043 16238
rect 14111 16182 14167 16238
rect 14235 16182 14291 16238
rect 14359 16182 14415 16238
rect 14483 16182 14539 16238
rect 14607 16182 14663 16238
rect 12871 16058 12927 16114
rect 12995 16058 13051 16114
rect 13119 16058 13175 16114
rect 13243 16058 13299 16114
rect 13367 16058 13423 16114
rect 13491 16058 13547 16114
rect 13615 16058 13671 16114
rect 13739 16058 13795 16114
rect 13863 16058 13919 16114
rect 13987 16058 14043 16114
rect 14111 16058 14167 16114
rect 14235 16058 14291 16114
rect 14359 16058 14415 16114
rect 14483 16058 14539 16114
rect 14607 16058 14663 16114
rect 12871 15934 12927 15990
rect 12995 15934 13051 15990
rect 13119 15934 13175 15990
rect 13243 15934 13299 15990
rect 13367 15934 13423 15990
rect 13491 15934 13547 15990
rect 13615 15934 13671 15990
rect 13739 15934 13795 15990
rect 13863 15934 13919 15990
rect 13987 15934 14043 15990
rect 14111 15934 14167 15990
rect 14235 15934 14291 15990
rect 14359 15934 14415 15990
rect 14483 15934 14539 15990
rect 14607 15934 14663 15990
rect 12871 15810 12927 15866
rect 12995 15810 13051 15866
rect 13119 15810 13175 15866
rect 13243 15810 13299 15866
rect 13367 15810 13423 15866
rect 13491 15810 13547 15866
rect 13615 15810 13671 15866
rect 13739 15810 13795 15866
rect 13863 15810 13919 15866
rect 13987 15810 14043 15866
rect 14111 15810 14167 15866
rect 14235 15810 14291 15866
rect 14359 15810 14415 15866
rect 14483 15810 14539 15866
rect 14607 15810 14663 15866
rect 12871 15686 12927 15742
rect 12995 15686 13051 15742
rect 13119 15686 13175 15742
rect 13243 15686 13299 15742
rect 13367 15686 13423 15742
rect 13491 15686 13547 15742
rect 13615 15686 13671 15742
rect 13739 15686 13795 15742
rect 13863 15686 13919 15742
rect 13987 15686 14043 15742
rect 14111 15686 14167 15742
rect 14235 15686 14291 15742
rect 14359 15686 14415 15742
rect 14483 15686 14539 15742
rect 14607 15686 14663 15742
rect 12871 15562 12927 15618
rect 12995 15562 13051 15618
rect 13119 15562 13175 15618
rect 13243 15562 13299 15618
rect 13367 15562 13423 15618
rect 13491 15562 13547 15618
rect 13615 15562 13671 15618
rect 13739 15562 13795 15618
rect 13863 15562 13919 15618
rect 13987 15562 14043 15618
rect 14111 15562 14167 15618
rect 14235 15562 14291 15618
rect 14359 15562 14415 15618
rect 14483 15562 14539 15618
rect 14607 15562 14663 15618
rect 12871 15438 12927 15494
rect 12995 15438 13051 15494
rect 13119 15438 13175 15494
rect 13243 15438 13299 15494
rect 13367 15438 13423 15494
rect 13491 15438 13547 15494
rect 13615 15438 13671 15494
rect 13739 15438 13795 15494
rect 13863 15438 13919 15494
rect 13987 15438 14043 15494
rect 14111 15438 14167 15494
rect 14235 15438 14291 15494
rect 14359 15438 14415 15494
rect 14483 15438 14539 15494
rect 14607 15438 14663 15494
rect 12871 15314 12927 15370
rect 12995 15314 13051 15370
rect 13119 15314 13175 15370
rect 13243 15314 13299 15370
rect 13367 15314 13423 15370
rect 13491 15314 13547 15370
rect 13615 15314 13671 15370
rect 13739 15314 13795 15370
rect 13863 15314 13919 15370
rect 13987 15314 14043 15370
rect 14111 15314 14167 15370
rect 14235 15314 14291 15370
rect 14359 15314 14415 15370
rect 14483 15314 14539 15370
rect 14607 15314 14663 15370
rect 12871 15190 12927 15246
rect 12995 15190 13051 15246
rect 13119 15190 13175 15246
rect 13243 15190 13299 15246
rect 13367 15190 13423 15246
rect 13491 15190 13547 15246
rect 13615 15190 13671 15246
rect 13739 15190 13795 15246
rect 13863 15190 13919 15246
rect 13987 15190 14043 15246
rect 14111 15190 14167 15246
rect 14235 15190 14291 15246
rect 14359 15190 14415 15246
rect 14483 15190 14539 15246
rect 14607 15190 14663 15246
rect 12871 15066 12927 15122
rect 12995 15066 13051 15122
rect 13119 15066 13175 15122
rect 13243 15066 13299 15122
rect 13367 15066 13423 15122
rect 13491 15066 13547 15122
rect 13615 15066 13671 15122
rect 13739 15066 13795 15122
rect 13863 15066 13919 15122
rect 13987 15066 14043 15122
rect 14111 15066 14167 15122
rect 14235 15066 14291 15122
rect 14359 15066 14415 15122
rect 14483 15066 14539 15122
rect 14607 15066 14663 15122
rect 12871 14942 12927 14998
rect 12995 14942 13051 14998
rect 13119 14942 13175 14998
rect 13243 14942 13299 14998
rect 13367 14942 13423 14998
rect 13491 14942 13547 14998
rect 13615 14942 13671 14998
rect 13739 14942 13795 14998
rect 13863 14942 13919 14998
rect 13987 14942 14043 14998
rect 14111 14942 14167 14998
rect 14235 14942 14291 14998
rect 14359 14942 14415 14998
rect 14483 14942 14539 14998
rect 14607 14942 14663 14998
rect 12871 14818 12927 14874
rect 12995 14818 13051 14874
rect 13119 14818 13175 14874
rect 13243 14818 13299 14874
rect 13367 14818 13423 14874
rect 13491 14818 13547 14874
rect 13615 14818 13671 14874
rect 13739 14818 13795 14874
rect 13863 14818 13919 14874
rect 13987 14818 14043 14874
rect 14111 14818 14167 14874
rect 14235 14818 14291 14874
rect 14359 14818 14415 14874
rect 14483 14818 14539 14874
rect 14607 14818 14663 14874
rect 12871 14694 12927 14750
rect 12995 14694 13051 14750
rect 13119 14694 13175 14750
rect 13243 14694 13299 14750
rect 13367 14694 13423 14750
rect 13491 14694 13547 14750
rect 13615 14694 13671 14750
rect 13739 14694 13795 14750
rect 13863 14694 13919 14750
rect 13987 14694 14043 14750
rect 14111 14694 14167 14750
rect 14235 14694 14291 14750
rect 14359 14694 14415 14750
rect 14483 14694 14539 14750
rect 14607 14694 14663 14750
rect 12871 14570 12927 14626
rect 12995 14570 13051 14626
rect 13119 14570 13175 14626
rect 13243 14570 13299 14626
rect 13367 14570 13423 14626
rect 13491 14570 13547 14626
rect 13615 14570 13671 14626
rect 13739 14570 13795 14626
rect 13863 14570 13919 14626
rect 13987 14570 14043 14626
rect 14111 14570 14167 14626
rect 14235 14570 14291 14626
rect 14359 14570 14415 14626
rect 14483 14570 14539 14626
rect 14607 14570 14663 14626
rect 12871 14446 12927 14502
rect 12995 14446 13051 14502
rect 13119 14446 13175 14502
rect 13243 14446 13299 14502
rect 13367 14446 13423 14502
rect 13491 14446 13547 14502
rect 13615 14446 13671 14502
rect 13739 14446 13795 14502
rect 13863 14446 13919 14502
rect 13987 14446 14043 14502
rect 14111 14446 14167 14502
rect 14235 14446 14291 14502
rect 14359 14446 14415 14502
rect 14483 14446 14539 14502
rect 14607 14446 14663 14502
rect 2491 14092 2547 14148
rect 2615 14092 2671 14148
rect 2491 13968 2547 14024
rect 2615 13968 2671 14024
rect 2491 13844 2547 13900
rect 2615 13844 2671 13900
rect 2491 13720 2547 13776
rect 2615 13720 2671 13776
rect 2491 13596 2547 13652
rect 2615 13596 2671 13652
rect 2491 13472 2547 13528
rect 2615 13472 2671 13528
rect 2491 13348 2547 13404
rect 2615 13348 2671 13404
rect 2491 13224 2547 13280
rect 2615 13224 2671 13280
rect 2491 13100 2547 13156
rect 2615 13100 2671 13156
rect 2491 12976 2547 13032
rect 2615 12976 2671 13032
rect 2491 12852 2547 12908
rect 2615 12852 2671 12908
rect 4861 14092 4917 14148
rect 4985 14092 5041 14148
rect 4861 13968 4917 14024
rect 4985 13968 5041 14024
rect 4861 13844 4917 13900
rect 4985 13844 5041 13900
rect 4861 13720 4917 13776
rect 4985 13720 5041 13776
rect 4861 13596 4917 13652
rect 4985 13596 5041 13652
rect 4861 13472 4917 13528
rect 4985 13472 5041 13528
rect 4861 13348 4917 13404
rect 4985 13348 5041 13404
rect 4861 13224 4917 13280
rect 4985 13224 5041 13280
rect 4861 13100 4917 13156
rect 4985 13100 5041 13156
rect 4861 12976 4917 13032
rect 4985 12976 5041 13032
rect 4861 12852 4917 12908
rect 4985 12852 5041 12908
rect 7275 14092 7331 14148
rect 7399 14092 7455 14148
rect 7523 14092 7579 14148
rect 7647 14092 7703 14148
rect 7275 13968 7331 14024
rect 7399 13968 7455 14024
rect 7523 13968 7579 14024
rect 7647 13968 7703 14024
rect 7275 13844 7331 13900
rect 7399 13844 7455 13900
rect 7523 13844 7579 13900
rect 7647 13844 7703 13900
rect 7275 13720 7331 13776
rect 7399 13720 7455 13776
rect 7523 13720 7579 13776
rect 7647 13720 7703 13776
rect 7275 13596 7331 13652
rect 7399 13596 7455 13652
rect 7523 13596 7579 13652
rect 7647 13596 7703 13652
rect 7275 13472 7331 13528
rect 7399 13472 7455 13528
rect 7523 13472 7579 13528
rect 7647 13472 7703 13528
rect 7275 13348 7331 13404
rect 7399 13348 7455 13404
rect 7523 13348 7579 13404
rect 7647 13348 7703 13404
rect 7275 13224 7331 13280
rect 7399 13224 7455 13280
rect 7523 13224 7579 13280
rect 7647 13224 7703 13280
rect 7275 13100 7331 13156
rect 7399 13100 7455 13156
rect 7523 13100 7579 13156
rect 7647 13100 7703 13156
rect 7275 12976 7331 13032
rect 7399 12976 7455 13032
rect 7523 12976 7579 13032
rect 7647 12976 7703 13032
rect 7275 12852 7331 12908
rect 7399 12852 7455 12908
rect 7523 12852 7579 12908
rect 7647 12852 7703 12908
rect 9937 14092 9993 14148
rect 10061 14092 10117 14148
rect 9937 13968 9993 14024
rect 10061 13968 10117 14024
rect 9937 13844 9993 13900
rect 10061 13844 10117 13900
rect 9937 13720 9993 13776
rect 10061 13720 10117 13776
rect 9937 13596 9993 13652
rect 10061 13596 10117 13652
rect 9937 13472 9993 13528
rect 10061 13472 10117 13528
rect 9937 13348 9993 13404
rect 10061 13348 10117 13404
rect 9937 13224 9993 13280
rect 10061 13224 10117 13280
rect 9937 13100 9993 13156
rect 10061 13100 10117 13156
rect 9937 12976 9993 13032
rect 10061 12976 10117 13032
rect 9937 12852 9993 12908
rect 10061 12852 10117 12908
rect 12307 14092 12363 14148
rect 12431 14092 12487 14148
rect 12307 13968 12363 14024
rect 12431 13968 12487 14024
rect 12307 13844 12363 13900
rect 12431 13844 12487 13900
rect 12307 13720 12363 13776
rect 12431 13720 12487 13776
rect 12307 13596 12363 13652
rect 12431 13596 12487 13652
rect 12307 13472 12363 13528
rect 12431 13472 12487 13528
rect 12307 13348 12363 13404
rect 12431 13348 12487 13404
rect 12307 13224 12363 13280
rect 12431 13224 12487 13280
rect 12307 13100 12363 13156
rect 12431 13100 12487 13156
rect 12307 12976 12363 13032
rect 12431 12976 12487 13032
rect 12307 12852 12363 12908
rect 12431 12852 12487 12908
rect 315 12492 371 12548
rect 439 12492 495 12548
rect 563 12492 619 12548
rect 687 12492 743 12548
rect 811 12492 867 12548
rect 935 12492 991 12548
rect 1059 12492 1115 12548
rect 1183 12492 1239 12548
rect 1307 12492 1363 12548
rect 1431 12492 1487 12548
rect 1555 12492 1611 12548
rect 1679 12492 1735 12548
rect 1803 12492 1859 12548
rect 1927 12492 1983 12548
rect 2051 12492 2107 12548
rect 315 12368 371 12424
rect 439 12368 495 12424
rect 563 12368 619 12424
rect 687 12368 743 12424
rect 811 12368 867 12424
rect 935 12368 991 12424
rect 1059 12368 1115 12424
rect 1183 12368 1239 12424
rect 1307 12368 1363 12424
rect 1431 12368 1487 12424
rect 1555 12368 1611 12424
rect 1679 12368 1735 12424
rect 1803 12368 1859 12424
rect 1927 12368 1983 12424
rect 2051 12368 2107 12424
rect 315 12244 371 12300
rect 439 12244 495 12300
rect 563 12244 619 12300
rect 687 12244 743 12300
rect 811 12244 867 12300
rect 935 12244 991 12300
rect 1059 12244 1115 12300
rect 1183 12244 1239 12300
rect 1307 12244 1363 12300
rect 1431 12244 1487 12300
rect 1555 12244 1611 12300
rect 1679 12244 1735 12300
rect 1803 12244 1859 12300
rect 1927 12244 1983 12300
rect 2051 12244 2107 12300
rect 315 12120 371 12176
rect 439 12120 495 12176
rect 563 12120 619 12176
rect 687 12120 743 12176
rect 811 12120 867 12176
rect 935 12120 991 12176
rect 1059 12120 1115 12176
rect 1183 12120 1239 12176
rect 1307 12120 1363 12176
rect 1431 12120 1487 12176
rect 1555 12120 1611 12176
rect 1679 12120 1735 12176
rect 1803 12120 1859 12176
rect 1927 12120 1983 12176
rect 2051 12120 2107 12176
rect 315 11996 371 12052
rect 439 11996 495 12052
rect 563 11996 619 12052
rect 687 11996 743 12052
rect 811 11996 867 12052
rect 935 11996 991 12052
rect 1059 11996 1115 12052
rect 1183 11996 1239 12052
rect 1307 11996 1363 12052
rect 1431 11996 1487 12052
rect 1555 11996 1611 12052
rect 1679 11996 1735 12052
rect 1803 11996 1859 12052
rect 1927 11996 1983 12052
rect 2051 11996 2107 12052
rect 315 11872 371 11928
rect 439 11872 495 11928
rect 563 11872 619 11928
rect 687 11872 743 11928
rect 811 11872 867 11928
rect 935 11872 991 11928
rect 1059 11872 1115 11928
rect 1183 11872 1239 11928
rect 1307 11872 1363 11928
rect 1431 11872 1487 11928
rect 1555 11872 1611 11928
rect 1679 11872 1735 11928
rect 1803 11872 1859 11928
rect 1927 11872 1983 11928
rect 2051 11872 2107 11928
rect 315 11748 371 11804
rect 439 11748 495 11804
rect 563 11748 619 11804
rect 687 11748 743 11804
rect 811 11748 867 11804
rect 935 11748 991 11804
rect 1059 11748 1115 11804
rect 1183 11748 1239 11804
rect 1307 11748 1363 11804
rect 1431 11748 1487 11804
rect 1555 11748 1611 11804
rect 1679 11748 1735 11804
rect 1803 11748 1859 11804
rect 1927 11748 1983 11804
rect 2051 11748 2107 11804
rect 315 11624 371 11680
rect 439 11624 495 11680
rect 563 11624 619 11680
rect 687 11624 743 11680
rect 811 11624 867 11680
rect 935 11624 991 11680
rect 1059 11624 1115 11680
rect 1183 11624 1239 11680
rect 1307 11624 1363 11680
rect 1431 11624 1487 11680
rect 1555 11624 1611 11680
rect 1679 11624 1735 11680
rect 1803 11624 1859 11680
rect 1927 11624 1983 11680
rect 2051 11624 2107 11680
rect 315 11500 371 11556
rect 439 11500 495 11556
rect 563 11500 619 11556
rect 687 11500 743 11556
rect 811 11500 867 11556
rect 935 11500 991 11556
rect 1059 11500 1115 11556
rect 1183 11500 1239 11556
rect 1307 11500 1363 11556
rect 1431 11500 1487 11556
rect 1555 11500 1611 11556
rect 1679 11500 1735 11556
rect 1803 11500 1859 11556
rect 1927 11500 1983 11556
rect 2051 11500 2107 11556
rect 315 11376 371 11432
rect 439 11376 495 11432
rect 563 11376 619 11432
rect 687 11376 743 11432
rect 811 11376 867 11432
rect 935 11376 991 11432
rect 1059 11376 1115 11432
rect 1183 11376 1239 11432
rect 1307 11376 1363 11432
rect 1431 11376 1487 11432
rect 1555 11376 1611 11432
rect 1679 11376 1735 11432
rect 1803 11376 1859 11432
rect 1927 11376 1983 11432
rect 2051 11376 2107 11432
rect 315 11252 371 11308
rect 439 11252 495 11308
rect 563 11252 619 11308
rect 687 11252 743 11308
rect 811 11252 867 11308
rect 935 11252 991 11308
rect 1059 11252 1115 11308
rect 1183 11252 1239 11308
rect 1307 11252 1363 11308
rect 1431 11252 1487 11308
rect 1555 11252 1611 11308
rect 1679 11252 1735 11308
rect 1803 11252 1859 11308
rect 1927 11252 1983 11308
rect 2051 11252 2107 11308
rect 2808 12492 2864 12548
rect 2932 12492 2988 12548
rect 3056 12492 3112 12548
rect 3180 12492 3236 12548
rect 3304 12492 3360 12548
rect 3428 12492 3484 12548
rect 3552 12492 3608 12548
rect 3676 12492 3732 12548
rect 3800 12492 3856 12548
rect 3924 12492 3980 12548
rect 4048 12492 4104 12548
rect 4172 12492 4228 12548
rect 4296 12492 4352 12548
rect 4420 12492 4476 12548
rect 4544 12492 4600 12548
rect 4668 12492 4724 12548
rect 2808 12368 2864 12424
rect 2932 12368 2988 12424
rect 3056 12368 3112 12424
rect 3180 12368 3236 12424
rect 3304 12368 3360 12424
rect 3428 12368 3484 12424
rect 3552 12368 3608 12424
rect 3676 12368 3732 12424
rect 3800 12368 3856 12424
rect 3924 12368 3980 12424
rect 4048 12368 4104 12424
rect 4172 12368 4228 12424
rect 4296 12368 4352 12424
rect 4420 12368 4476 12424
rect 4544 12368 4600 12424
rect 4668 12368 4724 12424
rect 2808 12244 2864 12300
rect 2932 12244 2988 12300
rect 3056 12244 3112 12300
rect 3180 12244 3236 12300
rect 3304 12244 3360 12300
rect 3428 12244 3484 12300
rect 3552 12244 3608 12300
rect 3676 12244 3732 12300
rect 3800 12244 3856 12300
rect 3924 12244 3980 12300
rect 4048 12244 4104 12300
rect 4172 12244 4228 12300
rect 4296 12244 4352 12300
rect 4420 12244 4476 12300
rect 4544 12244 4600 12300
rect 4668 12244 4724 12300
rect 2808 12120 2864 12176
rect 2932 12120 2988 12176
rect 3056 12120 3112 12176
rect 3180 12120 3236 12176
rect 3304 12120 3360 12176
rect 3428 12120 3484 12176
rect 3552 12120 3608 12176
rect 3676 12120 3732 12176
rect 3800 12120 3856 12176
rect 3924 12120 3980 12176
rect 4048 12120 4104 12176
rect 4172 12120 4228 12176
rect 4296 12120 4352 12176
rect 4420 12120 4476 12176
rect 4544 12120 4600 12176
rect 4668 12120 4724 12176
rect 2808 11996 2864 12052
rect 2932 11996 2988 12052
rect 3056 11996 3112 12052
rect 3180 11996 3236 12052
rect 3304 11996 3360 12052
rect 3428 11996 3484 12052
rect 3552 11996 3608 12052
rect 3676 11996 3732 12052
rect 3800 11996 3856 12052
rect 3924 11996 3980 12052
rect 4048 11996 4104 12052
rect 4172 11996 4228 12052
rect 4296 11996 4352 12052
rect 4420 11996 4476 12052
rect 4544 11996 4600 12052
rect 4668 11996 4724 12052
rect 2808 11872 2864 11928
rect 2932 11872 2988 11928
rect 3056 11872 3112 11928
rect 3180 11872 3236 11928
rect 3304 11872 3360 11928
rect 3428 11872 3484 11928
rect 3552 11872 3608 11928
rect 3676 11872 3732 11928
rect 3800 11872 3856 11928
rect 3924 11872 3980 11928
rect 4048 11872 4104 11928
rect 4172 11872 4228 11928
rect 4296 11872 4352 11928
rect 4420 11872 4476 11928
rect 4544 11872 4600 11928
rect 4668 11872 4724 11928
rect 2808 11748 2864 11804
rect 2932 11748 2988 11804
rect 3056 11748 3112 11804
rect 3180 11748 3236 11804
rect 3304 11748 3360 11804
rect 3428 11748 3484 11804
rect 3552 11748 3608 11804
rect 3676 11748 3732 11804
rect 3800 11748 3856 11804
rect 3924 11748 3980 11804
rect 4048 11748 4104 11804
rect 4172 11748 4228 11804
rect 4296 11748 4352 11804
rect 4420 11748 4476 11804
rect 4544 11748 4600 11804
rect 4668 11748 4724 11804
rect 2808 11624 2864 11680
rect 2932 11624 2988 11680
rect 3056 11624 3112 11680
rect 3180 11624 3236 11680
rect 3304 11624 3360 11680
rect 3428 11624 3484 11680
rect 3552 11624 3608 11680
rect 3676 11624 3732 11680
rect 3800 11624 3856 11680
rect 3924 11624 3980 11680
rect 4048 11624 4104 11680
rect 4172 11624 4228 11680
rect 4296 11624 4352 11680
rect 4420 11624 4476 11680
rect 4544 11624 4600 11680
rect 4668 11624 4724 11680
rect 2808 11500 2864 11556
rect 2932 11500 2988 11556
rect 3056 11500 3112 11556
rect 3180 11500 3236 11556
rect 3304 11500 3360 11556
rect 3428 11500 3484 11556
rect 3552 11500 3608 11556
rect 3676 11500 3732 11556
rect 3800 11500 3856 11556
rect 3924 11500 3980 11556
rect 4048 11500 4104 11556
rect 4172 11500 4228 11556
rect 4296 11500 4352 11556
rect 4420 11500 4476 11556
rect 4544 11500 4600 11556
rect 4668 11500 4724 11556
rect 2808 11376 2864 11432
rect 2932 11376 2988 11432
rect 3056 11376 3112 11432
rect 3180 11376 3236 11432
rect 3304 11376 3360 11432
rect 3428 11376 3484 11432
rect 3552 11376 3608 11432
rect 3676 11376 3732 11432
rect 3800 11376 3856 11432
rect 3924 11376 3980 11432
rect 4048 11376 4104 11432
rect 4172 11376 4228 11432
rect 4296 11376 4352 11432
rect 4420 11376 4476 11432
rect 4544 11376 4600 11432
rect 4668 11376 4724 11432
rect 2808 11252 2864 11308
rect 2932 11252 2988 11308
rect 3056 11252 3112 11308
rect 3180 11252 3236 11308
rect 3304 11252 3360 11308
rect 3428 11252 3484 11308
rect 3552 11252 3608 11308
rect 3676 11252 3732 11308
rect 3800 11252 3856 11308
rect 3924 11252 3980 11308
rect 4048 11252 4104 11308
rect 4172 11252 4228 11308
rect 4296 11252 4352 11308
rect 4420 11252 4476 11308
rect 4544 11252 4600 11308
rect 4668 11252 4724 11308
rect 5178 12492 5234 12548
rect 5302 12492 5358 12548
rect 5426 12492 5482 12548
rect 5550 12492 5606 12548
rect 5674 12492 5730 12548
rect 5798 12492 5854 12548
rect 5922 12492 5978 12548
rect 6046 12492 6102 12548
rect 6170 12492 6226 12548
rect 6294 12492 6350 12548
rect 6418 12492 6474 12548
rect 6542 12492 6598 12548
rect 6666 12492 6722 12548
rect 6790 12492 6846 12548
rect 6914 12492 6970 12548
rect 7038 12492 7094 12548
rect 5178 12368 5234 12424
rect 5302 12368 5358 12424
rect 5426 12368 5482 12424
rect 5550 12368 5606 12424
rect 5674 12368 5730 12424
rect 5798 12368 5854 12424
rect 5922 12368 5978 12424
rect 6046 12368 6102 12424
rect 6170 12368 6226 12424
rect 6294 12368 6350 12424
rect 6418 12368 6474 12424
rect 6542 12368 6598 12424
rect 6666 12368 6722 12424
rect 6790 12368 6846 12424
rect 6914 12368 6970 12424
rect 7038 12368 7094 12424
rect 5178 12244 5234 12300
rect 5302 12244 5358 12300
rect 5426 12244 5482 12300
rect 5550 12244 5606 12300
rect 5674 12244 5730 12300
rect 5798 12244 5854 12300
rect 5922 12244 5978 12300
rect 6046 12244 6102 12300
rect 6170 12244 6226 12300
rect 6294 12244 6350 12300
rect 6418 12244 6474 12300
rect 6542 12244 6598 12300
rect 6666 12244 6722 12300
rect 6790 12244 6846 12300
rect 6914 12244 6970 12300
rect 7038 12244 7094 12300
rect 5178 12120 5234 12176
rect 5302 12120 5358 12176
rect 5426 12120 5482 12176
rect 5550 12120 5606 12176
rect 5674 12120 5730 12176
rect 5798 12120 5854 12176
rect 5922 12120 5978 12176
rect 6046 12120 6102 12176
rect 6170 12120 6226 12176
rect 6294 12120 6350 12176
rect 6418 12120 6474 12176
rect 6542 12120 6598 12176
rect 6666 12120 6722 12176
rect 6790 12120 6846 12176
rect 6914 12120 6970 12176
rect 7038 12120 7094 12176
rect 5178 11996 5234 12052
rect 5302 11996 5358 12052
rect 5426 11996 5482 12052
rect 5550 11996 5606 12052
rect 5674 11996 5730 12052
rect 5798 11996 5854 12052
rect 5922 11996 5978 12052
rect 6046 11996 6102 12052
rect 6170 11996 6226 12052
rect 6294 11996 6350 12052
rect 6418 11996 6474 12052
rect 6542 11996 6598 12052
rect 6666 11996 6722 12052
rect 6790 11996 6846 12052
rect 6914 11996 6970 12052
rect 7038 11996 7094 12052
rect 5178 11872 5234 11928
rect 5302 11872 5358 11928
rect 5426 11872 5482 11928
rect 5550 11872 5606 11928
rect 5674 11872 5730 11928
rect 5798 11872 5854 11928
rect 5922 11872 5978 11928
rect 6046 11872 6102 11928
rect 6170 11872 6226 11928
rect 6294 11872 6350 11928
rect 6418 11872 6474 11928
rect 6542 11872 6598 11928
rect 6666 11872 6722 11928
rect 6790 11872 6846 11928
rect 6914 11872 6970 11928
rect 7038 11872 7094 11928
rect 5178 11748 5234 11804
rect 5302 11748 5358 11804
rect 5426 11748 5482 11804
rect 5550 11748 5606 11804
rect 5674 11748 5730 11804
rect 5798 11748 5854 11804
rect 5922 11748 5978 11804
rect 6046 11748 6102 11804
rect 6170 11748 6226 11804
rect 6294 11748 6350 11804
rect 6418 11748 6474 11804
rect 6542 11748 6598 11804
rect 6666 11748 6722 11804
rect 6790 11748 6846 11804
rect 6914 11748 6970 11804
rect 7038 11748 7094 11804
rect 5178 11624 5234 11680
rect 5302 11624 5358 11680
rect 5426 11624 5482 11680
rect 5550 11624 5606 11680
rect 5674 11624 5730 11680
rect 5798 11624 5854 11680
rect 5922 11624 5978 11680
rect 6046 11624 6102 11680
rect 6170 11624 6226 11680
rect 6294 11624 6350 11680
rect 6418 11624 6474 11680
rect 6542 11624 6598 11680
rect 6666 11624 6722 11680
rect 6790 11624 6846 11680
rect 6914 11624 6970 11680
rect 7038 11624 7094 11680
rect 5178 11500 5234 11556
rect 5302 11500 5358 11556
rect 5426 11500 5482 11556
rect 5550 11500 5606 11556
rect 5674 11500 5730 11556
rect 5798 11500 5854 11556
rect 5922 11500 5978 11556
rect 6046 11500 6102 11556
rect 6170 11500 6226 11556
rect 6294 11500 6350 11556
rect 6418 11500 6474 11556
rect 6542 11500 6598 11556
rect 6666 11500 6722 11556
rect 6790 11500 6846 11556
rect 6914 11500 6970 11556
rect 7038 11500 7094 11556
rect 5178 11376 5234 11432
rect 5302 11376 5358 11432
rect 5426 11376 5482 11432
rect 5550 11376 5606 11432
rect 5674 11376 5730 11432
rect 5798 11376 5854 11432
rect 5922 11376 5978 11432
rect 6046 11376 6102 11432
rect 6170 11376 6226 11432
rect 6294 11376 6350 11432
rect 6418 11376 6474 11432
rect 6542 11376 6598 11432
rect 6666 11376 6722 11432
rect 6790 11376 6846 11432
rect 6914 11376 6970 11432
rect 7038 11376 7094 11432
rect 5178 11252 5234 11308
rect 5302 11252 5358 11308
rect 5426 11252 5482 11308
rect 5550 11252 5606 11308
rect 5674 11252 5730 11308
rect 5798 11252 5854 11308
rect 5922 11252 5978 11308
rect 6046 11252 6102 11308
rect 6170 11252 6226 11308
rect 6294 11252 6350 11308
rect 6418 11252 6474 11308
rect 6542 11252 6598 11308
rect 6666 11252 6722 11308
rect 6790 11252 6846 11308
rect 6914 11252 6970 11308
rect 7038 11252 7094 11308
rect 7884 12492 7940 12548
rect 8008 12492 8064 12548
rect 8132 12492 8188 12548
rect 8256 12492 8312 12548
rect 8380 12492 8436 12548
rect 8504 12492 8560 12548
rect 8628 12492 8684 12548
rect 8752 12492 8808 12548
rect 8876 12492 8932 12548
rect 9000 12492 9056 12548
rect 9124 12492 9180 12548
rect 9248 12492 9304 12548
rect 9372 12492 9428 12548
rect 9496 12492 9552 12548
rect 9620 12492 9676 12548
rect 9744 12492 9800 12548
rect 7884 12368 7940 12424
rect 8008 12368 8064 12424
rect 8132 12368 8188 12424
rect 8256 12368 8312 12424
rect 8380 12368 8436 12424
rect 8504 12368 8560 12424
rect 8628 12368 8684 12424
rect 8752 12368 8808 12424
rect 8876 12368 8932 12424
rect 9000 12368 9056 12424
rect 9124 12368 9180 12424
rect 9248 12368 9304 12424
rect 9372 12368 9428 12424
rect 9496 12368 9552 12424
rect 9620 12368 9676 12424
rect 9744 12368 9800 12424
rect 7884 12244 7940 12300
rect 8008 12244 8064 12300
rect 8132 12244 8188 12300
rect 8256 12244 8312 12300
rect 8380 12244 8436 12300
rect 8504 12244 8560 12300
rect 8628 12244 8684 12300
rect 8752 12244 8808 12300
rect 8876 12244 8932 12300
rect 9000 12244 9056 12300
rect 9124 12244 9180 12300
rect 9248 12244 9304 12300
rect 9372 12244 9428 12300
rect 9496 12244 9552 12300
rect 9620 12244 9676 12300
rect 9744 12244 9800 12300
rect 7884 12120 7940 12176
rect 8008 12120 8064 12176
rect 8132 12120 8188 12176
rect 8256 12120 8312 12176
rect 8380 12120 8436 12176
rect 8504 12120 8560 12176
rect 8628 12120 8684 12176
rect 8752 12120 8808 12176
rect 8876 12120 8932 12176
rect 9000 12120 9056 12176
rect 9124 12120 9180 12176
rect 9248 12120 9304 12176
rect 9372 12120 9428 12176
rect 9496 12120 9552 12176
rect 9620 12120 9676 12176
rect 9744 12120 9800 12176
rect 7884 11996 7940 12052
rect 8008 11996 8064 12052
rect 8132 11996 8188 12052
rect 8256 11996 8312 12052
rect 8380 11996 8436 12052
rect 8504 11996 8560 12052
rect 8628 11996 8684 12052
rect 8752 11996 8808 12052
rect 8876 11996 8932 12052
rect 9000 11996 9056 12052
rect 9124 11996 9180 12052
rect 9248 11996 9304 12052
rect 9372 11996 9428 12052
rect 9496 11996 9552 12052
rect 9620 11996 9676 12052
rect 9744 11996 9800 12052
rect 7884 11872 7940 11928
rect 8008 11872 8064 11928
rect 8132 11872 8188 11928
rect 8256 11872 8312 11928
rect 8380 11872 8436 11928
rect 8504 11872 8560 11928
rect 8628 11872 8684 11928
rect 8752 11872 8808 11928
rect 8876 11872 8932 11928
rect 9000 11872 9056 11928
rect 9124 11872 9180 11928
rect 9248 11872 9304 11928
rect 9372 11872 9428 11928
rect 9496 11872 9552 11928
rect 9620 11872 9676 11928
rect 9744 11872 9800 11928
rect 7884 11748 7940 11804
rect 8008 11748 8064 11804
rect 8132 11748 8188 11804
rect 8256 11748 8312 11804
rect 8380 11748 8436 11804
rect 8504 11748 8560 11804
rect 8628 11748 8684 11804
rect 8752 11748 8808 11804
rect 8876 11748 8932 11804
rect 9000 11748 9056 11804
rect 9124 11748 9180 11804
rect 9248 11748 9304 11804
rect 9372 11748 9428 11804
rect 9496 11748 9552 11804
rect 9620 11748 9676 11804
rect 9744 11748 9800 11804
rect 7884 11624 7940 11680
rect 8008 11624 8064 11680
rect 8132 11624 8188 11680
rect 8256 11624 8312 11680
rect 8380 11624 8436 11680
rect 8504 11624 8560 11680
rect 8628 11624 8684 11680
rect 8752 11624 8808 11680
rect 8876 11624 8932 11680
rect 9000 11624 9056 11680
rect 9124 11624 9180 11680
rect 9248 11624 9304 11680
rect 9372 11624 9428 11680
rect 9496 11624 9552 11680
rect 9620 11624 9676 11680
rect 9744 11624 9800 11680
rect 7884 11500 7940 11556
rect 8008 11500 8064 11556
rect 8132 11500 8188 11556
rect 8256 11500 8312 11556
rect 8380 11500 8436 11556
rect 8504 11500 8560 11556
rect 8628 11500 8684 11556
rect 8752 11500 8808 11556
rect 8876 11500 8932 11556
rect 9000 11500 9056 11556
rect 9124 11500 9180 11556
rect 9248 11500 9304 11556
rect 9372 11500 9428 11556
rect 9496 11500 9552 11556
rect 9620 11500 9676 11556
rect 9744 11500 9800 11556
rect 7884 11376 7940 11432
rect 8008 11376 8064 11432
rect 8132 11376 8188 11432
rect 8256 11376 8312 11432
rect 8380 11376 8436 11432
rect 8504 11376 8560 11432
rect 8628 11376 8684 11432
rect 8752 11376 8808 11432
rect 8876 11376 8932 11432
rect 9000 11376 9056 11432
rect 9124 11376 9180 11432
rect 9248 11376 9304 11432
rect 9372 11376 9428 11432
rect 9496 11376 9552 11432
rect 9620 11376 9676 11432
rect 9744 11376 9800 11432
rect 7884 11252 7940 11308
rect 8008 11252 8064 11308
rect 8132 11252 8188 11308
rect 8256 11252 8312 11308
rect 8380 11252 8436 11308
rect 8504 11252 8560 11308
rect 8628 11252 8684 11308
rect 8752 11252 8808 11308
rect 8876 11252 8932 11308
rect 9000 11252 9056 11308
rect 9124 11252 9180 11308
rect 9248 11252 9304 11308
rect 9372 11252 9428 11308
rect 9496 11252 9552 11308
rect 9620 11252 9676 11308
rect 9744 11252 9800 11308
rect 10254 12492 10310 12548
rect 10378 12492 10434 12548
rect 10502 12492 10558 12548
rect 10626 12492 10682 12548
rect 10750 12492 10806 12548
rect 10874 12492 10930 12548
rect 10998 12492 11054 12548
rect 11122 12492 11178 12548
rect 11246 12492 11302 12548
rect 11370 12492 11426 12548
rect 11494 12492 11550 12548
rect 11618 12492 11674 12548
rect 11742 12492 11798 12548
rect 11866 12492 11922 12548
rect 11990 12492 12046 12548
rect 12114 12492 12170 12548
rect 10254 12368 10310 12424
rect 10378 12368 10434 12424
rect 10502 12368 10558 12424
rect 10626 12368 10682 12424
rect 10750 12368 10806 12424
rect 10874 12368 10930 12424
rect 10998 12368 11054 12424
rect 11122 12368 11178 12424
rect 11246 12368 11302 12424
rect 11370 12368 11426 12424
rect 11494 12368 11550 12424
rect 11618 12368 11674 12424
rect 11742 12368 11798 12424
rect 11866 12368 11922 12424
rect 11990 12368 12046 12424
rect 12114 12368 12170 12424
rect 10254 12244 10310 12300
rect 10378 12244 10434 12300
rect 10502 12244 10558 12300
rect 10626 12244 10682 12300
rect 10750 12244 10806 12300
rect 10874 12244 10930 12300
rect 10998 12244 11054 12300
rect 11122 12244 11178 12300
rect 11246 12244 11302 12300
rect 11370 12244 11426 12300
rect 11494 12244 11550 12300
rect 11618 12244 11674 12300
rect 11742 12244 11798 12300
rect 11866 12244 11922 12300
rect 11990 12244 12046 12300
rect 12114 12244 12170 12300
rect 10254 12120 10310 12176
rect 10378 12120 10434 12176
rect 10502 12120 10558 12176
rect 10626 12120 10682 12176
rect 10750 12120 10806 12176
rect 10874 12120 10930 12176
rect 10998 12120 11054 12176
rect 11122 12120 11178 12176
rect 11246 12120 11302 12176
rect 11370 12120 11426 12176
rect 11494 12120 11550 12176
rect 11618 12120 11674 12176
rect 11742 12120 11798 12176
rect 11866 12120 11922 12176
rect 11990 12120 12046 12176
rect 12114 12120 12170 12176
rect 10254 11996 10310 12052
rect 10378 11996 10434 12052
rect 10502 11996 10558 12052
rect 10626 11996 10682 12052
rect 10750 11996 10806 12052
rect 10874 11996 10930 12052
rect 10998 11996 11054 12052
rect 11122 11996 11178 12052
rect 11246 11996 11302 12052
rect 11370 11996 11426 12052
rect 11494 11996 11550 12052
rect 11618 11996 11674 12052
rect 11742 11996 11798 12052
rect 11866 11996 11922 12052
rect 11990 11996 12046 12052
rect 12114 11996 12170 12052
rect 10254 11872 10310 11928
rect 10378 11872 10434 11928
rect 10502 11872 10558 11928
rect 10626 11872 10682 11928
rect 10750 11872 10806 11928
rect 10874 11872 10930 11928
rect 10998 11872 11054 11928
rect 11122 11872 11178 11928
rect 11246 11872 11302 11928
rect 11370 11872 11426 11928
rect 11494 11872 11550 11928
rect 11618 11872 11674 11928
rect 11742 11872 11798 11928
rect 11866 11872 11922 11928
rect 11990 11872 12046 11928
rect 12114 11872 12170 11928
rect 10254 11748 10310 11804
rect 10378 11748 10434 11804
rect 10502 11748 10558 11804
rect 10626 11748 10682 11804
rect 10750 11748 10806 11804
rect 10874 11748 10930 11804
rect 10998 11748 11054 11804
rect 11122 11748 11178 11804
rect 11246 11748 11302 11804
rect 11370 11748 11426 11804
rect 11494 11748 11550 11804
rect 11618 11748 11674 11804
rect 11742 11748 11798 11804
rect 11866 11748 11922 11804
rect 11990 11748 12046 11804
rect 12114 11748 12170 11804
rect 10254 11624 10310 11680
rect 10378 11624 10434 11680
rect 10502 11624 10558 11680
rect 10626 11624 10682 11680
rect 10750 11624 10806 11680
rect 10874 11624 10930 11680
rect 10998 11624 11054 11680
rect 11122 11624 11178 11680
rect 11246 11624 11302 11680
rect 11370 11624 11426 11680
rect 11494 11624 11550 11680
rect 11618 11624 11674 11680
rect 11742 11624 11798 11680
rect 11866 11624 11922 11680
rect 11990 11624 12046 11680
rect 12114 11624 12170 11680
rect 10254 11500 10310 11556
rect 10378 11500 10434 11556
rect 10502 11500 10558 11556
rect 10626 11500 10682 11556
rect 10750 11500 10806 11556
rect 10874 11500 10930 11556
rect 10998 11500 11054 11556
rect 11122 11500 11178 11556
rect 11246 11500 11302 11556
rect 11370 11500 11426 11556
rect 11494 11500 11550 11556
rect 11618 11500 11674 11556
rect 11742 11500 11798 11556
rect 11866 11500 11922 11556
rect 11990 11500 12046 11556
rect 12114 11500 12170 11556
rect 10254 11376 10310 11432
rect 10378 11376 10434 11432
rect 10502 11376 10558 11432
rect 10626 11376 10682 11432
rect 10750 11376 10806 11432
rect 10874 11376 10930 11432
rect 10998 11376 11054 11432
rect 11122 11376 11178 11432
rect 11246 11376 11302 11432
rect 11370 11376 11426 11432
rect 11494 11376 11550 11432
rect 11618 11376 11674 11432
rect 11742 11376 11798 11432
rect 11866 11376 11922 11432
rect 11990 11376 12046 11432
rect 12114 11376 12170 11432
rect 10254 11252 10310 11308
rect 10378 11252 10434 11308
rect 10502 11252 10558 11308
rect 10626 11252 10682 11308
rect 10750 11252 10806 11308
rect 10874 11252 10930 11308
rect 10998 11252 11054 11308
rect 11122 11252 11178 11308
rect 11246 11252 11302 11308
rect 11370 11252 11426 11308
rect 11494 11252 11550 11308
rect 11618 11252 11674 11308
rect 11742 11252 11798 11308
rect 11866 11252 11922 11308
rect 11990 11252 12046 11308
rect 12114 11252 12170 11308
rect 12871 12492 12927 12548
rect 12995 12492 13051 12548
rect 13119 12492 13175 12548
rect 13243 12492 13299 12548
rect 13367 12492 13423 12548
rect 13491 12492 13547 12548
rect 13615 12492 13671 12548
rect 13739 12492 13795 12548
rect 13863 12492 13919 12548
rect 13987 12492 14043 12548
rect 14111 12492 14167 12548
rect 14235 12492 14291 12548
rect 14359 12492 14415 12548
rect 14483 12492 14539 12548
rect 14607 12492 14663 12548
rect 12871 12368 12927 12424
rect 12995 12368 13051 12424
rect 13119 12368 13175 12424
rect 13243 12368 13299 12424
rect 13367 12368 13423 12424
rect 13491 12368 13547 12424
rect 13615 12368 13671 12424
rect 13739 12368 13795 12424
rect 13863 12368 13919 12424
rect 13987 12368 14043 12424
rect 14111 12368 14167 12424
rect 14235 12368 14291 12424
rect 14359 12368 14415 12424
rect 14483 12368 14539 12424
rect 14607 12368 14663 12424
rect 12871 12244 12927 12300
rect 12995 12244 13051 12300
rect 13119 12244 13175 12300
rect 13243 12244 13299 12300
rect 13367 12244 13423 12300
rect 13491 12244 13547 12300
rect 13615 12244 13671 12300
rect 13739 12244 13795 12300
rect 13863 12244 13919 12300
rect 13987 12244 14043 12300
rect 14111 12244 14167 12300
rect 14235 12244 14291 12300
rect 14359 12244 14415 12300
rect 14483 12244 14539 12300
rect 14607 12244 14663 12300
rect 12871 12120 12927 12176
rect 12995 12120 13051 12176
rect 13119 12120 13175 12176
rect 13243 12120 13299 12176
rect 13367 12120 13423 12176
rect 13491 12120 13547 12176
rect 13615 12120 13671 12176
rect 13739 12120 13795 12176
rect 13863 12120 13919 12176
rect 13987 12120 14043 12176
rect 14111 12120 14167 12176
rect 14235 12120 14291 12176
rect 14359 12120 14415 12176
rect 14483 12120 14539 12176
rect 14607 12120 14663 12176
rect 12871 11996 12927 12052
rect 12995 11996 13051 12052
rect 13119 11996 13175 12052
rect 13243 11996 13299 12052
rect 13367 11996 13423 12052
rect 13491 11996 13547 12052
rect 13615 11996 13671 12052
rect 13739 11996 13795 12052
rect 13863 11996 13919 12052
rect 13987 11996 14043 12052
rect 14111 11996 14167 12052
rect 14235 11996 14291 12052
rect 14359 11996 14415 12052
rect 14483 11996 14539 12052
rect 14607 11996 14663 12052
rect 12871 11872 12927 11928
rect 12995 11872 13051 11928
rect 13119 11872 13175 11928
rect 13243 11872 13299 11928
rect 13367 11872 13423 11928
rect 13491 11872 13547 11928
rect 13615 11872 13671 11928
rect 13739 11872 13795 11928
rect 13863 11872 13919 11928
rect 13987 11872 14043 11928
rect 14111 11872 14167 11928
rect 14235 11872 14291 11928
rect 14359 11872 14415 11928
rect 14483 11872 14539 11928
rect 14607 11872 14663 11928
rect 12871 11748 12927 11804
rect 12995 11748 13051 11804
rect 13119 11748 13175 11804
rect 13243 11748 13299 11804
rect 13367 11748 13423 11804
rect 13491 11748 13547 11804
rect 13615 11748 13671 11804
rect 13739 11748 13795 11804
rect 13863 11748 13919 11804
rect 13987 11748 14043 11804
rect 14111 11748 14167 11804
rect 14235 11748 14291 11804
rect 14359 11748 14415 11804
rect 14483 11748 14539 11804
rect 14607 11748 14663 11804
rect 12871 11624 12927 11680
rect 12995 11624 13051 11680
rect 13119 11624 13175 11680
rect 13243 11624 13299 11680
rect 13367 11624 13423 11680
rect 13491 11624 13547 11680
rect 13615 11624 13671 11680
rect 13739 11624 13795 11680
rect 13863 11624 13919 11680
rect 13987 11624 14043 11680
rect 14111 11624 14167 11680
rect 14235 11624 14291 11680
rect 14359 11624 14415 11680
rect 14483 11624 14539 11680
rect 14607 11624 14663 11680
rect 12871 11500 12927 11556
rect 12995 11500 13051 11556
rect 13119 11500 13175 11556
rect 13243 11500 13299 11556
rect 13367 11500 13423 11556
rect 13491 11500 13547 11556
rect 13615 11500 13671 11556
rect 13739 11500 13795 11556
rect 13863 11500 13919 11556
rect 13987 11500 14043 11556
rect 14111 11500 14167 11556
rect 14235 11500 14291 11556
rect 14359 11500 14415 11556
rect 14483 11500 14539 11556
rect 14607 11500 14663 11556
rect 12871 11376 12927 11432
rect 12995 11376 13051 11432
rect 13119 11376 13175 11432
rect 13243 11376 13299 11432
rect 13367 11376 13423 11432
rect 13491 11376 13547 11432
rect 13615 11376 13671 11432
rect 13739 11376 13795 11432
rect 13863 11376 13919 11432
rect 13987 11376 14043 11432
rect 14111 11376 14167 11432
rect 14235 11376 14291 11432
rect 14359 11376 14415 11432
rect 14483 11376 14539 11432
rect 14607 11376 14663 11432
rect 12871 11252 12927 11308
rect 12995 11252 13051 11308
rect 13119 11252 13175 11308
rect 13243 11252 13299 11308
rect 13367 11252 13423 11308
rect 13491 11252 13547 11308
rect 13615 11252 13671 11308
rect 13739 11252 13795 11308
rect 13863 11252 13919 11308
rect 13987 11252 14043 11308
rect 14111 11252 14167 11308
rect 14235 11252 14291 11308
rect 14359 11252 14415 11308
rect 14483 11252 14539 11308
rect 14607 11252 14663 11308
rect 2491 10898 2547 10954
rect 2615 10898 2671 10954
rect 2491 10774 2547 10830
rect 2615 10774 2671 10830
rect 2491 10650 2547 10706
rect 2615 10650 2671 10706
rect 2491 10526 2547 10582
rect 2615 10526 2671 10582
rect 2491 10402 2547 10458
rect 2615 10402 2671 10458
rect 2491 10278 2547 10334
rect 2615 10278 2671 10334
rect 2491 10154 2547 10210
rect 2615 10154 2671 10210
rect 2491 10030 2547 10086
rect 2615 10030 2671 10086
rect 2491 9906 2547 9962
rect 2615 9906 2671 9962
rect 2491 9782 2547 9838
rect 2615 9782 2671 9838
rect 2491 9658 2547 9714
rect 2615 9658 2671 9714
rect 2491 9534 2547 9590
rect 2615 9534 2671 9590
rect 2491 9410 2547 9466
rect 2615 9410 2671 9466
rect 2491 9286 2547 9342
rect 2615 9286 2671 9342
rect 2491 9162 2547 9218
rect 2615 9162 2671 9218
rect 2491 9038 2547 9094
rect 2615 9038 2671 9094
rect 2491 8914 2547 8970
rect 2615 8914 2671 8970
rect 2491 8790 2547 8846
rect 2615 8790 2671 8846
rect 2491 8666 2547 8722
rect 2615 8666 2671 8722
rect 2491 8542 2547 8598
rect 2615 8542 2671 8598
rect 2491 8418 2547 8474
rect 2615 8418 2671 8474
rect 2491 8294 2547 8350
rect 2615 8294 2671 8350
rect 2491 8170 2547 8226
rect 2615 8170 2671 8226
rect 2491 8046 2547 8102
rect 2615 8046 2671 8102
rect 4861 10898 4917 10954
rect 4985 10898 5041 10954
rect 4861 10774 4917 10830
rect 4985 10774 5041 10830
rect 4861 10650 4917 10706
rect 4985 10650 5041 10706
rect 4861 10526 4917 10582
rect 4985 10526 5041 10582
rect 4861 10402 4917 10458
rect 4985 10402 5041 10458
rect 4861 10278 4917 10334
rect 4985 10278 5041 10334
rect 4861 10154 4917 10210
rect 4985 10154 5041 10210
rect 4861 10030 4917 10086
rect 4985 10030 5041 10086
rect 4861 9906 4917 9962
rect 4985 9906 5041 9962
rect 4861 9782 4917 9838
rect 4985 9782 5041 9838
rect 4861 9658 4917 9714
rect 4985 9658 5041 9714
rect 4861 9534 4917 9590
rect 4985 9534 5041 9590
rect 4861 9410 4917 9466
rect 4985 9410 5041 9466
rect 4861 9286 4917 9342
rect 4985 9286 5041 9342
rect 4861 9162 4917 9218
rect 4985 9162 5041 9218
rect 4861 9038 4917 9094
rect 4985 9038 5041 9094
rect 4861 8914 4917 8970
rect 4985 8914 5041 8970
rect 4861 8790 4917 8846
rect 4985 8790 5041 8846
rect 4861 8666 4917 8722
rect 4985 8666 5041 8722
rect 4861 8542 4917 8598
rect 4985 8542 5041 8598
rect 4861 8418 4917 8474
rect 4985 8418 5041 8474
rect 4861 8294 4917 8350
rect 4985 8294 5041 8350
rect 4861 8170 4917 8226
rect 4985 8170 5041 8226
rect 4861 8046 4917 8102
rect 4985 8046 5041 8102
rect 7275 10898 7331 10954
rect 7399 10898 7455 10954
rect 7523 10898 7579 10954
rect 7647 10898 7703 10954
rect 7275 10774 7331 10830
rect 7399 10774 7455 10830
rect 7523 10774 7579 10830
rect 7647 10774 7703 10830
rect 7275 10650 7331 10706
rect 7399 10650 7455 10706
rect 7523 10650 7579 10706
rect 7647 10650 7703 10706
rect 7275 10526 7331 10582
rect 7399 10526 7455 10582
rect 7523 10526 7579 10582
rect 7647 10526 7703 10582
rect 7275 10402 7331 10458
rect 7399 10402 7455 10458
rect 7523 10402 7579 10458
rect 7647 10402 7703 10458
rect 7275 10278 7331 10334
rect 7399 10278 7455 10334
rect 7523 10278 7579 10334
rect 7647 10278 7703 10334
rect 7275 10154 7331 10210
rect 7399 10154 7455 10210
rect 7523 10154 7579 10210
rect 7647 10154 7703 10210
rect 7275 10030 7331 10086
rect 7399 10030 7455 10086
rect 7523 10030 7579 10086
rect 7647 10030 7703 10086
rect 7275 9906 7331 9962
rect 7399 9906 7455 9962
rect 7523 9906 7579 9962
rect 7647 9906 7703 9962
rect 7275 9782 7331 9838
rect 7399 9782 7455 9838
rect 7523 9782 7579 9838
rect 7647 9782 7703 9838
rect 7275 9658 7331 9714
rect 7399 9658 7455 9714
rect 7523 9658 7579 9714
rect 7647 9658 7703 9714
rect 7275 9534 7331 9590
rect 7399 9534 7455 9590
rect 7523 9534 7579 9590
rect 7647 9534 7703 9590
rect 7275 9410 7331 9466
rect 7399 9410 7455 9466
rect 7523 9410 7579 9466
rect 7647 9410 7703 9466
rect 7275 9286 7331 9342
rect 7399 9286 7455 9342
rect 7523 9286 7579 9342
rect 7647 9286 7703 9342
rect 7275 9162 7331 9218
rect 7399 9162 7455 9218
rect 7523 9162 7579 9218
rect 7647 9162 7703 9218
rect 7275 9038 7331 9094
rect 7399 9038 7455 9094
rect 7523 9038 7579 9094
rect 7647 9038 7703 9094
rect 7275 8914 7331 8970
rect 7399 8914 7455 8970
rect 7523 8914 7579 8970
rect 7647 8914 7703 8970
rect 7275 8790 7331 8846
rect 7399 8790 7455 8846
rect 7523 8790 7579 8846
rect 7647 8790 7703 8846
rect 7275 8666 7331 8722
rect 7399 8666 7455 8722
rect 7523 8666 7579 8722
rect 7647 8666 7703 8722
rect 7275 8542 7331 8598
rect 7399 8542 7455 8598
rect 7523 8542 7579 8598
rect 7647 8542 7703 8598
rect 7275 8418 7331 8474
rect 7399 8418 7455 8474
rect 7523 8418 7579 8474
rect 7647 8418 7703 8474
rect 7275 8294 7331 8350
rect 7399 8294 7455 8350
rect 7523 8294 7579 8350
rect 7647 8294 7703 8350
rect 7275 8170 7331 8226
rect 7399 8170 7455 8226
rect 7523 8170 7579 8226
rect 7647 8170 7703 8226
rect 7275 8046 7331 8102
rect 7399 8046 7455 8102
rect 7523 8046 7579 8102
rect 7647 8046 7703 8102
rect 9937 10898 9993 10954
rect 10061 10898 10117 10954
rect 9937 10774 9993 10830
rect 10061 10774 10117 10830
rect 9937 10650 9993 10706
rect 10061 10650 10117 10706
rect 9937 10526 9993 10582
rect 10061 10526 10117 10582
rect 9937 10402 9993 10458
rect 10061 10402 10117 10458
rect 9937 10278 9993 10334
rect 10061 10278 10117 10334
rect 9937 10154 9993 10210
rect 10061 10154 10117 10210
rect 9937 10030 9993 10086
rect 10061 10030 10117 10086
rect 9937 9906 9993 9962
rect 10061 9906 10117 9962
rect 9937 9782 9993 9838
rect 10061 9782 10117 9838
rect 9937 9658 9993 9714
rect 10061 9658 10117 9714
rect 9937 9534 9993 9590
rect 10061 9534 10117 9590
rect 9937 9410 9993 9466
rect 10061 9410 10117 9466
rect 9937 9286 9993 9342
rect 10061 9286 10117 9342
rect 9937 9162 9993 9218
rect 10061 9162 10117 9218
rect 9937 9038 9993 9094
rect 10061 9038 10117 9094
rect 9937 8914 9993 8970
rect 10061 8914 10117 8970
rect 9937 8790 9993 8846
rect 10061 8790 10117 8846
rect 9937 8666 9993 8722
rect 10061 8666 10117 8722
rect 9937 8542 9993 8598
rect 10061 8542 10117 8598
rect 9937 8418 9993 8474
rect 10061 8418 10117 8474
rect 9937 8294 9993 8350
rect 10061 8294 10117 8350
rect 9937 8170 9993 8226
rect 10061 8170 10117 8226
rect 9937 8046 9993 8102
rect 10061 8046 10117 8102
rect 12307 10898 12363 10954
rect 12431 10898 12487 10954
rect 12307 10774 12363 10830
rect 12431 10774 12487 10830
rect 12307 10650 12363 10706
rect 12431 10650 12487 10706
rect 12307 10526 12363 10582
rect 12431 10526 12487 10582
rect 12307 10402 12363 10458
rect 12431 10402 12487 10458
rect 12307 10278 12363 10334
rect 12431 10278 12487 10334
rect 12307 10154 12363 10210
rect 12431 10154 12487 10210
rect 12307 10030 12363 10086
rect 12431 10030 12487 10086
rect 12307 9906 12363 9962
rect 12431 9906 12487 9962
rect 12307 9782 12363 9838
rect 12431 9782 12487 9838
rect 12307 9658 12363 9714
rect 12431 9658 12487 9714
rect 12307 9534 12363 9590
rect 12431 9534 12487 9590
rect 12307 9410 12363 9466
rect 12431 9410 12487 9466
rect 12307 9286 12363 9342
rect 12431 9286 12487 9342
rect 12307 9162 12363 9218
rect 12431 9162 12487 9218
rect 12307 9038 12363 9094
rect 12431 9038 12487 9094
rect 12307 8914 12363 8970
rect 12431 8914 12487 8970
rect 12307 8790 12363 8846
rect 12431 8790 12487 8846
rect 12307 8666 12363 8722
rect 12431 8666 12487 8722
rect 12307 8542 12363 8598
rect 12431 8542 12487 8598
rect 12307 8418 12363 8474
rect 12431 8418 12487 8474
rect 12307 8294 12363 8350
rect 12431 8294 12487 8350
rect 12307 8170 12363 8226
rect 12431 8170 12487 8226
rect 12307 8046 12363 8102
rect 12431 8046 12487 8102
rect 2491 7698 2547 7754
rect 2615 7698 2671 7754
rect 2491 7574 2547 7630
rect 2615 7574 2671 7630
rect 2491 7450 2547 7506
rect 2615 7450 2671 7506
rect 2491 7326 2547 7382
rect 2615 7326 2671 7382
rect 2491 7202 2547 7258
rect 2615 7202 2671 7258
rect 2491 7078 2547 7134
rect 2615 7078 2671 7134
rect 2491 6954 2547 7010
rect 2615 6954 2671 7010
rect 2491 6830 2547 6886
rect 2615 6830 2671 6886
rect 2491 6706 2547 6762
rect 2615 6706 2671 6762
rect 2491 6582 2547 6638
rect 2615 6582 2671 6638
rect 2491 6458 2547 6514
rect 2615 6458 2671 6514
rect 2491 6334 2547 6390
rect 2615 6334 2671 6390
rect 2491 6210 2547 6266
rect 2615 6210 2671 6266
rect 2491 6086 2547 6142
rect 2615 6086 2671 6142
rect 2491 5962 2547 6018
rect 2615 5962 2671 6018
rect 2491 5838 2547 5894
rect 2615 5838 2671 5894
rect 2491 5714 2547 5770
rect 2615 5714 2671 5770
rect 2491 5590 2547 5646
rect 2615 5590 2671 5646
rect 2491 5466 2547 5522
rect 2615 5466 2671 5522
rect 2491 5342 2547 5398
rect 2615 5342 2671 5398
rect 2491 5218 2547 5274
rect 2615 5218 2671 5274
rect 2491 5094 2547 5150
rect 2615 5094 2671 5150
rect 2491 4970 2547 5026
rect 2615 4970 2671 5026
rect 2491 4846 2547 4902
rect 2615 4846 2671 4902
rect 4861 7698 4917 7754
rect 4985 7698 5041 7754
rect 4861 7574 4917 7630
rect 4985 7574 5041 7630
rect 4861 7450 4917 7506
rect 4985 7450 5041 7506
rect 4861 7326 4917 7382
rect 4985 7326 5041 7382
rect 4861 7202 4917 7258
rect 4985 7202 5041 7258
rect 4861 7078 4917 7134
rect 4985 7078 5041 7134
rect 4861 6954 4917 7010
rect 4985 6954 5041 7010
rect 4861 6830 4917 6886
rect 4985 6830 5041 6886
rect 4861 6706 4917 6762
rect 4985 6706 5041 6762
rect 4861 6582 4917 6638
rect 4985 6582 5041 6638
rect 4861 6458 4917 6514
rect 4985 6458 5041 6514
rect 4861 6334 4917 6390
rect 4985 6334 5041 6390
rect 4861 6210 4917 6266
rect 4985 6210 5041 6266
rect 4861 6086 4917 6142
rect 4985 6086 5041 6142
rect 4861 5962 4917 6018
rect 4985 5962 5041 6018
rect 4861 5838 4917 5894
rect 4985 5838 5041 5894
rect 4861 5714 4917 5770
rect 4985 5714 5041 5770
rect 4861 5590 4917 5646
rect 4985 5590 5041 5646
rect 4861 5466 4917 5522
rect 4985 5466 5041 5522
rect 4861 5342 4917 5398
rect 4985 5342 5041 5398
rect 4861 5218 4917 5274
rect 4985 5218 5041 5274
rect 4861 5094 4917 5150
rect 4985 5094 5041 5150
rect 4861 4970 4917 5026
rect 4985 4970 5041 5026
rect 4861 4846 4917 4902
rect 4985 4846 5041 4902
rect 7275 7698 7331 7754
rect 7399 7698 7455 7754
rect 7523 7698 7579 7754
rect 7647 7698 7703 7754
rect 7275 7574 7331 7630
rect 7399 7574 7455 7630
rect 7523 7574 7579 7630
rect 7647 7574 7703 7630
rect 7275 7450 7331 7506
rect 7399 7450 7455 7506
rect 7523 7450 7579 7506
rect 7647 7450 7703 7506
rect 7275 7326 7331 7382
rect 7399 7326 7455 7382
rect 7523 7326 7579 7382
rect 7647 7326 7703 7382
rect 7275 7202 7331 7258
rect 7399 7202 7455 7258
rect 7523 7202 7579 7258
rect 7647 7202 7703 7258
rect 7275 7078 7331 7134
rect 7399 7078 7455 7134
rect 7523 7078 7579 7134
rect 7647 7078 7703 7134
rect 7275 6954 7331 7010
rect 7399 6954 7455 7010
rect 7523 6954 7579 7010
rect 7647 6954 7703 7010
rect 7275 6830 7331 6886
rect 7399 6830 7455 6886
rect 7523 6830 7579 6886
rect 7647 6830 7703 6886
rect 7275 6706 7331 6762
rect 7399 6706 7455 6762
rect 7523 6706 7579 6762
rect 7647 6706 7703 6762
rect 7275 6582 7331 6638
rect 7399 6582 7455 6638
rect 7523 6582 7579 6638
rect 7647 6582 7703 6638
rect 7275 6458 7331 6514
rect 7399 6458 7455 6514
rect 7523 6458 7579 6514
rect 7647 6458 7703 6514
rect 7275 6334 7331 6390
rect 7399 6334 7455 6390
rect 7523 6334 7579 6390
rect 7647 6334 7703 6390
rect 7275 6210 7331 6266
rect 7399 6210 7455 6266
rect 7523 6210 7579 6266
rect 7647 6210 7703 6266
rect 7275 6086 7331 6142
rect 7399 6086 7455 6142
rect 7523 6086 7579 6142
rect 7647 6086 7703 6142
rect 7275 5962 7331 6018
rect 7399 5962 7455 6018
rect 7523 5962 7579 6018
rect 7647 5962 7703 6018
rect 7275 5838 7331 5894
rect 7399 5838 7455 5894
rect 7523 5838 7579 5894
rect 7647 5838 7703 5894
rect 7275 5714 7331 5770
rect 7399 5714 7455 5770
rect 7523 5714 7579 5770
rect 7647 5714 7703 5770
rect 7275 5590 7331 5646
rect 7399 5590 7455 5646
rect 7523 5590 7579 5646
rect 7647 5590 7703 5646
rect 7275 5466 7331 5522
rect 7399 5466 7455 5522
rect 7523 5466 7579 5522
rect 7647 5466 7703 5522
rect 7275 5342 7331 5398
rect 7399 5342 7455 5398
rect 7523 5342 7579 5398
rect 7647 5342 7703 5398
rect 7275 5218 7331 5274
rect 7399 5218 7455 5274
rect 7523 5218 7579 5274
rect 7647 5218 7703 5274
rect 7275 5094 7331 5150
rect 7399 5094 7455 5150
rect 7523 5094 7579 5150
rect 7647 5094 7703 5150
rect 7275 4970 7331 5026
rect 7399 4970 7455 5026
rect 7523 4970 7579 5026
rect 7647 4970 7703 5026
rect 7275 4846 7331 4902
rect 7399 4846 7455 4902
rect 7523 4846 7579 4902
rect 7647 4846 7703 4902
rect 9937 7698 9993 7754
rect 10061 7698 10117 7754
rect 9937 7574 9993 7630
rect 10061 7574 10117 7630
rect 9937 7450 9993 7506
rect 10061 7450 10117 7506
rect 9937 7326 9993 7382
rect 10061 7326 10117 7382
rect 9937 7202 9993 7258
rect 10061 7202 10117 7258
rect 9937 7078 9993 7134
rect 10061 7078 10117 7134
rect 9937 6954 9993 7010
rect 10061 6954 10117 7010
rect 9937 6830 9993 6886
rect 10061 6830 10117 6886
rect 9937 6706 9993 6762
rect 10061 6706 10117 6762
rect 9937 6582 9993 6638
rect 10061 6582 10117 6638
rect 9937 6458 9993 6514
rect 10061 6458 10117 6514
rect 9937 6334 9993 6390
rect 10061 6334 10117 6390
rect 9937 6210 9993 6266
rect 10061 6210 10117 6266
rect 9937 6086 9993 6142
rect 10061 6086 10117 6142
rect 9937 5962 9993 6018
rect 10061 5962 10117 6018
rect 9937 5838 9993 5894
rect 10061 5838 10117 5894
rect 9937 5714 9993 5770
rect 10061 5714 10117 5770
rect 9937 5590 9993 5646
rect 10061 5590 10117 5646
rect 9937 5466 9993 5522
rect 10061 5466 10117 5522
rect 9937 5342 9993 5398
rect 10061 5342 10117 5398
rect 9937 5218 9993 5274
rect 10061 5218 10117 5274
rect 9937 5094 9993 5150
rect 10061 5094 10117 5150
rect 9937 4970 9993 5026
rect 10061 4970 10117 5026
rect 9937 4846 9993 4902
rect 10061 4846 10117 4902
rect 12307 7698 12363 7754
rect 12431 7698 12487 7754
rect 12307 7574 12363 7630
rect 12431 7574 12487 7630
rect 12307 7450 12363 7506
rect 12431 7450 12487 7506
rect 12307 7326 12363 7382
rect 12431 7326 12487 7382
rect 12307 7202 12363 7258
rect 12431 7202 12487 7258
rect 12307 7078 12363 7134
rect 12431 7078 12487 7134
rect 12307 6954 12363 7010
rect 12431 6954 12487 7010
rect 12307 6830 12363 6886
rect 12431 6830 12487 6886
rect 12307 6706 12363 6762
rect 12431 6706 12487 6762
rect 12307 6582 12363 6638
rect 12431 6582 12487 6638
rect 12307 6458 12363 6514
rect 12431 6458 12487 6514
rect 12307 6334 12363 6390
rect 12431 6334 12487 6390
rect 12307 6210 12363 6266
rect 12431 6210 12487 6266
rect 12307 6086 12363 6142
rect 12431 6086 12487 6142
rect 12307 5962 12363 6018
rect 12431 5962 12487 6018
rect 12307 5838 12363 5894
rect 12431 5838 12487 5894
rect 12307 5714 12363 5770
rect 12431 5714 12487 5770
rect 12307 5590 12363 5646
rect 12431 5590 12487 5646
rect 12307 5466 12363 5522
rect 12431 5466 12487 5522
rect 12307 5342 12363 5398
rect 12431 5342 12487 5398
rect 12307 5218 12363 5274
rect 12431 5218 12487 5274
rect 12307 5094 12363 5150
rect 12431 5094 12487 5150
rect 12307 4970 12363 5026
rect 12431 4970 12487 5026
rect 12307 4846 12363 4902
rect 12431 4846 12487 4902
rect 2491 4498 2547 4554
rect 2615 4498 2671 4554
rect 2491 4374 2547 4430
rect 2615 4374 2671 4430
rect 2491 4250 2547 4306
rect 2615 4250 2671 4306
rect 2491 4126 2547 4182
rect 2615 4126 2671 4182
rect 2491 4002 2547 4058
rect 2615 4002 2671 4058
rect 2491 3878 2547 3934
rect 2615 3878 2671 3934
rect 2491 3754 2547 3810
rect 2615 3754 2671 3810
rect 2491 3630 2547 3686
rect 2615 3630 2671 3686
rect 2491 3506 2547 3562
rect 2615 3506 2671 3562
rect 2491 3382 2547 3438
rect 2615 3382 2671 3438
rect 2491 3258 2547 3314
rect 2615 3258 2671 3314
rect 2491 3134 2547 3190
rect 2615 3134 2671 3190
rect 2491 3010 2547 3066
rect 2615 3010 2671 3066
rect 2491 2886 2547 2942
rect 2615 2886 2671 2942
rect 2491 2762 2547 2818
rect 2615 2762 2671 2818
rect 2491 2638 2547 2694
rect 2615 2638 2671 2694
rect 2491 2514 2547 2570
rect 2615 2514 2671 2570
rect 2491 2390 2547 2446
rect 2615 2390 2671 2446
rect 2491 2266 2547 2322
rect 2615 2266 2671 2322
rect 2491 2142 2547 2198
rect 2615 2142 2671 2198
rect 2491 2018 2547 2074
rect 2615 2018 2671 2074
rect 2491 1894 2547 1950
rect 2615 1894 2671 1950
rect 2491 1770 2547 1826
rect 2615 1770 2671 1826
rect 2491 1646 2547 1702
rect 2615 1646 2671 1702
rect 4861 4498 4917 4554
rect 4985 4498 5041 4554
rect 4861 4374 4917 4430
rect 4985 4374 5041 4430
rect 4861 4250 4917 4306
rect 4985 4250 5041 4306
rect 4861 4126 4917 4182
rect 4985 4126 5041 4182
rect 4861 4002 4917 4058
rect 4985 4002 5041 4058
rect 4861 3878 4917 3934
rect 4985 3878 5041 3934
rect 4861 3754 4917 3810
rect 4985 3754 5041 3810
rect 4861 3630 4917 3686
rect 4985 3630 5041 3686
rect 4861 3506 4917 3562
rect 4985 3506 5041 3562
rect 4861 3382 4917 3438
rect 4985 3382 5041 3438
rect 4861 3258 4917 3314
rect 4985 3258 5041 3314
rect 4861 3134 4917 3190
rect 4985 3134 5041 3190
rect 4861 3010 4917 3066
rect 4985 3010 5041 3066
rect 4861 2886 4917 2942
rect 4985 2886 5041 2942
rect 4861 2762 4917 2818
rect 4985 2762 5041 2818
rect 4861 2638 4917 2694
rect 4985 2638 5041 2694
rect 4861 2514 4917 2570
rect 4985 2514 5041 2570
rect 4861 2390 4917 2446
rect 4985 2390 5041 2446
rect 4861 2266 4917 2322
rect 4985 2266 5041 2322
rect 4861 2142 4917 2198
rect 4985 2142 5041 2198
rect 4861 2018 4917 2074
rect 4985 2018 5041 2074
rect 4861 1894 4917 1950
rect 4985 1894 5041 1950
rect 4861 1770 4917 1826
rect 4985 1770 5041 1826
rect 4861 1646 4917 1702
rect 4985 1646 5041 1702
rect 7275 4498 7331 4554
rect 7399 4498 7455 4554
rect 7523 4498 7579 4554
rect 7647 4498 7703 4554
rect 7275 4374 7331 4430
rect 7399 4374 7455 4430
rect 7523 4374 7579 4430
rect 7647 4374 7703 4430
rect 7275 4250 7331 4306
rect 7399 4250 7455 4306
rect 7523 4250 7579 4306
rect 7647 4250 7703 4306
rect 7275 4126 7331 4182
rect 7399 4126 7455 4182
rect 7523 4126 7579 4182
rect 7647 4126 7703 4182
rect 7275 4002 7331 4058
rect 7399 4002 7455 4058
rect 7523 4002 7579 4058
rect 7647 4002 7703 4058
rect 7275 3878 7331 3934
rect 7399 3878 7455 3934
rect 7523 3878 7579 3934
rect 7647 3878 7703 3934
rect 7275 3754 7331 3810
rect 7399 3754 7455 3810
rect 7523 3754 7579 3810
rect 7647 3754 7703 3810
rect 7275 3630 7331 3686
rect 7399 3630 7455 3686
rect 7523 3630 7579 3686
rect 7647 3630 7703 3686
rect 7275 3506 7331 3562
rect 7399 3506 7455 3562
rect 7523 3506 7579 3562
rect 7647 3506 7703 3562
rect 7275 3382 7331 3438
rect 7399 3382 7455 3438
rect 7523 3382 7579 3438
rect 7647 3382 7703 3438
rect 7275 3258 7331 3314
rect 7399 3258 7455 3314
rect 7523 3258 7579 3314
rect 7647 3258 7703 3314
rect 7275 3134 7331 3190
rect 7399 3134 7455 3190
rect 7523 3134 7579 3190
rect 7647 3134 7703 3190
rect 7275 3010 7331 3066
rect 7399 3010 7455 3066
rect 7523 3010 7579 3066
rect 7647 3010 7703 3066
rect 7275 2886 7331 2942
rect 7399 2886 7455 2942
rect 7523 2886 7579 2942
rect 7647 2886 7703 2942
rect 7275 2762 7331 2818
rect 7399 2762 7455 2818
rect 7523 2762 7579 2818
rect 7647 2762 7703 2818
rect 7275 2638 7331 2694
rect 7399 2638 7455 2694
rect 7523 2638 7579 2694
rect 7647 2638 7703 2694
rect 7275 2514 7331 2570
rect 7399 2514 7455 2570
rect 7523 2514 7579 2570
rect 7647 2514 7703 2570
rect 7275 2390 7331 2446
rect 7399 2390 7455 2446
rect 7523 2390 7579 2446
rect 7647 2390 7703 2446
rect 7275 2266 7331 2322
rect 7399 2266 7455 2322
rect 7523 2266 7579 2322
rect 7647 2266 7703 2322
rect 7275 2142 7331 2198
rect 7399 2142 7455 2198
rect 7523 2142 7579 2198
rect 7647 2142 7703 2198
rect 7275 2018 7331 2074
rect 7399 2018 7455 2074
rect 7523 2018 7579 2074
rect 7647 2018 7703 2074
rect 7275 1894 7331 1950
rect 7399 1894 7455 1950
rect 7523 1894 7579 1950
rect 7647 1894 7703 1950
rect 7275 1770 7331 1826
rect 7399 1770 7455 1826
rect 7523 1770 7579 1826
rect 7647 1770 7703 1826
rect 7275 1646 7331 1702
rect 7399 1646 7455 1702
rect 7523 1646 7579 1702
rect 7647 1646 7703 1702
rect 9937 4498 9993 4554
rect 10061 4498 10117 4554
rect 9937 4374 9993 4430
rect 10061 4374 10117 4430
rect 9937 4250 9993 4306
rect 10061 4250 10117 4306
rect 9937 4126 9993 4182
rect 10061 4126 10117 4182
rect 9937 4002 9993 4058
rect 10061 4002 10117 4058
rect 9937 3878 9993 3934
rect 10061 3878 10117 3934
rect 9937 3754 9993 3810
rect 10061 3754 10117 3810
rect 9937 3630 9993 3686
rect 10061 3630 10117 3686
rect 9937 3506 9993 3562
rect 10061 3506 10117 3562
rect 9937 3382 9993 3438
rect 10061 3382 10117 3438
rect 9937 3258 9993 3314
rect 10061 3258 10117 3314
rect 9937 3134 9993 3190
rect 10061 3134 10117 3190
rect 9937 3010 9993 3066
rect 10061 3010 10117 3066
rect 9937 2886 9993 2942
rect 10061 2886 10117 2942
rect 9937 2762 9993 2818
rect 10061 2762 10117 2818
rect 9937 2638 9993 2694
rect 10061 2638 10117 2694
rect 9937 2514 9993 2570
rect 10061 2514 10117 2570
rect 9937 2390 9993 2446
rect 10061 2390 10117 2446
rect 9937 2266 9993 2322
rect 10061 2266 10117 2322
rect 9937 2142 9993 2198
rect 10061 2142 10117 2198
rect 9937 2018 9993 2074
rect 10061 2018 10117 2074
rect 9937 1894 9993 1950
rect 10061 1894 10117 1950
rect 9937 1770 9993 1826
rect 10061 1770 10117 1826
rect 9937 1646 9993 1702
rect 10061 1646 10117 1702
rect 12307 4498 12363 4554
rect 12431 4498 12487 4554
rect 12307 4374 12363 4430
rect 12431 4374 12487 4430
rect 12307 4250 12363 4306
rect 12431 4250 12487 4306
rect 12307 4126 12363 4182
rect 12431 4126 12487 4182
rect 12307 4002 12363 4058
rect 12431 4002 12487 4058
rect 12307 3878 12363 3934
rect 12431 3878 12487 3934
rect 12307 3754 12363 3810
rect 12431 3754 12487 3810
rect 12307 3630 12363 3686
rect 12431 3630 12487 3686
rect 12307 3506 12363 3562
rect 12431 3506 12487 3562
rect 12307 3382 12363 3438
rect 12431 3382 12487 3438
rect 12307 3258 12363 3314
rect 12431 3258 12487 3314
rect 12307 3134 12363 3190
rect 12431 3134 12487 3190
rect 12307 3010 12363 3066
rect 12431 3010 12487 3066
rect 12307 2886 12363 2942
rect 12431 2886 12487 2942
rect 12307 2762 12363 2818
rect 12431 2762 12487 2818
rect 12307 2638 12363 2694
rect 12431 2638 12487 2694
rect 12307 2514 12363 2570
rect 12431 2514 12487 2570
rect 12307 2390 12363 2446
rect 12431 2390 12487 2446
rect 12307 2266 12363 2322
rect 12431 2266 12487 2322
rect 12307 2142 12363 2198
rect 12431 2142 12487 2198
rect 12307 2018 12363 2074
rect 12431 2018 12487 2074
rect 12307 1894 12363 1950
rect 12431 1894 12487 1950
rect 12307 1770 12363 1826
rect 12431 1770 12487 1826
rect 12307 1646 12363 1702
rect 12431 1646 12487 1702
<< metal3 >>
rect 2481 57225 2681 57235
rect 2481 57169 2491 57225
rect 2547 57169 2615 57225
rect 2671 57169 2681 57225
rect 2481 57101 2681 57169
rect 2481 57045 2491 57101
rect 2547 57045 2615 57101
rect 2671 57045 2681 57101
rect 2481 56977 2681 57045
rect 2481 56921 2491 56977
rect 2547 56921 2615 56977
rect 2671 56921 2681 56977
rect 2481 56853 2681 56921
rect 2481 56797 2491 56853
rect 2547 56797 2615 56853
rect 2671 56797 2681 56853
rect 2481 56729 2681 56797
rect 2481 56673 2491 56729
rect 2547 56673 2615 56729
rect 2671 56673 2681 56729
rect 2481 56605 2681 56673
rect 2481 56549 2491 56605
rect 2547 56549 2615 56605
rect 2671 56549 2681 56605
rect 2481 56481 2681 56549
rect 2481 56425 2491 56481
rect 2547 56425 2615 56481
rect 2671 56425 2681 56481
rect 2481 56357 2681 56425
rect 2481 56301 2491 56357
rect 2547 56301 2615 56357
rect 2671 56301 2681 56357
rect 2481 56233 2681 56301
rect 2481 56177 2491 56233
rect 2547 56177 2615 56233
rect 2671 56177 2681 56233
rect 2481 56109 2681 56177
rect 2481 56053 2491 56109
rect 2547 56053 2615 56109
rect 2671 56053 2681 56109
rect 2481 56043 2681 56053
rect 4851 57225 5051 57235
rect 4851 57169 4861 57225
rect 4917 57169 4985 57225
rect 5041 57169 5051 57225
rect 4851 57101 5051 57169
rect 4851 57045 4861 57101
rect 4917 57045 4985 57101
rect 5041 57045 5051 57101
rect 4851 56977 5051 57045
rect 4851 56921 4861 56977
rect 4917 56921 4985 56977
rect 5041 56921 5051 56977
rect 4851 56853 5051 56921
rect 4851 56797 4861 56853
rect 4917 56797 4985 56853
rect 5041 56797 5051 56853
rect 4851 56729 5051 56797
rect 4851 56673 4861 56729
rect 4917 56673 4985 56729
rect 5041 56673 5051 56729
rect 4851 56605 5051 56673
rect 4851 56549 4861 56605
rect 4917 56549 4985 56605
rect 5041 56549 5051 56605
rect 4851 56481 5051 56549
rect 4851 56425 4861 56481
rect 4917 56425 4985 56481
rect 5041 56425 5051 56481
rect 4851 56357 5051 56425
rect 4851 56301 4861 56357
rect 4917 56301 4985 56357
rect 5041 56301 5051 56357
rect 4851 56233 5051 56301
rect 4851 56177 4861 56233
rect 4917 56177 4985 56233
rect 5041 56177 5051 56233
rect 4851 56109 5051 56177
rect 4851 56053 4861 56109
rect 4917 56053 4985 56109
rect 5041 56053 5051 56109
rect 4851 56043 5051 56053
rect 7265 57225 7713 57235
rect 7265 57169 7275 57225
rect 7331 57169 7399 57225
rect 7455 57169 7523 57225
rect 7579 57169 7647 57225
rect 7703 57169 7713 57225
rect 7265 57101 7713 57169
rect 7265 57045 7275 57101
rect 7331 57045 7399 57101
rect 7455 57045 7523 57101
rect 7579 57045 7647 57101
rect 7703 57045 7713 57101
rect 7265 56977 7713 57045
rect 7265 56921 7275 56977
rect 7331 56921 7399 56977
rect 7455 56921 7523 56977
rect 7579 56921 7647 56977
rect 7703 56921 7713 56977
rect 7265 56853 7713 56921
rect 7265 56797 7275 56853
rect 7331 56797 7399 56853
rect 7455 56797 7523 56853
rect 7579 56797 7647 56853
rect 7703 56797 7713 56853
rect 7265 56729 7713 56797
rect 7265 56673 7275 56729
rect 7331 56673 7399 56729
rect 7455 56673 7523 56729
rect 7579 56673 7647 56729
rect 7703 56673 7713 56729
rect 7265 56605 7713 56673
rect 7265 56549 7275 56605
rect 7331 56549 7399 56605
rect 7455 56549 7523 56605
rect 7579 56549 7647 56605
rect 7703 56549 7713 56605
rect 7265 56481 7713 56549
rect 7265 56425 7275 56481
rect 7331 56425 7399 56481
rect 7455 56425 7523 56481
rect 7579 56425 7647 56481
rect 7703 56425 7713 56481
rect 7265 56357 7713 56425
rect 7265 56301 7275 56357
rect 7331 56301 7399 56357
rect 7455 56301 7523 56357
rect 7579 56301 7647 56357
rect 7703 56301 7713 56357
rect 7265 56233 7713 56301
rect 7265 56177 7275 56233
rect 7331 56177 7399 56233
rect 7455 56177 7523 56233
rect 7579 56177 7647 56233
rect 7703 56177 7713 56233
rect 7265 56109 7713 56177
rect 7265 56053 7275 56109
rect 7331 56053 7399 56109
rect 7455 56053 7523 56109
rect 7579 56053 7647 56109
rect 7703 56053 7713 56109
rect 7265 56043 7713 56053
rect 9927 57225 10127 57235
rect 9927 57169 9937 57225
rect 9993 57169 10061 57225
rect 10117 57169 10127 57225
rect 9927 57101 10127 57169
rect 9927 57045 9937 57101
rect 9993 57045 10061 57101
rect 10117 57045 10127 57101
rect 9927 56977 10127 57045
rect 9927 56921 9937 56977
rect 9993 56921 10061 56977
rect 10117 56921 10127 56977
rect 9927 56853 10127 56921
rect 9927 56797 9937 56853
rect 9993 56797 10061 56853
rect 10117 56797 10127 56853
rect 9927 56729 10127 56797
rect 9927 56673 9937 56729
rect 9993 56673 10061 56729
rect 10117 56673 10127 56729
rect 9927 56605 10127 56673
rect 9927 56549 9937 56605
rect 9993 56549 10061 56605
rect 10117 56549 10127 56605
rect 9927 56481 10127 56549
rect 9927 56425 9937 56481
rect 9993 56425 10061 56481
rect 10117 56425 10127 56481
rect 9927 56357 10127 56425
rect 9927 56301 9937 56357
rect 9993 56301 10061 56357
rect 10117 56301 10127 56357
rect 9927 56233 10127 56301
rect 9927 56177 9937 56233
rect 9993 56177 10061 56233
rect 10117 56177 10127 56233
rect 9927 56109 10127 56177
rect 9927 56053 9937 56109
rect 9993 56053 10061 56109
rect 10117 56053 10127 56109
rect 9927 56043 10127 56053
rect 12297 57225 12497 57235
rect 12297 57169 12307 57225
rect 12363 57169 12431 57225
rect 12487 57169 12497 57225
rect 12297 57101 12497 57169
rect 12297 57045 12307 57101
rect 12363 57045 12431 57101
rect 12487 57045 12497 57101
rect 12297 56977 12497 57045
rect 12297 56921 12307 56977
rect 12363 56921 12431 56977
rect 12487 56921 12497 56977
rect 12297 56853 12497 56921
rect 12297 56797 12307 56853
rect 12363 56797 12431 56853
rect 12487 56797 12497 56853
rect 12297 56729 12497 56797
rect 12297 56673 12307 56729
rect 12363 56673 12431 56729
rect 12487 56673 12497 56729
rect 12297 56605 12497 56673
rect 12297 56549 12307 56605
rect 12363 56549 12431 56605
rect 12487 56549 12497 56605
rect 12297 56481 12497 56549
rect 12297 56425 12307 56481
rect 12363 56425 12431 56481
rect 12487 56425 12497 56481
rect 12297 56357 12497 56425
rect 12297 56301 12307 56357
rect 12363 56301 12431 56357
rect 12487 56301 12497 56357
rect 12297 56233 12497 56301
rect 12297 56177 12307 56233
rect 12363 56177 12431 56233
rect 12487 56177 12497 56233
rect 12297 56109 12497 56177
rect 12297 56053 12307 56109
rect 12363 56053 12431 56109
rect 12487 56053 12497 56109
rect 12297 56043 12497 56053
rect 305 55748 2117 55758
rect 305 55692 315 55748
rect 371 55692 439 55748
rect 495 55692 563 55748
rect 619 55692 687 55748
rect 743 55692 811 55748
rect 867 55692 935 55748
rect 991 55692 1059 55748
rect 1115 55692 1183 55748
rect 1239 55692 1307 55748
rect 1363 55692 1431 55748
rect 1487 55692 1555 55748
rect 1611 55692 1679 55748
rect 1735 55692 1803 55748
rect 1859 55692 1927 55748
rect 1983 55692 2051 55748
rect 2107 55692 2117 55748
rect 305 55624 2117 55692
rect 305 55568 315 55624
rect 371 55568 439 55624
rect 495 55568 563 55624
rect 619 55568 687 55624
rect 743 55568 811 55624
rect 867 55568 935 55624
rect 991 55568 1059 55624
rect 1115 55568 1183 55624
rect 1239 55568 1307 55624
rect 1363 55568 1431 55624
rect 1487 55568 1555 55624
rect 1611 55568 1679 55624
rect 1735 55568 1803 55624
rect 1859 55568 1927 55624
rect 1983 55568 2051 55624
rect 2107 55568 2117 55624
rect 305 55500 2117 55568
rect 305 55444 315 55500
rect 371 55444 439 55500
rect 495 55444 563 55500
rect 619 55444 687 55500
rect 743 55444 811 55500
rect 867 55444 935 55500
rect 991 55444 1059 55500
rect 1115 55444 1183 55500
rect 1239 55444 1307 55500
rect 1363 55444 1431 55500
rect 1487 55444 1555 55500
rect 1611 55444 1679 55500
rect 1735 55444 1803 55500
rect 1859 55444 1927 55500
rect 1983 55444 2051 55500
rect 2107 55444 2117 55500
rect 305 55376 2117 55444
rect 305 55320 315 55376
rect 371 55320 439 55376
rect 495 55320 563 55376
rect 619 55320 687 55376
rect 743 55320 811 55376
rect 867 55320 935 55376
rect 991 55320 1059 55376
rect 1115 55320 1183 55376
rect 1239 55320 1307 55376
rect 1363 55320 1431 55376
rect 1487 55320 1555 55376
rect 1611 55320 1679 55376
rect 1735 55320 1803 55376
rect 1859 55320 1927 55376
rect 1983 55320 2051 55376
rect 2107 55320 2117 55376
rect 305 55252 2117 55320
rect 305 55196 315 55252
rect 371 55196 439 55252
rect 495 55196 563 55252
rect 619 55196 687 55252
rect 743 55196 811 55252
rect 867 55196 935 55252
rect 991 55196 1059 55252
rect 1115 55196 1183 55252
rect 1239 55196 1307 55252
rect 1363 55196 1431 55252
rect 1487 55196 1555 55252
rect 1611 55196 1679 55252
rect 1735 55196 1803 55252
rect 1859 55196 1927 55252
rect 1983 55196 2051 55252
rect 2107 55196 2117 55252
rect 305 55128 2117 55196
rect 305 55072 315 55128
rect 371 55072 439 55128
rect 495 55072 563 55128
rect 619 55072 687 55128
rect 743 55072 811 55128
rect 867 55072 935 55128
rect 991 55072 1059 55128
rect 1115 55072 1183 55128
rect 1239 55072 1307 55128
rect 1363 55072 1431 55128
rect 1487 55072 1555 55128
rect 1611 55072 1679 55128
rect 1735 55072 1803 55128
rect 1859 55072 1927 55128
rect 1983 55072 2051 55128
rect 2107 55072 2117 55128
rect 305 55004 2117 55072
rect 305 54948 315 55004
rect 371 54948 439 55004
rect 495 54948 563 55004
rect 619 54948 687 55004
rect 743 54948 811 55004
rect 867 54948 935 55004
rect 991 54948 1059 55004
rect 1115 54948 1183 55004
rect 1239 54948 1307 55004
rect 1363 54948 1431 55004
rect 1487 54948 1555 55004
rect 1611 54948 1679 55004
rect 1735 54948 1803 55004
rect 1859 54948 1927 55004
rect 1983 54948 2051 55004
rect 2107 54948 2117 55004
rect 305 54880 2117 54948
rect 305 54824 315 54880
rect 371 54824 439 54880
rect 495 54824 563 54880
rect 619 54824 687 54880
rect 743 54824 811 54880
rect 867 54824 935 54880
rect 991 54824 1059 54880
rect 1115 54824 1183 54880
rect 1239 54824 1307 54880
rect 1363 54824 1431 54880
rect 1487 54824 1555 54880
rect 1611 54824 1679 54880
rect 1735 54824 1803 54880
rect 1859 54824 1927 54880
rect 1983 54824 2051 54880
rect 2107 54824 2117 54880
rect 305 54756 2117 54824
rect 305 54700 315 54756
rect 371 54700 439 54756
rect 495 54700 563 54756
rect 619 54700 687 54756
rect 743 54700 811 54756
rect 867 54700 935 54756
rect 991 54700 1059 54756
rect 1115 54700 1183 54756
rect 1239 54700 1307 54756
rect 1363 54700 1431 54756
rect 1487 54700 1555 54756
rect 1611 54700 1679 54756
rect 1735 54700 1803 54756
rect 1859 54700 1927 54756
rect 1983 54700 2051 54756
rect 2107 54700 2117 54756
rect 305 54632 2117 54700
rect 305 54576 315 54632
rect 371 54576 439 54632
rect 495 54576 563 54632
rect 619 54576 687 54632
rect 743 54576 811 54632
rect 867 54576 935 54632
rect 991 54576 1059 54632
rect 1115 54576 1183 54632
rect 1239 54576 1307 54632
rect 1363 54576 1431 54632
rect 1487 54576 1555 54632
rect 1611 54576 1679 54632
rect 1735 54576 1803 54632
rect 1859 54576 1927 54632
rect 1983 54576 2051 54632
rect 2107 54576 2117 54632
rect 305 54508 2117 54576
rect 305 54452 315 54508
rect 371 54452 439 54508
rect 495 54452 563 54508
rect 619 54452 687 54508
rect 743 54452 811 54508
rect 867 54452 935 54508
rect 991 54452 1059 54508
rect 1115 54452 1183 54508
rect 1239 54452 1307 54508
rect 1363 54452 1431 54508
rect 1487 54452 1555 54508
rect 1611 54452 1679 54508
rect 1735 54452 1803 54508
rect 1859 54452 1927 54508
rect 1983 54452 2051 54508
rect 2107 54452 2117 54508
rect 305 54442 2117 54452
rect 2798 55748 4734 55758
rect 2798 55692 2808 55748
rect 2864 55692 2932 55748
rect 2988 55692 3056 55748
rect 3112 55692 3180 55748
rect 3236 55692 3304 55748
rect 3360 55692 3428 55748
rect 3484 55692 3552 55748
rect 3608 55692 3676 55748
rect 3732 55692 3800 55748
rect 3856 55692 3924 55748
rect 3980 55692 4048 55748
rect 4104 55692 4172 55748
rect 4228 55692 4296 55748
rect 4352 55692 4420 55748
rect 4476 55692 4544 55748
rect 4600 55692 4668 55748
rect 4724 55692 4734 55748
rect 2798 55624 4734 55692
rect 2798 55568 2808 55624
rect 2864 55568 2932 55624
rect 2988 55568 3056 55624
rect 3112 55568 3180 55624
rect 3236 55568 3304 55624
rect 3360 55568 3428 55624
rect 3484 55568 3552 55624
rect 3608 55568 3676 55624
rect 3732 55568 3800 55624
rect 3856 55568 3924 55624
rect 3980 55568 4048 55624
rect 4104 55568 4172 55624
rect 4228 55568 4296 55624
rect 4352 55568 4420 55624
rect 4476 55568 4544 55624
rect 4600 55568 4668 55624
rect 4724 55568 4734 55624
rect 2798 55500 4734 55568
rect 2798 55444 2808 55500
rect 2864 55444 2932 55500
rect 2988 55444 3056 55500
rect 3112 55444 3180 55500
rect 3236 55444 3304 55500
rect 3360 55444 3428 55500
rect 3484 55444 3552 55500
rect 3608 55444 3676 55500
rect 3732 55444 3800 55500
rect 3856 55444 3924 55500
rect 3980 55444 4048 55500
rect 4104 55444 4172 55500
rect 4228 55444 4296 55500
rect 4352 55444 4420 55500
rect 4476 55444 4544 55500
rect 4600 55444 4668 55500
rect 4724 55444 4734 55500
rect 2798 55376 4734 55444
rect 2798 55320 2808 55376
rect 2864 55320 2932 55376
rect 2988 55320 3056 55376
rect 3112 55320 3180 55376
rect 3236 55320 3304 55376
rect 3360 55320 3428 55376
rect 3484 55320 3552 55376
rect 3608 55320 3676 55376
rect 3732 55320 3800 55376
rect 3856 55320 3924 55376
rect 3980 55320 4048 55376
rect 4104 55320 4172 55376
rect 4228 55320 4296 55376
rect 4352 55320 4420 55376
rect 4476 55320 4544 55376
rect 4600 55320 4668 55376
rect 4724 55320 4734 55376
rect 2798 55252 4734 55320
rect 2798 55196 2808 55252
rect 2864 55196 2932 55252
rect 2988 55196 3056 55252
rect 3112 55196 3180 55252
rect 3236 55196 3304 55252
rect 3360 55196 3428 55252
rect 3484 55196 3552 55252
rect 3608 55196 3676 55252
rect 3732 55196 3800 55252
rect 3856 55196 3924 55252
rect 3980 55196 4048 55252
rect 4104 55196 4172 55252
rect 4228 55196 4296 55252
rect 4352 55196 4420 55252
rect 4476 55196 4544 55252
rect 4600 55196 4668 55252
rect 4724 55196 4734 55252
rect 2798 55128 4734 55196
rect 2798 55072 2808 55128
rect 2864 55072 2932 55128
rect 2988 55072 3056 55128
rect 3112 55072 3180 55128
rect 3236 55072 3304 55128
rect 3360 55072 3428 55128
rect 3484 55072 3552 55128
rect 3608 55072 3676 55128
rect 3732 55072 3800 55128
rect 3856 55072 3924 55128
rect 3980 55072 4048 55128
rect 4104 55072 4172 55128
rect 4228 55072 4296 55128
rect 4352 55072 4420 55128
rect 4476 55072 4544 55128
rect 4600 55072 4668 55128
rect 4724 55072 4734 55128
rect 2798 55004 4734 55072
rect 2798 54948 2808 55004
rect 2864 54948 2932 55004
rect 2988 54948 3056 55004
rect 3112 54948 3180 55004
rect 3236 54948 3304 55004
rect 3360 54948 3428 55004
rect 3484 54948 3552 55004
rect 3608 54948 3676 55004
rect 3732 54948 3800 55004
rect 3856 54948 3924 55004
rect 3980 54948 4048 55004
rect 4104 54948 4172 55004
rect 4228 54948 4296 55004
rect 4352 54948 4420 55004
rect 4476 54948 4544 55004
rect 4600 54948 4668 55004
rect 4724 54948 4734 55004
rect 2798 54880 4734 54948
rect 2798 54824 2808 54880
rect 2864 54824 2932 54880
rect 2988 54824 3056 54880
rect 3112 54824 3180 54880
rect 3236 54824 3304 54880
rect 3360 54824 3428 54880
rect 3484 54824 3552 54880
rect 3608 54824 3676 54880
rect 3732 54824 3800 54880
rect 3856 54824 3924 54880
rect 3980 54824 4048 54880
rect 4104 54824 4172 54880
rect 4228 54824 4296 54880
rect 4352 54824 4420 54880
rect 4476 54824 4544 54880
rect 4600 54824 4668 54880
rect 4724 54824 4734 54880
rect 2798 54756 4734 54824
rect 2798 54700 2808 54756
rect 2864 54700 2932 54756
rect 2988 54700 3056 54756
rect 3112 54700 3180 54756
rect 3236 54700 3304 54756
rect 3360 54700 3428 54756
rect 3484 54700 3552 54756
rect 3608 54700 3676 54756
rect 3732 54700 3800 54756
rect 3856 54700 3924 54756
rect 3980 54700 4048 54756
rect 4104 54700 4172 54756
rect 4228 54700 4296 54756
rect 4352 54700 4420 54756
rect 4476 54700 4544 54756
rect 4600 54700 4668 54756
rect 4724 54700 4734 54756
rect 2798 54632 4734 54700
rect 2798 54576 2808 54632
rect 2864 54576 2932 54632
rect 2988 54576 3056 54632
rect 3112 54576 3180 54632
rect 3236 54576 3304 54632
rect 3360 54576 3428 54632
rect 3484 54576 3552 54632
rect 3608 54576 3676 54632
rect 3732 54576 3800 54632
rect 3856 54576 3924 54632
rect 3980 54576 4048 54632
rect 4104 54576 4172 54632
rect 4228 54576 4296 54632
rect 4352 54576 4420 54632
rect 4476 54576 4544 54632
rect 4600 54576 4668 54632
rect 4724 54576 4734 54632
rect 2798 54508 4734 54576
rect 2798 54452 2808 54508
rect 2864 54452 2932 54508
rect 2988 54452 3056 54508
rect 3112 54452 3180 54508
rect 3236 54452 3304 54508
rect 3360 54452 3428 54508
rect 3484 54452 3552 54508
rect 3608 54452 3676 54508
rect 3732 54452 3800 54508
rect 3856 54452 3924 54508
rect 3980 54452 4048 54508
rect 4104 54452 4172 54508
rect 4228 54452 4296 54508
rect 4352 54452 4420 54508
rect 4476 54452 4544 54508
rect 4600 54452 4668 54508
rect 4724 54452 4734 54508
rect 2798 54442 4734 54452
rect 5168 55748 7104 55758
rect 5168 55692 5178 55748
rect 5234 55692 5302 55748
rect 5358 55692 5426 55748
rect 5482 55692 5550 55748
rect 5606 55692 5674 55748
rect 5730 55692 5798 55748
rect 5854 55692 5922 55748
rect 5978 55692 6046 55748
rect 6102 55692 6170 55748
rect 6226 55692 6294 55748
rect 6350 55692 6418 55748
rect 6474 55692 6542 55748
rect 6598 55692 6666 55748
rect 6722 55692 6790 55748
rect 6846 55692 6914 55748
rect 6970 55692 7038 55748
rect 7094 55692 7104 55748
rect 5168 55624 7104 55692
rect 5168 55568 5178 55624
rect 5234 55568 5302 55624
rect 5358 55568 5426 55624
rect 5482 55568 5550 55624
rect 5606 55568 5674 55624
rect 5730 55568 5798 55624
rect 5854 55568 5922 55624
rect 5978 55568 6046 55624
rect 6102 55568 6170 55624
rect 6226 55568 6294 55624
rect 6350 55568 6418 55624
rect 6474 55568 6542 55624
rect 6598 55568 6666 55624
rect 6722 55568 6790 55624
rect 6846 55568 6914 55624
rect 6970 55568 7038 55624
rect 7094 55568 7104 55624
rect 5168 55500 7104 55568
rect 5168 55444 5178 55500
rect 5234 55444 5302 55500
rect 5358 55444 5426 55500
rect 5482 55444 5550 55500
rect 5606 55444 5674 55500
rect 5730 55444 5798 55500
rect 5854 55444 5922 55500
rect 5978 55444 6046 55500
rect 6102 55444 6170 55500
rect 6226 55444 6294 55500
rect 6350 55444 6418 55500
rect 6474 55444 6542 55500
rect 6598 55444 6666 55500
rect 6722 55444 6790 55500
rect 6846 55444 6914 55500
rect 6970 55444 7038 55500
rect 7094 55444 7104 55500
rect 5168 55376 7104 55444
rect 5168 55320 5178 55376
rect 5234 55320 5302 55376
rect 5358 55320 5426 55376
rect 5482 55320 5550 55376
rect 5606 55320 5674 55376
rect 5730 55320 5798 55376
rect 5854 55320 5922 55376
rect 5978 55320 6046 55376
rect 6102 55320 6170 55376
rect 6226 55320 6294 55376
rect 6350 55320 6418 55376
rect 6474 55320 6542 55376
rect 6598 55320 6666 55376
rect 6722 55320 6790 55376
rect 6846 55320 6914 55376
rect 6970 55320 7038 55376
rect 7094 55320 7104 55376
rect 5168 55252 7104 55320
rect 5168 55196 5178 55252
rect 5234 55196 5302 55252
rect 5358 55196 5426 55252
rect 5482 55196 5550 55252
rect 5606 55196 5674 55252
rect 5730 55196 5798 55252
rect 5854 55196 5922 55252
rect 5978 55196 6046 55252
rect 6102 55196 6170 55252
rect 6226 55196 6294 55252
rect 6350 55196 6418 55252
rect 6474 55196 6542 55252
rect 6598 55196 6666 55252
rect 6722 55196 6790 55252
rect 6846 55196 6914 55252
rect 6970 55196 7038 55252
rect 7094 55196 7104 55252
rect 5168 55128 7104 55196
rect 5168 55072 5178 55128
rect 5234 55072 5302 55128
rect 5358 55072 5426 55128
rect 5482 55072 5550 55128
rect 5606 55072 5674 55128
rect 5730 55072 5798 55128
rect 5854 55072 5922 55128
rect 5978 55072 6046 55128
rect 6102 55072 6170 55128
rect 6226 55072 6294 55128
rect 6350 55072 6418 55128
rect 6474 55072 6542 55128
rect 6598 55072 6666 55128
rect 6722 55072 6790 55128
rect 6846 55072 6914 55128
rect 6970 55072 7038 55128
rect 7094 55072 7104 55128
rect 5168 55004 7104 55072
rect 5168 54948 5178 55004
rect 5234 54948 5302 55004
rect 5358 54948 5426 55004
rect 5482 54948 5550 55004
rect 5606 54948 5674 55004
rect 5730 54948 5798 55004
rect 5854 54948 5922 55004
rect 5978 54948 6046 55004
rect 6102 54948 6170 55004
rect 6226 54948 6294 55004
rect 6350 54948 6418 55004
rect 6474 54948 6542 55004
rect 6598 54948 6666 55004
rect 6722 54948 6790 55004
rect 6846 54948 6914 55004
rect 6970 54948 7038 55004
rect 7094 54948 7104 55004
rect 5168 54880 7104 54948
rect 5168 54824 5178 54880
rect 5234 54824 5302 54880
rect 5358 54824 5426 54880
rect 5482 54824 5550 54880
rect 5606 54824 5674 54880
rect 5730 54824 5798 54880
rect 5854 54824 5922 54880
rect 5978 54824 6046 54880
rect 6102 54824 6170 54880
rect 6226 54824 6294 54880
rect 6350 54824 6418 54880
rect 6474 54824 6542 54880
rect 6598 54824 6666 54880
rect 6722 54824 6790 54880
rect 6846 54824 6914 54880
rect 6970 54824 7038 54880
rect 7094 54824 7104 54880
rect 5168 54756 7104 54824
rect 5168 54700 5178 54756
rect 5234 54700 5302 54756
rect 5358 54700 5426 54756
rect 5482 54700 5550 54756
rect 5606 54700 5674 54756
rect 5730 54700 5798 54756
rect 5854 54700 5922 54756
rect 5978 54700 6046 54756
rect 6102 54700 6170 54756
rect 6226 54700 6294 54756
rect 6350 54700 6418 54756
rect 6474 54700 6542 54756
rect 6598 54700 6666 54756
rect 6722 54700 6790 54756
rect 6846 54700 6914 54756
rect 6970 54700 7038 54756
rect 7094 54700 7104 54756
rect 5168 54632 7104 54700
rect 5168 54576 5178 54632
rect 5234 54576 5302 54632
rect 5358 54576 5426 54632
rect 5482 54576 5550 54632
rect 5606 54576 5674 54632
rect 5730 54576 5798 54632
rect 5854 54576 5922 54632
rect 5978 54576 6046 54632
rect 6102 54576 6170 54632
rect 6226 54576 6294 54632
rect 6350 54576 6418 54632
rect 6474 54576 6542 54632
rect 6598 54576 6666 54632
rect 6722 54576 6790 54632
rect 6846 54576 6914 54632
rect 6970 54576 7038 54632
rect 7094 54576 7104 54632
rect 5168 54508 7104 54576
rect 5168 54452 5178 54508
rect 5234 54452 5302 54508
rect 5358 54452 5426 54508
rect 5482 54452 5550 54508
rect 5606 54452 5674 54508
rect 5730 54452 5798 54508
rect 5854 54452 5922 54508
rect 5978 54452 6046 54508
rect 6102 54452 6170 54508
rect 6226 54452 6294 54508
rect 6350 54452 6418 54508
rect 6474 54452 6542 54508
rect 6598 54452 6666 54508
rect 6722 54452 6790 54508
rect 6846 54452 6914 54508
rect 6970 54452 7038 54508
rect 7094 54452 7104 54508
rect 5168 54442 7104 54452
rect 7874 55748 9810 55758
rect 7874 55692 7884 55748
rect 7940 55692 8008 55748
rect 8064 55692 8132 55748
rect 8188 55692 8256 55748
rect 8312 55692 8380 55748
rect 8436 55692 8504 55748
rect 8560 55692 8628 55748
rect 8684 55692 8752 55748
rect 8808 55692 8876 55748
rect 8932 55692 9000 55748
rect 9056 55692 9124 55748
rect 9180 55692 9248 55748
rect 9304 55692 9372 55748
rect 9428 55692 9496 55748
rect 9552 55692 9620 55748
rect 9676 55692 9744 55748
rect 9800 55692 9810 55748
rect 7874 55624 9810 55692
rect 7874 55568 7884 55624
rect 7940 55568 8008 55624
rect 8064 55568 8132 55624
rect 8188 55568 8256 55624
rect 8312 55568 8380 55624
rect 8436 55568 8504 55624
rect 8560 55568 8628 55624
rect 8684 55568 8752 55624
rect 8808 55568 8876 55624
rect 8932 55568 9000 55624
rect 9056 55568 9124 55624
rect 9180 55568 9248 55624
rect 9304 55568 9372 55624
rect 9428 55568 9496 55624
rect 9552 55568 9620 55624
rect 9676 55568 9744 55624
rect 9800 55568 9810 55624
rect 7874 55500 9810 55568
rect 7874 55444 7884 55500
rect 7940 55444 8008 55500
rect 8064 55444 8132 55500
rect 8188 55444 8256 55500
rect 8312 55444 8380 55500
rect 8436 55444 8504 55500
rect 8560 55444 8628 55500
rect 8684 55444 8752 55500
rect 8808 55444 8876 55500
rect 8932 55444 9000 55500
rect 9056 55444 9124 55500
rect 9180 55444 9248 55500
rect 9304 55444 9372 55500
rect 9428 55444 9496 55500
rect 9552 55444 9620 55500
rect 9676 55444 9744 55500
rect 9800 55444 9810 55500
rect 7874 55376 9810 55444
rect 7874 55320 7884 55376
rect 7940 55320 8008 55376
rect 8064 55320 8132 55376
rect 8188 55320 8256 55376
rect 8312 55320 8380 55376
rect 8436 55320 8504 55376
rect 8560 55320 8628 55376
rect 8684 55320 8752 55376
rect 8808 55320 8876 55376
rect 8932 55320 9000 55376
rect 9056 55320 9124 55376
rect 9180 55320 9248 55376
rect 9304 55320 9372 55376
rect 9428 55320 9496 55376
rect 9552 55320 9620 55376
rect 9676 55320 9744 55376
rect 9800 55320 9810 55376
rect 7874 55252 9810 55320
rect 7874 55196 7884 55252
rect 7940 55196 8008 55252
rect 8064 55196 8132 55252
rect 8188 55196 8256 55252
rect 8312 55196 8380 55252
rect 8436 55196 8504 55252
rect 8560 55196 8628 55252
rect 8684 55196 8752 55252
rect 8808 55196 8876 55252
rect 8932 55196 9000 55252
rect 9056 55196 9124 55252
rect 9180 55196 9248 55252
rect 9304 55196 9372 55252
rect 9428 55196 9496 55252
rect 9552 55196 9620 55252
rect 9676 55196 9744 55252
rect 9800 55196 9810 55252
rect 7874 55128 9810 55196
rect 7874 55072 7884 55128
rect 7940 55072 8008 55128
rect 8064 55072 8132 55128
rect 8188 55072 8256 55128
rect 8312 55072 8380 55128
rect 8436 55072 8504 55128
rect 8560 55072 8628 55128
rect 8684 55072 8752 55128
rect 8808 55072 8876 55128
rect 8932 55072 9000 55128
rect 9056 55072 9124 55128
rect 9180 55072 9248 55128
rect 9304 55072 9372 55128
rect 9428 55072 9496 55128
rect 9552 55072 9620 55128
rect 9676 55072 9744 55128
rect 9800 55072 9810 55128
rect 7874 55004 9810 55072
rect 7874 54948 7884 55004
rect 7940 54948 8008 55004
rect 8064 54948 8132 55004
rect 8188 54948 8256 55004
rect 8312 54948 8380 55004
rect 8436 54948 8504 55004
rect 8560 54948 8628 55004
rect 8684 54948 8752 55004
rect 8808 54948 8876 55004
rect 8932 54948 9000 55004
rect 9056 54948 9124 55004
rect 9180 54948 9248 55004
rect 9304 54948 9372 55004
rect 9428 54948 9496 55004
rect 9552 54948 9620 55004
rect 9676 54948 9744 55004
rect 9800 54948 9810 55004
rect 7874 54880 9810 54948
rect 7874 54824 7884 54880
rect 7940 54824 8008 54880
rect 8064 54824 8132 54880
rect 8188 54824 8256 54880
rect 8312 54824 8380 54880
rect 8436 54824 8504 54880
rect 8560 54824 8628 54880
rect 8684 54824 8752 54880
rect 8808 54824 8876 54880
rect 8932 54824 9000 54880
rect 9056 54824 9124 54880
rect 9180 54824 9248 54880
rect 9304 54824 9372 54880
rect 9428 54824 9496 54880
rect 9552 54824 9620 54880
rect 9676 54824 9744 54880
rect 9800 54824 9810 54880
rect 7874 54756 9810 54824
rect 7874 54700 7884 54756
rect 7940 54700 8008 54756
rect 8064 54700 8132 54756
rect 8188 54700 8256 54756
rect 8312 54700 8380 54756
rect 8436 54700 8504 54756
rect 8560 54700 8628 54756
rect 8684 54700 8752 54756
rect 8808 54700 8876 54756
rect 8932 54700 9000 54756
rect 9056 54700 9124 54756
rect 9180 54700 9248 54756
rect 9304 54700 9372 54756
rect 9428 54700 9496 54756
rect 9552 54700 9620 54756
rect 9676 54700 9744 54756
rect 9800 54700 9810 54756
rect 7874 54632 9810 54700
rect 7874 54576 7884 54632
rect 7940 54576 8008 54632
rect 8064 54576 8132 54632
rect 8188 54576 8256 54632
rect 8312 54576 8380 54632
rect 8436 54576 8504 54632
rect 8560 54576 8628 54632
rect 8684 54576 8752 54632
rect 8808 54576 8876 54632
rect 8932 54576 9000 54632
rect 9056 54576 9124 54632
rect 9180 54576 9248 54632
rect 9304 54576 9372 54632
rect 9428 54576 9496 54632
rect 9552 54576 9620 54632
rect 9676 54576 9744 54632
rect 9800 54576 9810 54632
rect 7874 54508 9810 54576
rect 7874 54452 7884 54508
rect 7940 54452 8008 54508
rect 8064 54452 8132 54508
rect 8188 54452 8256 54508
rect 8312 54452 8380 54508
rect 8436 54452 8504 54508
rect 8560 54452 8628 54508
rect 8684 54452 8752 54508
rect 8808 54452 8876 54508
rect 8932 54452 9000 54508
rect 9056 54452 9124 54508
rect 9180 54452 9248 54508
rect 9304 54452 9372 54508
rect 9428 54452 9496 54508
rect 9552 54452 9620 54508
rect 9676 54452 9744 54508
rect 9800 54452 9810 54508
rect 7874 54442 9810 54452
rect 10244 55748 12180 55758
rect 10244 55692 10254 55748
rect 10310 55692 10378 55748
rect 10434 55692 10502 55748
rect 10558 55692 10626 55748
rect 10682 55692 10750 55748
rect 10806 55692 10874 55748
rect 10930 55692 10998 55748
rect 11054 55692 11122 55748
rect 11178 55692 11246 55748
rect 11302 55692 11370 55748
rect 11426 55692 11494 55748
rect 11550 55692 11618 55748
rect 11674 55692 11742 55748
rect 11798 55692 11866 55748
rect 11922 55692 11990 55748
rect 12046 55692 12114 55748
rect 12170 55692 12180 55748
rect 10244 55624 12180 55692
rect 10244 55568 10254 55624
rect 10310 55568 10378 55624
rect 10434 55568 10502 55624
rect 10558 55568 10626 55624
rect 10682 55568 10750 55624
rect 10806 55568 10874 55624
rect 10930 55568 10998 55624
rect 11054 55568 11122 55624
rect 11178 55568 11246 55624
rect 11302 55568 11370 55624
rect 11426 55568 11494 55624
rect 11550 55568 11618 55624
rect 11674 55568 11742 55624
rect 11798 55568 11866 55624
rect 11922 55568 11990 55624
rect 12046 55568 12114 55624
rect 12170 55568 12180 55624
rect 10244 55500 12180 55568
rect 10244 55444 10254 55500
rect 10310 55444 10378 55500
rect 10434 55444 10502 55500
rect 10558 55444 10626 55500
rect 10682 55444 10750 55500
rect 10806 55444 10874 55500
rect 10930 55444 10998 55500
rect 11054 55444 11122 55500
rect 11178 55444 11246 55500
rect 11302 55444 11370 55500
rect 11426 55444 11494 55500
rect 11550 55444 11618 55500
rect 11674 55444 11742 55500
rect 11798 55444 11866 55500
rect 11922 55444 11990 55500
rect 12046 55444 12114 55500
rect 12170 55444 12180 55500
rect 10244 55376 12180 55444
rect 10244 55320 10254 55376
rect 10310 55320 10378 55376
rect 10434 55320 10502 55376
rect 10558 55320 10626 55376
rect 10682 55320 10750 55376
rect 10806 55320 10874 55376
rect 10930 55320 10998 55376
rect 11054 55320 11122 55376
rect 11178 55320 11246 55376
rect 11302 55320 11370 55376
rect 11426 55320 11494 55376
rect 11550 55320 11618 55376
rect 11674 55320 11742 55376
rect 11798 55320 11866 55376
rect 11922 55320 11990 55376
rect 12046 55320 12114 55376
rect 12170 55320 12180 55376
rect 10244 55252 12180 55320
rect 10244 55196 10254 55252
rect 10310 55196 10378 55252
rect 10434 55196 10502 55252
rect 10558 55196 10626 55252
rect 10682 55196 10750 55252
rect 10806 55196 10874 55252
rect 10930 55196 10998 55252
rect 11054 55196 11122 55252
rect 11178 55196 11246 55252
rect 11302 55196 11370 55252
rect 11426 55196 11494 55252
rect 11550 55196 11618 55252
rect 11674 55196 11742 55252
rect 11798 55196 11866 55252
rect 11922 55196 11990 55252
rect 12046 55196 12114 55252
rect 12170 55196 12180 55252
rect 10244 55128 12180 55196
rect 10244 55072 10254 55128
rect 10310 55072 10378 55128
rect 10434 55072 10502 55128
rect 10558 55072 10626 55128
rect 10682 55072 10750 55128
rect 10806 55072 10874 55128
rect 10930 55072 10998 55128
rect 11054 55072 11122 55128
rect 11178 55072 11246 55128
rect 11302 55072 11370 55128
rect 11426 55072 11494 55128
rect 11550 55072 11618 55128
rect 11674 55072 11742 55128
rect 11798 55072 11866 55128
rect 11922 55072 11990 55128
rect 12046 55072 12114 55128
rect 12170 55072 12180 55128
rect 10244 55004 12180 55072
rect 10244 54948 10254 55004
rect 10310 54948 10378 55004
rect 10434 54948 10502 55004
rect 10558 54948 10626 55004
rect 10682 54948 10750 55004
rect 10806 54948 10874 55004
rect 10930 54948 10998 55004
rect 11054 54948 11122 55004
rect 11178 54948 11246 55004
rect 11302 54948 11370 55004
rect 11426 54948 11494 55004
rect 11550 54948 11618 55004
rect 11674 54948 11742 55004
rect 11798 54948 11866 55004
rect 11922 54948 11990 55004
rect 12046 54948 12114 55004
rect 12170 54948 12180 55004
rect 10244 54880 12180 54948
rect 10244 54824 10254 54880
rect 10310 54824 10378 54880
rect 10434 54824 10502 54880
rect 10558 54824 10626 54880
rect 10682 54824 10750 54880
rect 10806 54824 10874 54880
rect 10930 54824 10998 54880
rect 11054 54824 11122 54880
rect 11178 54824 11246 54880
rect 11302 54824 11370 54880
rect 11426 54824 11494 54880
rect 11550 54824 11618 54880
rect 11674 54824 11742 54880
rect 11798 54824 11866 54880
rect 11922 54824 11990 54880
rect 12046 54824 12114 54880
rect 12170 54824 12180 54880
rect 10244 54756 12180 54824
rect 10244 54700 10254 54756
rect 10310 54700 10378 54756
rect 10434 54700 10502 54756
rect 10558 54700 10626 54756
rect 10682 54700 10750 54756
rect 10806 54700 10874 54756
rect 10930 54700 10998 54756
rect 11054 54700 11122 54756
rect 11178 54700 11246 54756
rect 11302 54700 11370 54756
rect 11426 54700 11494 54756
rect 11550 54700 11618 54756
rect 11674 54700 11742 54756
rect 11798 54700 11866 54756
rect 11922 54700 11990 54756
rect 12046 54700 12114 54756
rect 12170 54700 12180 54756
rect 10244 54632 12180 54700
rect 10244 54576 10254 54632
rect 10310 54576 10378 54632
rect 10434 54576 10502 54632
rect 10558 54576 10626 54632
rect 10682 54576 10750 54632
rect 10806 54576 10874 54632
rect 10930 54576 10998 54632
rect 11054 54576 11122 54632
rect 11178 54576 11246 54632
rect 11302 54576 11370 54632
rect 11426 54576 11494 54632
rect 11550 54576 11618 54632
rect 11674 54576 11742 54632
rect 11798 54576 11866 54632
rect 11922 54576 11990 54632
rect 12046 54576 12114 54632
rect 12170 54576 12180 54632
rect 10244 54508 12180 54576
rect 10244 54452 10254 54508
rect 10310 54452 10378 54508
rect 10434 54452 10502 54508
rect 10558 54452 10626 54508
rect 10682 54452 10750 54508
rect 10806 54452 10874 54508
rect 10930 54452 10998 54508
rect 11054 54452 11122 54508
rect 11178 54452 11246 54508
rect 11302 54452 11370 54508
rect 11426 54452 11494 54508
rect 11550 54452 11618 54508
rect 11674 54452 11742 54508
rect 11798 54452 11866 54508
rect 11922 54452 11990 54508
rect 12046 54452 12114 54508
rect 12170 54452 12180 54508
rect 10244 54442 12180 54452
rect 12861 55748 14673 55758
rect 12861 55692 12871 55748
rect 12927 55692 12995 55748
rect 13051 55692 13119 55748
rect 13175 55692 13243 55748
rect 13299 55692 13367 55748
rect 13423 55692 13491 55748
rect 13547 55692 13615 55748
rect 13671 55692 13739 55748
rect 13795 55692 13863 55748
rect 13919 55692 13987 55748
rect 14043 55692 14111 55748
rect 14167 55692 14235 55748
rect 14291 55692 14359 55748
rect 14415 55692 14483 55748
rect 14539 55692 14607 55748
rect 14663 55692 14673 55748
rect 12861 55624 14673 55692
rect 12861 55568 12871 55624
rect 12927 55568 12995 55624
rect 13051 55568 13119 55624
rect 13175 55568 13243 55624
rect 13299 55568 13367 55624
rect 13423 55568 13491 55624
rect 13547 55568 13615 55624
rect 13671 55568 13739 55624
rect 13795 55568 13863 55624
rect 13919 55568 13987 55624
rect 14043 55568 14111 55624
rect 14167 55568 14235 55624
rect 14291 55568 14359 55624
rect 14415 55568 14483 55624
rect 14539 55568 14607 55624
rect 14663 55568 14673 55624
rect 12861 55500 14673 55568
rect 12861 55444 12871 55500
rect 12927 55444 12995 55500
rect 13051 55444 13119 55500
rect 13175 55444 13243 55500
rect 13299 55444 13367 55500
rect 13423 55444 13491 55500
rect 13547 55444 13615 55500
rect 13671 55444 13739 55500
rect 13795 55444 13863 55500
rect 13919 55444 13987 55500
rect 14043 55444 14111 55500
rect 14167 55444 14235 55500
rect 14291 55444 14359 55500
rect 14415 55444 14483 55500
rect 14539 55444 14607 55500
rect 14663 55444 14673 55500
rect 12861 55376 14673 55444
rect 12861 55320 12871 55376
rect 12927 55320 12995 55376
rect 13051 55320 13119 55376
rect 13175 55320 13243 55376
rect 13299 55320 13367 55376
rect 13423 55320 13491 55376
rect 13547 55320 13615 55376
rect 13671 55320 13739 55376
rect 13795 55320 13863 55376
rect 13919 55320 13987 55376
rect 14043 55320 14111 55376
rect 14167 55320 14235 55376
rect 14291 55320 14359 55376
rect 14415 55320 14483 55376
rect 14539 55320 14607 55376
rect 14663 55320 14673 55376
rect 12861 55252 14673 55320
rect 12861 55196 12871 55252
rect 12927 55196 12995 55252
rect 13051 55196 13119 55252
rect 13175 55196 13243 55252
rect 13299 55196 13367 55252
rect 13423 55196 13491 55252
rect 13547 55196 13615 55252
rect 13671 55196 13739 55252
rect 13795 55196 13863 55252
rect 13919 55196 13987 55252
rect 14043 55196 14111 55252
rect 14167 55196 14235 55252
rect 14291 55196 14359 55252
rect 14415 55196 14483 55252
rect 14539 55196 14607 55252
rect 14663 55196 14673 55252
rect 12861 55128 14673 55196
rect 12861 55072 12871 55128
rect 12927 55072 12995 55128
rect 13051 55072 13119 55128
rect 13175 55072 13243 55128
rect 13299 55072 13367 55128
rect 13423 55072 13491 55128
rect 13547 55072 13615 55128
rect 13671 55072 13739 55128
rect 13795 55072 13863 55128
rect 13919 55072 13987 55128
rect 14043 55072 14111 55128
rect 14167 55072 14235 55128
rect 14291 55072 14359 55128
rect 14415 55072 14483 55128
rect 14539 55072 14607 55128
rect 14663 55072 14673 55128
rect 12861 55004 14673 55072
rect 12861 54948 12871 55004
rect 12927 54948 12995 55004
rect 13051 54948 13119 55004
rect 13175 54948 13243 55004
rect 13299 54948 13367 55004
rect 13423 54948 13491 55004
rect 13547 54948 13615 55004
rect 13671 54948 13739 55004
rect 13795 54948 13863 55004
rect 13919 54948 13987 55004
rect 14043 54948 14111 55004
rect 14167 54948 14235 55004
rect 14291 54948 14359 55004
rect 14415 54948 14483 55004
rect 14539 54948 14607 55004
rect 14663 54948 14673 55004
rect 12861 54880 14673 54948
rect 12861 54824 12871 54880
rect 12927 54824 12995 54880
rect 13051 54824 13119 54880
rect 13175 54824 13243 54880
rect 13299 54824 13367 54880
rect 13423 54824 13491 54880
rect 13547 54824 13615 54880
rect 13671 54824 13739 54880
rect 13795 54824 13863 54880
rect 13919 54824 13987 54880
rect 14043 54824 14111 54880
rect 14167 54824 14235 54880
rect 14291 54824 14359 54880
rect 14415 54824 14483 54880
rect 14539 54824 14607 54880
rect 14663 54824 14673 54880
rect 12861 54756 14673 54824
rect 12861 54700 12871 54756
rect 12927 54700 12995 54756
rect 13051 54700 13119 54756
rect 13175 54700 13243 54756
rect 13299 54700 13367 54756
rect 13423 54700 13491 54756
rect 13547 54700 13615 54756
rect 13671 54700 13739 54756
rect 13795 54700 13863 54756
rect 13919 54700 13987 54756
rect 14043 54700 14111 54756
rect 14167 54700 14235 54756
rect 14291 54700 14359 54756
rect 14415 54700 14483 54756
rect 14539 54700 14607 54756
rect 14663 54700 14673 54756
rect 12861 54632 14673 54700
rect 12861 54576 12871 54632
rect 12927 54576 12995 54632
rect 13051 54576 13119 54632
rect 13175 54576 13243 54632
rect 13299 54576 13367 54632
rect 13423 54576 13491 54632
rect 13547 54576 13615 54632
rect 13671 54576 13739 54632
rect 13795 54576 13863 54632
rect 13919 54576 13987 54632
rect 14043 54576 14111 54632
rect 14167 54576 14235 54632
rect 14291 54576 14359 54632
rect 14415 54576 14483 54632
rect 14539 54576 14607 54632
rect 14663 54576 14673 54632
rect 12861 54508 14673 54576
rect 12861 54452 12871 54508
rect 12927 54452 12995 54508
rect 13051 54452 13119 54508
rect 13175 54452 13243 54508
rect 13299 54452 13367 54508
rect 13423 54452 13491 54508
rect 13547 54452 13615 54508
rect 13671 54452 13739 54508
rect 13795 54452 13863 54508
rect 13919 54452 13987 54508
rect 14043 54452 14111 54508
rect 14167 54452 14235 54508
rect 14291 54452 14359 54508
rect 14415 54452 14483 54508
rect 14539 54452 14607 54508
rect 14663 54452 14673 54508
rect 12861 54442 14673 54452
rect 2481 54148 2681 54158
rect 2481 54092 2491 54148
rect 2547 54092 2615 54148
rect 2671 54092 2681 54148
rect 2481 54024 2681 54092
rect 2481 53968 2491 54024
rect 2547 53968 2615 54024
rect 2671 53968 2681 54024
rect 2481 53900 2681 53968
rect 2481 53844 2491 53900
rect 2547 53844 2615 53900
rect 2671 53844 2681 53900
rect 2481 53776 2681 53844
rect 2481 53720 2491 53776
rect 2547 53720 2615 53776
rect 2671 53720 2681 53776
rect 2481 53652 2681 53720
rect 2481 53596 2491 53652
rect 2547 53596 2615 53652
rect 2671 53596 2681 53652
rect 2481 53528 2681 53596
rect 2481 53472 2491 53528
rect 2547 53472 2615 53528
rect 2671 53472 2681 53528
rect 2481 53404 2681 53472
rect 2481 53348 2491 53404
rect 2547 53348 2615 53404
rect 2671 53348 2681 53404
rect 2481 53280 2681 53348
rect 2481 53224 2491 53280
rect 2547 53224 2615 53280
rect 2671 53224 2681 53280
rect 2481 53156 2681 53224
rect 2481 53100 2491 53156
rect 2547 53100 2615 53156
rect 2671 53100 2681 53156
rect 2481 53032 2681 53100
rect 2481 52976 2491 53032
rect 2547 52976 2615 53032
rect 2671 52976 2681 53032
rect 2481 52908 2681 52976
rect 2481 52852 2491 52908
rect 2547 52852 2615 52908
rect 2671 52852 2681 52908
rect 2481 52842 2681 52852
rect 4851 54148 5051 54158
rect 4851 54092 4861 54148
rect 4917 54092 4985 54148
rect 5041 54092 5051 54148
rect 4851 54024 5051 54092
rect 4851 53968 4861 54024
rect 4917 53968 4985 54024
rect 5041 53968 5051 54024
rect 4851 53900 5051 53968
rect 4851 53844 4861 53900
rect 4917 53844 4985 53900
rect 5041 53844 5051 53900
rect 4851 53776 5051 53844
rect 4851 53720 4861 53776
rect 4917 53720 4985 53776
rect 5041 53720 5051 53776
rect 4851 53652 5051 53720
rect 4851 53596 4861 53652
rect 4917 53596 4985 53652
rect 5041 53596 5051 53652
rect 4851 53528 5051 53596
rect 4851 53472 4861 53528
rect 4917 53472 4985 53528
rect 5041 53472 5051 53528
rect 4851 53404 5051 53472
rect 4851 53348 4861 53404
rect 4917 53348 4985 53404
rect 5041 53348 5051 53404
rect 4851 53280 5051 53348
rect 4851 53224 4861 53280
rect 4917 53224 4985 53280
rect 5041 53224 5051 53280
rect 4851 53156 5051 53224
rect 4851 53100 4861 53156
rect 4917 53100 4985 53156
rect 5041 53100 5051 53156
rect 4851 53032 5051 53100
rect 4851 52976 4861 53032
rect 4917 52976 4985 53032
rect 5041 52976 5051 53032
rect 4851 52908 5051 52976
rect 4851 52852 4861 52908
rect 4917 52852 4985 52908
rect 5041 52852 5051 52908
rect 4851 52842 5051 52852
rect 7265 54148 7713 54158
rect 7265 54092 7275 54148
rect 7331 54092 7399 54148
rect 7455 54092 7523 54148
rect 7579 54092 7647 54148
rect 7703 54092 7713 54148
rect 7265 54024 7713 54092
rect 7265 53968 7275 54024
rect 7331 53968 7399 54024
rect 7455 53968 7523 54024
rect 7579 53968 7647 54024
rect 7703 53968 7713 54024
rect 7265 53900 7713 53968
rect 7265 53844 7275 53900
rect 7331 53844 7399 53900
rect 7455 53844 7523 53900
rect 7579 53844 7647 53900
rect 7703 53844 7713 53900
rect 7265 53776 7713 53844
rect 7265 53720 7275 53776
rect 7331 53720 7399 53776
rect 7455 53720 7523 53776
rect 7579 53720 7647 53776
rect 7703 53720 7713 53776
rect 7265 53652 7713 53720
rect 7265 53596 7275 53652
rect 7331 53596 7399 53652
rect 7455 53596 7523 53652
rect 7579 53596 7647 53652
rect 7703 53596 7713 53652
rect 7265 53528 7713 53596
rect 7265 53472 7275 53528
rect 7331 53472 7399 53528
rect 7455 53472 7523 53528
rect 7579 53472 7647 53528
rect 7703 53472 7713 53528
rect 7265 53404 7713 53472
rect 7265 53348 7275 53404
rect 7331 53348 7399 53404
rect 7455 53348 7523 53404
rect 7579 53348 7647 53404
rect 7703 53348 7713 53404
rect 7265 53280 7713 53348
rect 7265 53224 7275 53280
rect 7331 53224 7399 53280
rect 7455 53224 7523 53280
rect 7579 53224 7647 53280
rect 7703 53224 7713 53280
rect 7265 53156 7713 53224
rect 7265 53100 7275 53156
rect 7331 53100 7399 53156
rect 7455 53100 7523 53156
rect 7579 53100 7647 53156
rect 7703 53100 7713 53156
rect 7265 53032 7713 53100
rect 7265 52976 7275 53032
rect 7331 52976 7399 53032
rect 7455 52976 7523 53032
rect 7579 52976 7647 53032
rect 7703 52976 7713 53032
rect 7265 52908 7713 52976
rect 7265 52852 7275 52908
rect 7331 52852 7399 52908
rect 7455 52852 7523 52908
rect 7579 52852 7647 52908
rect 7703 52852 7713 52908
rect 7265 52842 7713 52852
rect 9927 54148 10127 54158
rect 9927 54092 9937 54148
rect 9993 54092 10061 54148
rect 10117 54092 10127 54148
rect 9927 54024 10127 54092
rect 9927 53968 9937 54024
rect 9993 53968 10061 54024
rect 10117 53968 10127 54024
rect 9927 53900 10127 53968
rect 9927 53844 9937 53900
rect 9993 53844 10061 53900
rect 10117 53844 10127 53900
rect 9927 53776 10127 53844
rect 9927 53720 9937 53776
rect 9993 53720 10061 53776
rect 10117 53720 10127 53776
rect 9927 53652 10127 53720
rect 9927 53596 9937 53652
rect 9993 53596 10061 53652
rect 10117 53596 10127 53652
rect 9927 53528 10127 53596
rect 9927 53472 9937 53528
rect 9993 53472 10061 53528
rect 10117 53472 10127 53528
rect 9927 53404 10127 53472
rect 9927 53348 9937 53404
rect 9993 53348 10061 53404
rect 10117 53348 10127 53404
rect 9927 53280 10127 53348
rect 9927 53224 9937 53280
rect 9993 53224 10061 53280
rect 10117 53224 10127 53280
rect 9927 53156 10127 53224
rect 9927 53100 9937 53156
rect 9993 53100 10061 53156
rect 10117 53100 10127 53156
rect 9927 53032 10127 53100
rect 9927 52976 9937 53032
rect 9993 52976 10061 53032
rect 10117 52976 10127 53032
rect 9927 52908 10127 52976
rect 9927 52852 9937 52908
rect 9993 52852 10061 52908
rect 10117 52852 10127 52908
rect 9927 52842 10127 52852
rect 12297 54148 12497 54158
rect 12297 54092 12307 54148
rect 12363 54092 12431 54148
rect 12487 54092 12497 54148
rect 12297 54024 12497 54092
rect 12297 53968 12307 54024
rect 12363 53968 12431 54024
rect 12487 53968 12497 54024
rect 12297 53900 12497 53968
rect 12297 53844 12307 53900
rect 12363 53844 12431 53900
rect 12487 53844 12497 53900
rect 12297 53776 12497 53844
rect 12297 53720 12307 53776
rect 12363 53720 12431 53776
rect 12487 53720 12497 53776
rect 12297 53652 12497 53720
rect 12297 53596 12307 53652
rect 12363 53596 12431 53652
rect 12487 53596 12497 53652
rect 12297 53528 12497 53596
rect 12297 53472 12307 53528
rect 12363 53472 12431 53528
rect 12487 53472 12497 53528
rect 12297 53404 12497 53472
rect 12297 53348 12307 53404
rect 12363 53348 12431 53404
rect 12487 53348 12497 53404
rect 12297 53280 12497 53348
rect 12297 53224 12307 53280
rect 12363 53224 12431 53280
rect 12487 53224 12497 53280
rect 12297 53156 12497 53224
rect 12297 53100 12307 53156
rect 12363 53100 12431 53156
rect 12487 53100 12497 53156
rect 12297 53032 12497 53100
rect 12297 52976 12307 53032
rect 12363 52976 12431 53032
rect 12487 52976 12497 53032
rect 12297 52908 12497 52976
rect 12297 52852 12307 52908
rect 12363 52852 12431 52908
rect 12487 52852 12497 52908
rect 12297 52842 12497 52852
rect 10 52576 86 52586
rect 10 51224 20 52576
rect 76 51224 86 52576
rect 14892 52576 14968 52586
rect 2279 52521 2355 52531
rect 2279 52465 2289 52521
rect 2345 52465 2355 52521
rect 2279 52389 2355 52465
rect 2279 52333 2289 52389
rect 2345 52333 2355 52389
rect 2279 52257 2355 52333
rect 2279 52201 2289 52257
rect 2345 52201 2355 52257
rect 2279 52125 2355 52201
rect 2279 52069 2289 52125
rect 2345 52069 2355 52125
rect 2279 51993 2355 52069
rect 2279 51937 2289 51993
rect 2345 51937 2355 51993
rect 2279 51861 2355 51937
rect 2279 51805 2289 51861
rect 2345 51805 2355 51861
rect 2279 51729 2355 51805
rect 2279 51673 2289 51729
rect 2345 51673 2355 51729
rect 2279 51597 2355 51673
rect 2279 51541 2289 51597
rect 2345 51541 2355 51597
rect 2279 51465 2355 51541
rect 2279 51409 2289 51465
rect 2345 51409 2355 51465
rect 2279 51333 2355 51409
rect 2279 51277 2289 51333
rect 2345 51277 2355 51333
rect 2279 51267 2355 51277
rect 10 51214 86 51224
rect 14892 51224 14902 52576
rect 14958 51224 14968 52576
rect 14892 51214 14968 51224
rect 305 50948 2117 50958
rect 305 50892 315 50948
rect 371 50892 439 50948
rect 495 50892 563 50948
rect 619 50892 687 50948
rect 743 50892 811 50948
rect 867 50892 935 50948
rect 991 50892 1059 50948
rect 1115 50892 1183 50948
rect 1239 50892 1307 50948
rect 1363 50892 1431 50948
rect 1487 50892 1555 50948
rect 1611 50892 1679 50948
rect 1735 50892 1803 50948
rect 1859 50892 1927 50948
rect 1983 50892 2051 50948
rect 2107 50892 2117 50948
rect 305 50824 2117 50892
rect 305 50768 315 50824
rect 371 50768 439 50824
rect 495 50768 563 50824
rect 619 50768 687 50824
rect 743 50768 811 50824
rect 867 50768 935 50824
rect 991 50768 1059 50824
rect 1115 50768 1183 50824
rect 1239 50768 1307 50824
rect 1363 50768 1431 50824
rect 1487 50768 1555 50824
rect 1611 50768 1679 50824
rect 1735 50768 1803 50824
rect 1859 50768 1927 50824
rect 1983 50768 2051 50824
rect 2107 50768 2117 50824
rect 305 50700 2117 50768
rect 305 50644 315 50700
rect 371 50644 439 50700
rect 495 50644 563 50700
rect 619 50644 687 50700
rect 743 50644 811 50700
rect 867 50644 935 50700
rect 991 50644 1059 50700
rect 1115 50644 1183 50700
rect 1239 50644 1307 50700
rect 1363 50644 1431 50700
rect 1487 50644 1555 50700
rect 1611 50644 1679 50700
rect 1735 50644 1803 50700
rect 1859 50644 1927 50700
rect 1983 50644 2051 50700
rect 2107 50644 2117 50700
rect 305 50576 2117 50644
rect 305 50520 315 50576
rect 371 50520 439 50576
rect 495 50520 563 50576
rect 619 50520 687 50576
rect 743 50520 811 50576
rect 867 50520 935 50576
rect 991 50520 1059 50576
rect 1115 50520 1183 50576
rect 1239 50520 1307 50576
rect 1363 50520 1431 50576
rect 1487 50520 1555 50576
rect 1611 50520 1679 50576
rect 1735 50520 1803 50576
rect 1859 50520 1927 50576
rect 1983 50520 2051 50576
rect 2107 50520 2117 50576
rect 305 50452 2117 50520
rect 305 50396 315 50452
rect 371 50396 439 50452
rect 495 50396 563 50452
rect 619 50396 687 50452
rect 743 50396 811 50452
rect 867 50396 935 50452
rect 991 50396 1059 50452
rect 1115 50396 1183 50452
rect 1239 50396 1307 50452
rect 1363 50396 1431 50452
rect 1487 50396 1555 50452
rect 1611 50396 1679 50452
rect 1735 50396 1803 50452
rect 1859 50396 1927 50452
rect 1983 50396 2051 50452
rect 2107 50396 2117 50452
rect 305 50328 2117 50396
rect 305 50272 315 50328
rect 371 50272 439 50328
rect 495 50272 563 50328
rect 619 50272 687 50328
rect 743 50272 811 50328
rect 867 50272 935 50328
rect 991 50272 1059 50328
rect 1115 50272 1183 50328
rect 1239 50272 1307 50328
rect 1363 50272 1431 50328
rect 1487 50272 1555 50328
rect 1611 50272 1679 50328
rect 1735 50272 1803 50328
rect 1859 50272 1927 50328
rect 1983 50272 2051 50328
rect 2107 50272 2117 50328
rect 305 50204 2117 50272
rect 305 50148 315 50204
rect 371 50148 439 50204
rect 495 50148 563 50204
rect 619 50148 687 50204
rect 743 50148 811 50204
rect 867 50148 935 50204
rect 991 50148 1059 50204
rect 1115 50148 1183 50204
rect 1239 50148 1307 50204
rect 1363 50148 1431 50204
rect 1487 50148 1555 50204
rect 1611 50148 1679 50204
rect 1735 50148 1803 50204
rect 1859 50148 1927 50204
rect 1983 50148 2051 50204
rect 2107 50148 2117 50204
rect 305 50080 2117 50148
rect 305 50024 315 50080
rect 371 50024 439 50080
rect 495 50024 563 50080
rect 619 50024 687 50080
rect 743 50024 811 50080
rect 867 50024 935 50080
rect 991 50024 1059 50080
rect 1115 50024 1183 50080
rect 1239 50024 1307 50080
rect 1363 50024 1431 50080
rect 1487 50024 1555 50080
rect 1611 50024 1679 50080
rect 1735 50024 1803 50080
rect 1859 50024 1927 50080
rect 1983 50024 2051 50080
rect 2107 50024 2117 50080
rect 305 49956 2117 50024
rect 305 49900 315 49956
rect 371 49900 439 49956
rect 495 49900 563 49956
rect 619 49900 687 49956
rect 743 49900 811 49956
rect 867 49900 935 49956
rect 991 49900 1059 49956
rect 1115 49900 1183 49956
rect 1239 49900 1307 49956
rect 1363 49900 1431 49956
rect 1487 49900 1555 49956
rect 1611 49900 1679 49956
rect 1735 49900 1803 49956
rect 1859 49900 1927 49956
rect 1983 49900 2051 49956
rect 2107 49900 2117 49956
rect 305 49832 2117 49900
rect 305 49776 315 49832
rect 371 49776 439 49832
rect 495 49776 563 49832
rect 619 49776 687 49832
rect 743 49776 811 49832
rect 867 49776 935 49832
rect 991 49776 1059 49832
rect 1115 49776 1183 49832
rect 1239 49776 1307 49832
rect 1363 49776 1431 49832
rect 1487 49776 1555 49832
rect 1611 49776 1679 49832
rect 1735 49776 1803 49832
rect 1859 49776 1927 49832
rect 1983 49776 2051 49832
rect 2107 49776 2117 49832
rect 305 49708 2117 49776
rect 305 49652 315 49708
rect 371 49652 439 49708
rect 495 49652 563 49708
rect 619 49652 687 49708
rect 743 49652 811 49708
rect 867 49652 935 49708
rect 991 49652 1059 49708
rect 1115 49652 1183 49708
rect 1239 49652 1307 49708
rect 1363 49652 1431 49708
rect 1487 49652 1555 49708
rect 1611 49652 1679 49708
rect 1735 49652 1803 49708
rect 1859 49652 1927 49708
rect 1983 49652 2051 49708
rect 2107 49652 2117 49708
rect 305 49642 2117 49652
rect 2798 50948 4734 50958
rect 2798 50892 2808 50948
rect 2864 50892 2932 50948
rect 2988 50892 3056 50948
rect 3112 50892 3180 50948
rect 3236 50892 3304 50948
rect 3360 50892 3428 50948
rect 3484 50892 3552 50948
rect 3608 50892 3676 50948
rect 3732 50892 3800 50948
rect 3856 50892 3924 50948
rect 3980 50892 4048 50948
rect 4104 50892 4172 50948
rect 4228 50892 4296 50948
rect 4352 50892 4420 50948
rect 4476 50892 4544 50948
rect 4600 50892 4668 50948
rect 4724 50892 4734 50948
rect 2798 50824 4734 50892
rect 2798 50768 2808 50824
rect 2864 50768 2932 50824
rect 2988 50768 3056 50824
rect 3112 50768 3180 50824
rect 3236 50768 3304 50824
rect 3360 50768 3428 50824
rect 3484 50768 3552 50824
rect 3608 50768 3676 50824
rect 3732 50768 3800 50824
rect 3856 50768 3924 50824
rect 3980 50768 4048 50824
rect 4104 50768 4172 50824
rect 4228 50768 4296 50824
rect 4352 50768 4420 50824
rect 4476 50768 4544 50824
rect 4600 50768 4668 50824
rect 4724 50768 4734 50824
rect 2798 50700 4734 50768
rect 2798 50644 2808 50700
rect 2864 50644 2932 50700
rect 2988 50644 3056 50700
rect 3112 50644 3180 50700
rect 3236 50644 3304 50700
rect 3360 50644 3428 50700
rect 3484 50644 3552 50700
rect 3608 50644 3676 50700
rect 3732 50644 3800 50700
rect 3856 50644 3924 50700
rect 3980 50644 4048 50700
rect 4104 50644 4172 50700
rect 4228 50644 4296 50700
rect 4352 50644 4420 50700
rect 4476 50644 4544 50700
rect 4600 50644 4668 50700
rect 4724 50644 4734 50700
rect 2798 50576 4734 50644
rect 2798 50520 2808 50576
rect 2864 50520 2932 50576
rect 2988 50520 3056 50576
rect 3112 50520 3180 50576
rect 3236 50520 3304 50576
rect 3360 50520 3428 50576
rect 3484 50520 3552 50576
rect 3608 50520 3676 50576
rect 3732 50520 3800 50576
rect 3856 50520 3924 50576
rect 3980 50520 4048 50576
rect 4104 50520 4172 50576
rect 4228 50520 4296 50576
rect 4352 50520 4420 50576
rect 4476 50520 4544 50576
rect 4600 50520 4668 50576
rect 4724 50520 4734 50576
rect 2798 50452 4734 50520
rect 2798 50396 2808 50452
rect 2864 50396 2932 50452
rect 2988 50396 3056 50452
rect 3112 50396 3180 50452
rect 3236 50396 3304 50452
rect 3360 50396 3428 50452
rect 3484 50396 3552 50452
rect 3608 50396 3676 50452
rect 3732 50396 3800 50452
rect 3856 50396 3924 50452
rect 3980 50396 4048 50452
rect 4104 50396 4172 50452
rect 4228 50396 4296 50452
rect 4352 50396 4420 50452
rect 4476 50396 4544 50452
rect 4600 50396 4668 50452
rect 4724 50396 4734 50452
rect 2798 50328 4734 50396
rect 2798 50272 2808 50328
rect 2864 50272 2932 50328
rect 2988 50272 3056 50328
rect 3112 50272 3180 50328
rect 3236 50272 3304 50328
rect 3360 50272 3428 50328
rect 3484 50272 3552 50328
rect 3608 50272 3676 50328
rect 3732 50272 3800 50328
rect 3856 50272 3924 50328
rect 3980 50272 4048 50328
rect 4104 50272 4172 50328
rect 4228 50272 4296 50328
rect 4352 50272 4420 50328
rect 4476 50272 4544 50328
rect 4600 50272 4668 50328
rect 4724 50272 4734 50328
rect 2798 50204 4734 50272
rect 2798 50148 2808 50204
rect 2864 50148 2932 50204
rect 2988 50148 3056 50204
rect 3112 50148 3180 50204
rect 3236 50148 3304 50204
rect 3360 50148 3428 50204
rect 3484 50148 3552 50204
rect 3608 50148 3676 50204
rect 3732 50148 3800 50204
rect 3856 50148 3924 50204
rect 3980 50148 4048 50204
rect 4104 50148 4172 50204
rect 4228 50148 4296 50204
rect 4352 50148 4420 50204
rect 4476 50148 4544 50204
rect 4600 50148 4668 50204
rect 4724 50148 4734 50204
rect 2798 50080 4734 50148
rect 2798 50024 2808 50080
rect 2864 50024 2932 50080
rect 2988 50024 3056 50080
rect 3112 50024 3180 50080
rect 3236 50024 3304 50080
rect 3360 50024 3428 50080
rect 3484 50024 3552 50080
rect 3608 50024 3676 50080
rect 3732 50024 3800 50080
rect 3856 50024 3924 50080
rect 3980 50024 4048 50080
rect 4104 50024 4172 50080
rect 4228 50024 4296 50080
rect 4352 50024 4420 50080
rect 4476 50024 4544 50080
rect 4600 50024 4668 50080
rect 4724 50024 4734 50080
rect 2798 49956 4734 50024
rect 2798 49900 2808 49956
rect 2864 49900 2932 49956
rect 2988 49900 3056 49956
rect 3112 49900 3180 49956
rect 3236 49900 3304 49956
rect 3360 49900 3428 49956
rect 3484 49900 3552 49956
rect 3608 49900 3676 49956
rect 3732 49900 3800 49956
rect 3856 49900 3924 49956
rect 3980 49900 4048 49956
rect 4104 49900 4172 49956
rect 4228 49900 4296 49956
rect 4352 49900 4420 49956
rect 4476 49900 4544 49956
rect 4600 49900 4668 49956
rect 4724 49900 4734 49956
rect 2798 49832 4734 49900
rect 2798 49776 2808 49832
rect 2864 49776 2932 49832
rect 2988 49776 3056 49832
rect 3112 49776 3180 49832
rect 3236 49776 3304 49832
rect 3360 49776 3428 49832
rect 3484 49776 3552 49832
rect 3608 49776 3676 49832
rect 3732 49776 3800 49832
rect 3856 49776 3924 49832
rect 3980 49776 4048 49832
rect 4104 49776 4172 49832
rect 4228 49776 4296 49832
rect 4352 49776 4420 49832
rect 4476 49776 4544 49832
rect 4600 49776 4668 49832
rect 4724 49776 4734 49832
rect 2798 49708 4734 49776
rect 2798 49652 2808 49708
rect 2864 49652 2932 49708
rect 2988 49652 3056 49708
rect 3112 49652 3180 49708
rect 3236 49652 3304 49708
rect 3360 49652 3428 49708
rect 3484 49652 3552 49708
rect 3608 49652 3676 49708
rect 3732 49652 3800 49708
rect 3856 49652 3924 49708
rect 3980 49652 4048 49708
rect 4104 49652 4172 49708
rect 4228 49652 4296 49708
rect 4352 49652 4420 49708
rect 4476 49652 4544 49708
rect 4600 49652 4668 49708
rect 4724 49652 4734 49708
rect 2798 49642 4734 49652
rect 5168 50948 7104 50958
rect 5168 50892 5178 50948
rect 5234 50892 5302 50948
rect 5358 50892 5426 50948
rect 5482 50892 5550 50948
rect 5606 50892 5674 50948
rect 5730 50892 5798 50948
rect 5854 50892 5922 50948
rect 5978 50892 6046 50948
rect 6102 50892 6170 50948
rect 6226 50892 6294 50948
rect 6350 50892 6418 50948
rect 6474 50892 6542 50948
rect 6598 50892 6666 50948
rect 6722 50892 6790 50948
rect 6846 50892 6914 50948
rect 6970 50892 7038 50948
rect 7094 50892 7104 50948
rect 5168 50824 7104 50892
rect 5168 50768 5178 50824
rect 5234 50768 5302 50824
rect 5358 50768 5426 50824
rect 5482 50768 5550 50824
rect 5606 50768 5674 50824
rect 5730 50768 5798 50824
rect 5854 50768 5922 50824
rect 5978 50768 6046 50824
rect 6102 50768 6170 50824
rect 6226 50768 6294 50824
rect 6350 50768 6418 50824
rect 6474 50768 6542 50824
rect 6598 50768 6666 50824
rect 6722 50768 6790 50824
rect 6846 50768 6914 50824
rect 6970 50768 7038 50824
rect 7094 50768 7104 50824
rect 5168 50700 7104 50768
rect 5168 50644 5178 50700
rect 5234 50644 5302 50700
rect 5358 50644 5426 50700
rect 5482 50644 5550 50700
rect 5606 50644 5674 50700
rect 5730 50644 5798 50700
rect 5854 50644 5922 50700
rect 5978 50644 6046 50700
rect 6102 50644 6170 50700
rect 6226 50644 6294 50700
rect 6350 50644 6418 50700
rect 6474 50644 6542 50700
rect 6598 50644 6666 50700
rect 6722 50644 6790 50700
rect 6846 50644 6914 50700
rect 6970 50644 7038 50700
rect 7094 50644 7104 50700
rect 5168 50576 7104 50644
rect 5168 50520 5178 50576
rect 5234 50520 5302 50576
rect 5358 50520 5426 50576
rect 5482 50520 5550 50576
rect 5606 50520 5674 50576
rect 5730 50520 5798 50576
rect 5854 50520 5922 50576
rect 5978 50520 6046 50576
rect 6102 50520 6170 50576
rect 6226 50520 6294 50576
rect 6350 50520 6418 50576
rect 6474 50520 6542 50576
rect 6598 50520 6666 50576
rect 6722 50520 6790 50576
rect 6846 50520 6914 50576
rect 6970 50520 7038 50576
rect 7094 50520 7104 50576
rect 5168 50452 7104 50520
rect 5168 50396 5178 50452
rect 5234 50396 5302 50452
rect 5358 50396 5426 50452
rect 5482 50396 5550 50452
rect 5606 50396 5674 50452
rect 5730 50396 5798 50452
rect 5854 50396 5922 50452
rect 5978 50396 6046 50452
rect 6102 50396 6170 50452
rect 6226 50396 6294 50452
rect 6350 50396 6418 50452
rect 6474 50396 6542 50452
rect 6598 50396 6666 50452
rect 6722 50396 6790 50452
rect 6846 50396 6914 50452
rect 6970 50396 7038 50452
rect 7094 50396 7104 50452
rect 5168 50328 7104 50396
rect 5168 50272 5178 50328
rect 5234 50272 5302 50328
rect 5358 50272 5426 50328
rect 5482 50272 5550 50328
rect 5606 50272 5674 50328
rect 5730 50272 5798 50328
rect 5854 50272 5922 50328
rect 5978 50272 6046 50328
rect 6102 50272 6170 50328
rect 6226 50272 6294 50328
rect 6350 50272 6418 50328
rect 6474 50272 6542 50328
rect 6598 50272 6666 50328
rect 6722 50272 6790 50328
rect 6846 50272 6914 50328
rect 6970 50272 7038 50328
rect 7094 50272 7104 50328
rect 5168 50204 7104 50272
rect 5168 50148 5178 50204
rect 5234 50148 5302 50204
rect 5358 50148 5426 50204
rect 5482 50148 5550 50204
rect 5606 50148 5674 50204
rect 5730 50148 5798 50204
rect 5854 50148 5922 50204
rect 5978 50148 6046 50204
rect 6102 50148 6170 50204
rect 6226 50148 6294 50204
rect 6350 50148 6418 50204
rect 6474 50148 6542 50204
rect 6598 50148 6666 50204
rect 6722 50148 6790 50204
rect 6846 50148 6914 50204
rect 6970 50148 7038 50204
rect 7094 50148 7104 50204
rect 5168 50080 7104 50148
rect 5168 50024 5178 50080
rect 5234 50024 5302 50080
rect 5358 50024 5426 50080
rect 5482 50024 5550 50080
rect 5606 50024 5674 50080
rect 5730 50024 5798 50080
rect 5854 50024 5922 50080
rect 5978 50024 6046 50080
rect 6102 50024 6170 50080
rect 6226 50024 6294 50080
rect 6350 50024 6418 50080
rect 6474 50024 6542 50080
rect 6598 50024 6666 50080
rect 6722 50024 6790 50080
rect 6846 50024 6914 50080
rect 6970 50024 7038 50080
rect 7094 50024 7104 50080
rect 5168 49956 7104 50024
rect 5168 49900 5178 49956
rect 5234 49900 5302 49956
rect 5358 49900 5426 49956
rect 5482 49900 5550 49956
rect 5606 49900 5674 49956
rect 5730 49900 5798 49956
rect 5854 49900 5922 49956
rect 5978 49900 6046 49956
rect 6102 49900 6170 49956
rect 6226 49900 6294 49956
rect 6350 49900 6418 49956
rect 6474 49900 6542 49956
rect 6598 49900 6666 49956
rect 6722 49900 6790 49956
rect 6846 49900 6914 49956
rect 6970 49900 7038 49956
rect 7094 49900 7104 49956
rect 5168 49832 7104 49900
rect 5168 49776 5178 49832
rect 5234 49776 5302 49832
rect 5358 49776 5426 49832
rect 5482 49776 5550 49832
rect 5606 49776 5674 49832
rect 5730 49776 5798 49832
rect 5854 49776 5922 49832
rect 5978 49776 6046 49832
rect 6102 49776 6170 49832
rect 6226 49776 6294 49832
rect 6350 49776 6418 49832
rect 6474 49776 6542 49832
rect 6598 49776 6666 49832
rect 6722 49776 6790 49832
rect 6846 49776 6914 49832
rect 6970 49776 7038 49832
rect 7094 49776 7104 49832
rect 5168 49708 7104 49776
rect 5168 49652 5178 49708
rect 5234 49652 5302 49708
rect 5358 49652 5426 49708
rect 5482 49652 5550 49708
rect 5606 49652 5674 49708
rect 5730 49652 5798 49708
rect 5854 49652 5922 49708
rect 5978 49652 6046 49708
rect 6102 49652 6170 49708
rect 6226 49652 6294 49708
rect 6350 49652 6418 49708
rect 6474 49652 6542 49708
rect 6598 49652 6666 49708
rect 6722 49652 6790 49708
rect 6846 49652 6914 49708
rect 6970 49652 7038 49708
rect 7094 49652 7104 49708
rect 5168 49642 7104 49652
rect 7874 50948 9810 50958
rect 7874 50892 7884 50948
rect 7940 50892 8008 50948
rect 8064 50892 8132 50948
rect 8188 50892 8256 50948
rect 8312 50892 8380 50948
rect 8436 50892 8504 50948
rect 8560 50892 8628 50948
rect 8684 50892 8752 50948
rect 8808 50892 8876 50948
rect 8932 50892 9000 50948
rect 9056 50892 9124 50948
rect 9180 50892 9248 50948
rect 9304 50892 9372 50948
rect 9428 50892 9496 50948
rect 9552 50892 9620 50948
rect 9676 50892 9744 50948
rect 9800 50892 9810 50948
rect 7874 50824 9810 50892
rect 7874 50768 7884 50824
rect 7940 50768 8008 50824
rect 8064 50768 8132 50824
rect 8188 50768 8256 50824
rect 8312 50768 8380 50824
rect 8436 50768 8504 50824
rect 8560 50768 8628 50824
rect 8684 50768 8752 50824
rect 8808 50768 8876 50824
rect 8932 50768 9000 50824
rect 9056 50768 9124 50824
rect 9180 50768 9248 50824
rect 9304 50768 9372 50824
rect 9428 50768 9496 50824
rect 9552 50768 9620 50824
rect 9676 50768 9744 50824
rect 9800 50768 9810 50824
rect 7874 50700 9810 50768
rect 7874 50644 7884 50700
rect 7940 50644 8008 50700
rect 8064 50644 8132 50700
rect 8188 50644 8256 50700
rect 8312 50644 8380 50700
rect 8436 50644 8504 50700
rect 8560 50644 8628 50700
rect 8684 50644 8752 50700
rect 8808 50644 8876 50700
rect 8932 50644 9000 50700
rect 9056 50644 9124 50700
rect 9180 50644 9248 50700
rect 9304 50644 9372 50700
rect 9428 50644 9496 50700
rect 9552 50644 9620 50700
rect 9676 50644 9744 50700
rect 9800 50644 9810 50700
rect 7874 50576 9810 50644
rect 7874 50520 7884 50576
rect 7940 50520 8008 50576
rect 8064 50520 8132 50576
rect 8188 50520 8256 50576
rect 8312 50520 8380 50576
rect 8436 50520 8504 50576
rect 8560 50520 8628 50576
rect 8684 50520 8752 50576
rect 8808 50520 8876 50576
rect 8932 50520 9000 50576
rect 9056 50520 9124 50576
rect 9180 50520 9248 50576
rect 9304 50520 9372 50576
rect 9428 50520 9496 50576
rect 9552 50520 9620 50576
rect 9676 50520 9744 50576
rect 9800 50520 9810 50576
rect 7874 50452 9810 50520
rect 7874 50396 7884 50452
rect 7940 50396 8008 50452
rect 8064 50396 8132 50452
rect 8188 50396 8256 50452
rect 8312 50396 8380 50452
rect 8436 50396 8504 50452
rect 8560 50396 8628 50452
rect 8684 50396 8752 50452
rect 8808 50396 8876 50452
rect 8932 50396 9000 50452
rect 9056 50396 9124 50452
rect 9180 50396 9248 50452
rect 9304 50396 9372 50452
rect 9428 50396 9496 50452
rect 9552 50396 9620 50452
rect 9676 50396 9744 50452
rect 9800 50396 9810 50452
rect 7874 50328 9810 50396
rect 7874 50272 7884 50328
rect 7940 50272 8008 50328
rect 8064 50272 8132 50328
rect 8188 50272 8256 50328
rect 8312 50272 8380 50328
rect 8436 50272 8504 50328
rect 8560 50272 8628 50328
rect 8684 50272 8752 50328
rect 8808 50272 8876 50328
rect 8932 50272 9000 50328
rect 9056 50272 9124 50328
rect 9180 50272 9248 50328
rect 9304 50272 9372 50328
rect 9428 50272 9496 50328
rect 9552 50272 9620 50328
rect 9676 50272 9744 50328
rect 9800 50272 9810 50328
rect 7874 50204 9810 50272
rect 7874 50148 7884 50204
rect 7940 50148 8008 50204
rect 8064 50148 8132 50204
rect 8188 50148 8256 50204
rect 8312 50148 8380 50204
rect 8436 50148 8504 50204
rect 8560 50148 8628 50204
rect 8684 50148 8752 50204
rect 8808 50148 8876 50204
rect 8932 50148 9000 50204
rect 9056 50148 9124 50204
rect 9180 50148 9248 50204
rect 9304 50148 9372 50204
rect 9428 50148 9496 50204
rect 9552 50148 9620 50204
rect 9676 50148 9744 50204
rect 9800 50148 9810 50204
rect 7874 50080 9810 50148
rect 7874 50024 7884 50080
rect 7940 50024 8008 50080
rect 8064 50024 8132 50080
rect 8188 50024 8256 50080
rect 8312 50024 8380 50080
rect 8436 50024 8504 50080
rect 8560 50024 8628 50080
rect 8684 50024 8752 50080
rect 8808 50024 8876 50080
rect 8932 50024 9000 50080
rect 9056 50024 9124 50080
rect 9180 50024 9248 50080
rect 9304 50024 9372 50080
rect 9428 50024 9496 50080
rect 9552 50024 9620 50080
rect 9676 50024 9744 50080
rect 9800 50024 9810 50080
rect 7874 49956 9810 50024
rect 7874 49900 7884 49956
rect 7940 49900 8008 49956
rect 8064 49900 8132 49956
rect 8188 49900 8256 49956
rect 8312 49900 8380 49956
rect 8436 49900 8504 49956
rect 8560 49900 8628 49956
rect 8684 49900 8752 49956
rect 8808 49900 8876 49956
rect 8932 49900 9000 49956
rect 9056 49900 9124 49956
rect 9180 49900 9248 49956
rect 9304 49900 9372 49956
rect 9428 49900 9496 49956
rect 9552 49900 9620 49956
rect 9676 49900 9744 49956
rect 9800 49900 9810 49956
rect 7874 49832 9810 49900
rect 7874 49776 7884 49832
rect 7940 49776 8008 49832
rect 8064 49776 8132 49832
rect 8188 49776 8256 49832
rect 8312 49776 8380 49832
rect 8436 49776 8504 49832
rect 8560 49776 8628 49832
rect 8684 49776 8752 49832
rect 8808 49776 8876 49832
rect 8932 49776 9000 49832
rect 9056 49776 9124 49832
rect 9180 49776 9248 49832
rect 9304 49776 9372 49832
rect 9428 49776 9496 49832
rect 9552 49776 9620 49832
rect 9676 49776 9744 49832
rect 9800 49776 9810 49832
rect 7874 49708 9810 49776
rect 7874 49652 7884 49708
rect 7940 49652 8008 49708
rect 8064 49652 8132 49708
rect 8188 49652 8256 49708
rect 8312 49652 8380 49708
rect 8436 49652 8504 49708
rect 8560 49652 8628 49708
rect 8684 49652 8752 49708
rect 8808 49652 8876 49708
rect 8932 49652 9000 49708
rect 9056 49652 9124 49708
rect 9180 49652 9248 49708
rect 9304 49652 9372 49708
rect 9428 49652 9496 49708
rect 9552 49652 9620 49708
rect 9676 49652 9744 49708
rect 9800 49652 9810 49708
rect 7874 49642 9810 49652
rect 10244 50948 12180 50958
rect 10244 50892 10254 50948
rect 10310 50892 10378 50948
rect 10434 50892 10502 50948
rect 10558 50892 10626 50948
rect 10682 50892 10750 50948
rect 10806 50892 10874 50948
rect 10930 50892 10998 50948
rect 11054 50892 11122 50948
rect 11178 50892 11246 50948
rect 11302 50892 11370 50948
rect 11426 50892 11494 50948
rect 11550 50892 11618 50948
rect 11674 50892 11742 50948
rect 11798 50892 11866 50948
rect 11922 50892 11990 50948
rect 12046 50892 12114 50948
rect 12170 50892 12180 50948
rect 10244 50824 12180 50892
rect 10244 50768 10254 50824
rect 10310 50768 10378 50824
rect 10434 50768 10502 50824
rect 10558 50768 10626 50824
rect 10682 50768 10750 50824
rect 10806 50768 10874 50824
rect 10930 50768 10998 50824
rect 11054 50768 11122 50824
rect 11178 50768 11246 50824
rect 11302 50768 11370 50824
rect 11426 50768 11494 50824
rect 11550 50768 11618 50824
rect 11674 50768 11742 50824
rect 11798 50768 11866 50824
rect 11922 50768 11990 50824
rect 12046 50768 12114 50824
rect 12170 50768 12180 50824
rect 10244 50700 12180 50768
rect 10244 50644 10254 50700
rect 10310 50644 10378 50700
rect 10434 50644 10502 50700
rect 10558 50644 10626 50700
rect 10682 50644 10750 50700
rect 10806 50644 10874 50700
rect 10930 50644 10998 50700
rect 11054 50644 11122 50700
rect 11178 50644 11246 50700
rect 11302 50644 11370 50700
rect 11426 50644 11494 50700
rect 11550 50644 11618 50700
rect 11674 50644 11742 50700
rect 11798 50644 11866 50700
rect 11922 50644 11990 50700
rect 12046 50644 12114 50700
rect 12170 50644 12180 50700
rect 10244 50576 12180 50644
rect 10244 50520 10254 50576
rect 10310 50520 10378 50576
rect 10434 50520 10502 50576
rect 10558 50520 10626 50576
rect 10682 50520 10750 50576
rect 10806 50520 10874 50576
rect 10930 50520 10998 50576
rect 11054 50520 11122 50576
rect 11178 50520 11246 50576
rect 11302 50520 11370 50576
rect 11426 50520 11494 50576
rect 11550 50520 11618 50576
rect 11674 50520 11742 50576
rect 11798 50520 11866 50576
rect 11922 50520 11990 50576
rect 12046 50520 12114 50576
rect 12170 50520 12180 50576
rect 10244 50452 12180 50520
rect 10244 50396 10254 50452
rect 10310 50396 10378 50452
rect 10434 50396 10502 50452
rect 10558 50396 10626 50452
rect 10682 50396 10750 50452
rect 10806 50396 10874 50452
rect 10930 50396 10998 50452
rect 11054 50396 11122 50452
rect 11178 50396 11246 50452
rect 11302 50396 11370 50452
rect 11426 50396 11494 50452
rect 11550 50396 11618 50452
rect 11674 50396 11742 50452
rect 11798 50396 11866 50452
rect 11922 50396 11990 50452
rect 12046 50396 12114 50452
rect 12170 50396 12180 50452
rect 10244 50328 12180 50396
rect 10244 50272 10254 50328
rect 10310 50272 10378 50328
rect 10434 50272 10502 50328
rect 10558 50272 10626 50328
rect 10682 50272 10750 50328
rect 10806 50272 10874 50328
rect 10930 50272 10998 50328
rect 11054 50272 11122 50328
rect 11178 50272 11246 50328
rect 11302 50272 11370 50328
rect 11426 50272 11494 50328
rect 11550 50272 11618 50328
rect 11674 50272 11742 50328
rect 11798 50272 11866 50328
rect 11922 50272 11990 50328
rect 12046 50272 12114 50328
rect 12170 50272 12180 50328
rect 10244 50204 12180 50272
rect 10244 50148 10254 50204
rect 10310 50148 10378 50204
rect 10434 50148 10502 50204
rect 10558 50148 10626 50204
rect 10682 50148 10750 50204
rect 10806 50148 10874 50204
rect 10930 50148 10998 50204
rect 11054 50148 11122 50204
rect 11178 50148 11246 50204
rect 11302 50148 11370 50204
rect 11426 50148 11494 50204
rect 11550 50148 11618 50204
rect 11674 50148 11742 50204
rect 11798 50148 11866 50204
rect 11922 50148 11990 50204
rect 12046 50148 12114 50204
rect 12170 50148 12180 50204
rect 10244 50080 12180 50148
rect 10244 50024 10254 50080
rect 10310 50024 10378 50080
rect 10434 50024 10502 50080
rect 10558 50024 10626 50080
rect 10682 50024 10750 50080
rect 10806 50024 10874 50080
rect 10930 50024 10998 50080
rect 11054 50024 11122 50080
rect 11178 50024 11246 50080
rect 11302 50024 11370 50080
rect 11426 50024 11494 50080
rect 11550 50024 11618 50080
rect 11674 50024 11742 50080
rect 11798 50024 11866 50080
rect 11922 50024 11990 50080
rect 12046 50024 12114 50080
rect 12170 50024 12180 50080
rect 10244 49956 12180 50024
rect 10244 49900 10254 49956
rect 10310 49900 10378 49956
rect 10434 49900 10502 49956
rect 10558 49900 10626 49956
rect 10682 49900 10750 49956
rect 10806 49900 10874 49956
rect 10930 49900 10998 49956
rect 11054 49900 11122 49956
rect 11178 49900 11246 49956
rect 11302 49900 11370 49956
rect 11426 49900 11494 49956
rect 11550 49900 11618 49956
rect 11674 49900 11742 49956
rect 11798 49900 11866 49956
rect 11922 49900 11990 49956
rect 12046 49900 12114 49956
rect 12170 49900 12180 49956
rect 10244 49832 12180 49900
rect 10244 49776 10254 49832
rect 10310 49776 10378 49832
rect 10434 49776 10502 49832
rect 10558 49776 10626 49832
rect 10682 49776 10750 49832
rect 10806 49776 10874 49832
rect 10930 49776 10998 49832
rect 11054 49776 11122 49832
rect 11178 49776 11246 49832
rect 11302 49776 11370 49832
rect 11426 49776 11494 49832
rect 11550 49776 11618 49832
rect 11674 49776 11742 49832
rect 11798 49776 11866 49832
rect 11922 49776 11990 49832
rect 12046 49776 12114 49832
rect 12170 49776 12180 49832
rect 10244 49708 12180 49776
rect 10244 49652 10254 49708
rect 10310 49652 10378 49708
rect 10434 49652 10502 49708
rect 10558 49652 10626 49708
rect 10682 49652 10750 49708
rect 10806 49652 10874 49708
rect 10930 49652 10998 49708
rect 11054 49652 11122 49708
rect 11178 49652 11246 49708
rect 11302 49652 11370 49708
rect 11426 49652 11494 49708
rect 11550 49652 11618 49708
rect 11674 49652 11742 49708
rect 11798 49652 11866 49708
rect 11922 49652 11990 49708
rect 12046 49652 12114 49708
rect 12170 49652 12180 49708
rect 10244 49642 12180 49652
rect 12861 50948 14673 50958
rect 12861 50892 12871 50948
rect 12927 50892 12995 50948
rect 13051 50892 13119 50948
rect 13175 50892 13243 50948
rect 13299 50892 13367 50948
rect 13423 50892 13491 50948
rect 13547 50892 13615 50948
rect 13671 50892 13739 50948
rect 13795 50892 13863 50948
rect 13919 50892 13987 50948
rect 14043 50892 14111 50948
rect 14167 50892 14235 50948
rect 14291 50892 14359 50948
rect 14415 50892 14483 50948
rect 14539 50892 14607 50948
rect 14663 50892 14673 50948
rect 12861 50824 14673 50892
rect 12861 50768 12871 50824
rect 12927 50768 12995 50824
rect 13051 50768 13119 50824
rect 13175 50768 13243 50824
rect 13299 50768 13367 50824
rect 13423 50768 13491 50824
rect 13547 50768 13615 50824
rect 13671 50768 13739 50824
rect 13795 50768 13863 50824
rect 13919 50768 13987 50824
rect 14043 50768 14111 50824
rect 14167 50768 14235 50824
rect 14291 50768 14359 50824
rect 14415 50768 14483 50824
rect 14539 50768 14607 50824
rect 14663 50768 14673 50824
rect 12861 50700 14673 50768
rect 12861 50644 12871 50700
rect 12927 50644 12995 50700
rect 13051 50644 13119 50700
rect 13175 50644 13243 50700
rect 13299 50644 13367 50700
rect 13423 50644 13491 50700
rect 13547 50644 13615 50700
rect 13671 50644 13739 50700
rect 13795 50644 13863 50700
rect 13919 50644 13987 50700
rect 14043 50644 14111 50700
rect 14167 50644 14235 50700
rect 14291 50644 14359 50700
rect 14415 50644 14483 50700
rect 14539 50644 14607 50700
rect 14663 50644 14673 50700
rect 12861 50576 14673 50644
rect 12861 50520 12871 50576
rect 12927 50520 12995 50576
rect 13051 50520 13119 50576
rect 13175 50520 13243 50576
rect 13299 50520 13367 50576
rect 13423 50520 13491 50576
rect 13547 50520 13615 50576
rect 13671 50520 13739 50576
rect 13795 50520 13863 50576
rect 13919 50520 13987 50576
rect 14043 50520 14111 50576
rect 14167 50520 14235 50576
rect 14291 50520 14359 50576
rect 14415 50520 14483 50576
rect 14539 50520 14607 50576
rect 14663 50520 14673 50576
rect 12861 50452 14673 50520
rect 12861 50396 12871 50452
rect 12927 50396 12995 50452
rect 13051 50396 13119 50452
rect 13175 50396 13243 50452
rect 13299 50396 13367 50452
rect 13423 50396 13491 50452
rect 13547 50396 13615 50452
rect 13671 50396 13739 50452
rect 13795 50396 13863 50452
rect 13919 50396 13987 50452
rect 14043 50396 14111 50452
rect 14167 50396 14235 50452
rect 14291 50396 14359 50452
rect 14415 50396 14483 50452
rect 14539 50396 14607 50452
rect 14663 50396 14673 50452
rect 12861 50328 14673 50396
rect 12861 50272 12871 50328
rect 12927 50272 12995 50328
rect 13051 50272 13119 50328
rect 13175 50272 13243 50328
rect 13299 50272 13367 50328
rect 13423 50272 13491 50328
rect 13547 50272 13615 50328
rect 13671 50272 13739 50328
rect 13795 50272 13863 50328
rect 13919 50272 13987 50328
rect 14043 50272 14111 50328
rect 14167 50272 14235 50328
rect 14291 50272 14359 50328
rect 14415 50272 14483 50328
rect 14539 50272 14607 50328
rect 14663 50272 14673 50328
rect 12861 50204 14673 50272
rect 12861 50148 12871 50204
rect 12927 50148 12995 50204
rect 13051 50148 13119 50204
rect 13175 50148 13243 50204
rect 13299 50148 13367 50204
rect 13423 50148 13491 50204
rect 13547 50148 13615 50204
rect 13671 50148 13739 50204
rect 13795 50148 13863 50204
rect 13919 50148 13987 50204
rect 14043 50148 14111 50204
rect 14167 50148 14235 50204
rect 14291 50148 14359 50204
rect 14415 50148 14483 50204
rect 14539 50148 14607 50204
rect 14663 50148 14673 50204
rect 12861 50080 14673 50148
rect 12861 50024 12871 50080
rect 12927 50024 12995 50080
rect 13051 50024 13119 50080
rect 13175 50024 13243 50080
rect 13299 50024 13367 50080
rect 13423 50024 13491 50080
rect 13547 50024 13615 50080
rect 13671 50024 13739 50080
rect 13795 50024 13863 50080
rect 13919 50024 13987 50080
rect 14043 50024 14111 50080
rect 14167 50024 14235 50080
rect 14291 50024 14359 50080
rect 14415 50024 14483 50080
rect 14539 50024 14607 50080
rect 14663 50024 14673 50080
rect 12861 49956 14673 50024
rect 12861 49900 12871 49956
rect 12927 49900 12995 49956
rect 13051 49900 13119 49956
rect 13175 49900 13243 49956
rect 13299 49900 13367 49956
rect 13423 49900 13491 49956
rect 13547 49900 13615 49956
rect 13671 49900 13739 49956
rect 13795 49900 13863 49956
rect 13919 49900 13987 49956
rect 14043 49900 14111 49956
rect 14167 49900 14235 49956
rect 14291 49900 14359 49956
rect 14415 49900 14483 49956
rect 14539 49900 14607 49956
rect 14663 49900 14673 49956
rect 12861 49832 14673 49900
rect 12861 49776 12871 49832
rect 12927 49776 12995 49832
rect 13051 49776 13119 49832
rect 13175 49776 13243 49832
rect 13299 49776 13367 49832
rect 13423 49776 13491 49832
rect 13547 49776 13615 49832
rect 13671 49776 13739 49832
rect 13795 49776 13863 49832
rect 13919 49776 13987 49832
rect 14043 49776 14111 49832
rect 14167 49776 14235 49832
rect 14291 49776 14359 49832
rect 14415 49776 14483 49832
rect 14539 49776 14607 49832
rect 14663 49776 14673 49832
rect 12861 49708 14673 49776
rect 12861 49652 12871 49708
rect 12927 49652 12995 49708
rect 13051 49652 13119 49708
rect 13175 49652 13243 49708
rect 13299 49652 13367 49708
rect 13423 49652 13491 49708
rect 13547 49652 13615 49708
rect 13671 49652 13739 49708
rect 13795 49652 13863 49708
rect 13919 49652 13987 49708
rect 14043 49652 14111 49708
rect 14167 49652 14235 49708
rect 14291 49652 14359 49708
rect 14415 49652 14483 49708
rect 14539 49652 14607 49708
rect 14663 49652 14673 49708
rect 12861 49642 14673 49652
rect 2481 49348 2681 49358
rect 2481 49292 2491 49348
rect 2547 49292 2615 49348
rect 2671 49292 2681 49348
rect 2481 49224 2681 49292
rect 2481 49168 2491 49224
rect 2547 49168 2615 49224
rect 2671 49168 2681 49224
rect 2481 49100 2681 49168
rect 2481 49044 2491 49100
rect 2547 49044 2615 49100
rect 2671 49044 2681 49100
rect 2481 48976 2681 49044
rect 2481 48920 2491 48976
rect 2547 48920 2615 48976
rect 2671 48920 2681 48976
rect 2481 48852 2681 48920
rect 2481 48796 2491 48852
rect 2547 48796 2615 48852
rect 2671 48796 2681 48852
rect 2481 48728 2681 48796
rect 2481 48672 2491 48728
rect 2547 48672 2615 48728
rect 2671 48672 2681 48728
rect 2481 48604 2681 48672
rect 2481 48548 2491 48604
rect 2547 48548 2615 48604
rect 2671 48548 2681 48604
rect 2481 48480 2681 48548
rect 2481 48424 2491 48480
rect 2547 48424 2615 48480
rect 2671 48424 2681 48480
rect 2481 48356 2681 48424
rect 2481 48300 2491 48356
rect 2547 48300 2615 48356
rect 2671 48300 2681 48356
rect 2481 48232 2681 48300
rect 2481 48176 2491 48232
rect 2547 48176 2615 48232
rect 2671 48176 2681 48232
rect 2481 48108 2681 48176
rect 2481 48052 2491 48108
rect 2547 48052 2615 48108
rect 2671 48052 2681 48108
rect 2481 48042 2681 48052
rect 4851 49348 5051 49358
rect 4851 49292 4861 49348
rect 4917 49292 4985 49348
rect 5041 49292 5051 49348
rect 4851 49224 5051 49292
rect 4851 49168 4861 49224
rect 4917 49168 4985 49224
rect 5041 49168 5051 49224
rect 4851 49100 5051 49168
rect 4851 49044 4861 49100
rect 4917 49044 4985 49100
rect 5041 49044 5051 49100
rect 4851 48976 5051 49044
rect 4851 48920 4861 48976
rect 4917 48920 4985 48976
rect 5041 48920 5051 48976
rect 4851 48852 5051 48920
rect 4851 48796 4861 48852
rect 4917 48796 4985 48852
rect 5041 48796 5051 48852
rect 4851 48728 5051 48796
rect 4851 48672 4861 48728
rect 4917 48672 4985 48728
rect 5041 48672 5051 48728
rect 4851 48604 5051 48672
rect 4851 48548 4861 48604
rect 4917 48548 4985 48604
rect 5041 48548 5051 48604
rect 4851 48480 5051 48548
rect 4851 48424 4861 48480
rect 4917 48424 4985 48480
rect 5041 48424 5051 48480
rect 4851 48356 5051 48424
rect 4851 48300 4861 48356
rect 4917 48300 4985 48356
rect 5041 48300 5051 48356
rect 4851 48232 5051 48300
rect 4851 48176 4861 48232
rect 4917 48176 4985 48232
rect 5041 48176 5051 48232
rect 4851 48108 5051 48176
rect 4851 48052 4861 48108
rect 4917 48052 4985 48108
rect 5041 48052 5051 48108
rect 4851 48042 5051 48052
rect 7265 49348 7713 49358
rect 7265 49292 7275 49348
rect 7331 49292 7399 49348
rect 7455 49292 7523 49348
rect 7579 49292 7647 49348
rect 7703 49292 7713 49348
rect 7265 49224 7713 49292
rect 7265 49168 7275 49224
rect 7331 49168 7399 49224
rect 7455 49168 7523 49224
rect 7579 49168 7647 49224
rect 7703 49168 7713 49224
rect 7265 49100 7713 49168
rect 7265 49044 7275 49100
rect 7331 49044 7399 49100
rect 7455 49044 7523 49100
rect 7579 49044 7647 49100
rect 7703 49044 7713 49100
rect 7265 48976 7713 49044
rect 7265 48920 7275 48976
rect 7331 48920 7399 48976
rect 7455 48920 7523 48976
rect 7579 48920 7647 48976
rect 7703 48920 7713 48976
rect 7265 48852 7713 48920
rect 7265 48796 7275 48852
rect 7331 48796 7399 48852
rect 7455 48796 7523 48852
rect 7579 48796 7647 48852
rect 7703 48796 7713 48852
rect 7265 48728 7713 48796
rect 7265 48672 7275 48728
rect 7331 48672 7399 48728
rect 7455 48672 7523 48728
rect 7579 48672 7647 48728
rect 7703 48672 7713 48728
rect 7265 48604 7713 48672
rect 7265 48548 7275 48604
rect 7331 48548 7399 48604
rect 7455 48548 7523 48604
rect 7579 48548 7647 48604
rect 7703 48548 7713 48604
rect 7265 48480 7713 48548
rect 7265 48424 7275 48480
rect 7331 48424 7399 48480
rect 7455 48424 7523 48480
rect 7579 48424 7647 48480
rect 7703 48424 7713 48480
rect 7265 48356 7713 48424
rect 7265 48300 7275 48356
rect 7331 48300 7399 48356
rect 7455 48300 7523 48356
rect 7579 48300 7647 48356
rect 7703 48300 7713 48356
rect 7265 48232 7713 48300
rect 7265 48176 7275 48232
rect 7331 48176 7399 48232
rect 7455 48176 7523 48232
rect 7579 48176 7647 48232
rect 7703 48176 7713 48232
rect 7265 48108 7713 48176
rect 7265 48052 7275 48108
rect 7331 48052 7399 48108
rect 7455 48052 7523 48108
rect 7579 48052 7647 48108
rect 7703 48052 7713 48108
rect 7265 48042 7713 48052
rect 9927 49348 10127 49358
rect 9927 49292 9937 49348
rect 9993 49292 10061 49348
rect 10117 49292 10127 49348
rect 9927 49224 10127 49292
rect 9927 49168 9937 49224
rect 9993 49168 10061 49224
rect 10117 49168 10127 49224
rect 9927 49100 10127 49168
rect 9927 49044 9937 49100
rect 9993 49044 10061 49100
rect 10117 49044 10127 49100
rect 9927 48976 10127 49044
rect 9927 48920 9937 48976
rect 9993 48920 10061 48976
rect 10117 48920 10127 48976
rect 9927 48852 10127 48920
rect 9927 48796 9937 48852
rect 9993 48796 10061 48852
rect 10117 48796 10127 48852
rect 9927 48728 10127 48796
rect 9927 48672 9937 48728
rect 9993 48672 10061 48728
rect 10117 48672 10127 48728
rect 9927 48604 10127 48672
rect 9927 48548 9937 48604
rect 9993 48548 10061 48604
rect 10117 48548 10127 48604
rect 9927 48480 10127 48548
rect 9927 48424 9937 48480
rect 9993 48424 10061 48480
rect 10117 48424 10127 48480
rect 9927 48356 10127 48424
rect 9927 48300 9937 48356
rect 9993 48300 10061 48356
rect 10117 48300 10127 48356
rect 9927 48232 10127 48300
rect 9927 48176 9937 48232
rect 9993 48176 10061 48232
rect 10117 48176 10127 48232
rect 9927 48108 10127 48176
rect 9927 48052 9937 48108
rect 9993 48052 10061 48108
rect 10117 48052 10127 48108
rect 9927 48042 10127 48052
rect 12297 49348 12497 49358
rect 12297 49292 12307 49348
rect 12363 49292 12431 49348
rect 12487 49292 12497 49348
rect 12297 49224 12497 49292
rect 12297 49168 12307 49224
rect 12363 49168 12431 49224
rect 12487 49168 12497 49224
rect 12297 49100 12497 49168
rect 12297 49044 12307 49100
rect 12363 49044 12431 49100
rect 12487 49044 12497 49100
rect 12297 48976 12497 49044
rect 12297 48920 12307 48976
rect 12363 48920 12431 48976
rect 12487 48920 12497 48976
rect 12297 48852 12497 48920
rect 12297 48796 12307 48852
rect 12363 48796 12431 48852
rect 12487 48796 12497 48852
rect 12297 48728 12497 48796
rect 12297 48672 12307 48728
rect 12363 48672 12431 48728
rect 12487 48672 12497 48728
rect 12297 48604 12497 48672
rect 12297 48548 12307 48604
rect 12363 48548 12431 48604
rect 12487 48548 12497 48604
rect 12297 48480 12497 48548
rect 12297 48424 12307 48480
rect 12363 48424 12431 48480
rect 12487 48424 12497 48480
rect 12297 48356 12497 48424
rect 12297 48300 12307 48356
rect 12363 48300 12431 48356
rect 12487 48300 12497 48356
rect 12297 48232 12497 48300
rect 12297 48176 12307 48232
rect 12363 48176 12431 48232
rect 12487 48176 12497 48232
rect 12297 48108 12497 48176
rect 12297 48052 12307 48108
rect 12363 48052 12431 48108
rect 12487 48052 12497 48108
rect 12297 48042 12497 48052
rect 305 47748 2117 47758
rect 305 47692 315 47748
rect 371 47692 439 47748
rect 495 47692 563 47748
rect 619 47692 687 47748
rect 743 47692 811 47748
rect 867 47692 935 47748
rect 991 47692 1059 47748
rect 1115 47692 1183 47748
rect 1239 47692 1307 47748
rect 1363 47692 1431 47748
rect 1487 47692 1555 47748
rect 1611 47692 1679 47748
rect 1735 47692 1803 47748
rect 1859 47692 1927 47748
rect 1983 47692 2051 47748
rect 2107 47692 2117 47748
rect 305 47624 2117 47692
rect 305 47568 315 47624
rect 371 47568 439 47624
rect 495 47568 563 47624
rect 619 47568 687 47624
rect 743 47568 811 47624
rect 867 47568 935 47624
rect 991 47568 1059 47624
rect 1115 47568 1183 47624
rect 1239 47568 1307 47624
rect 1363 47568 1431 47624
rect 1487 47568 1555 47624
rect 1611 47568 1679 47624
rect 1735 47568 1803 47624
rect 1859 47568 1927 47624
rect 1983 47568 2051 47624
rect 2107 47568 2117 47624
rect 305 47500 2117 47568
rect 305 47444 315 47500
rect 371 47444 439 47500
rect 495 47444 563 47500
rect 619 47444 687 47500
rect 743 47444 811 47500
rect 867 47444 935 47500
rect 991 47444 1059 47500
rect 1115 47444 1183 47500
rect 1239 47444 1307 47500
rect 1363 47444 1431 47500
rect 1487 47444 1555 47500
rect 1611 47444 1679 47500
rect 1735 47444 1803 47500
rect 1859 47444 1927 47500
rect 1983 47444 2051 47500
rect 2107 47444 2117 47500
rect 305 47376 2117 47444
rect 305 47320 315 47376
rect 371 47320 439 47376
rect 495 47320 563 47376
rect 619 47320 687 47376
rect 743 47320 811 47376
rect 867 47320 935 47376
rect 991 47320 1059 47376
rect 1115 47320 1183 47376
rect 1239 47320 1307 47376
rect 1363 47320 1431 47376
rect 1487 47320 1555 47376
rect 1611 47320 1679 47376
rect 1735 47320 1803 47376
rect 1859 47320 1927 47376
rect 1983 47320 2051 47376
rect 2107 47320 2117 47376
rect 305 47252 2117 47320
rect 305 47196 315 47252
rect 371 47196 439 47252
rect 495 47196 563 47252
rect 619 47196 687 47252
rect 743 47196 811 47252
rect 867 47196 935 47252
rect 991 47196 1059 47252
rect 1115 47196 1183 47252
rect 1239 47196 1307 47252
rect 1363 47196 1431 47252
rect 1487 47196 1555 47252
rect 1611 47196 1679 47252
rect 1735 47196 1803 47252
rect 1859 47196 1927 47252
rect 1983 47196 2051 47252
rect 2107 47196 2117 47252
rect 305 47128 2117 47196
rect 305 47072 315 47128
rect 371 47072 439 47128
rect 495 47072 563 47128
rect 619 47072 687 47128
rect 743 47072 811 47128
rect 867 47072 935 47128
rect 991 47072 1059 47128
rect 1115 47072 1183 47128
rect 1239 47072 1307 47128
rect 1363 47072 1431 47128
rect 1487 47072 1555 47128
rect 1611 47072 1679 47128
rect 1735 47072 1803 47128
rect 1859 47072 1927 47128
rect 1983 47072 2051 47128
rect 2107 47072 2117 47128
rect 305 47004 2117 47072
rect 305 46948 315 47004
rect 371 46948 439 47004
rect 495 46948 563 47004
rect 619 46948 687 47004
rect 743 46948 811 47004
rect 867 46948 935 47004
rect 991 46948 1059 47004
rect 1115 46948 1183 47004
rect 1239 46948 1307 47004
rect 1363 46948 1431 47004
rect 1487 46948 1555 47004
rect 1611 46948 1679 47004
rect 1735 46948 1803 47004
rect 1859 46948 1927 47004
rect 1983 46948 2051 47004
rect 2107 46948 2117 47004
rect 305 46880 2117 46948
rect 305 46824 315 46880
rect 371 46824 439 46880
rect 495 46824 563 46880
rect 619 46824 687 46880
rect 743 46824 811 46880
rect 867 46824 935 46880
rect 991 46824 1059 46880
rect 1115 46824 1183 46880
rect 1239 46824 1307 46880
rect 1363 46824 1431 46880
rect 1487 46824 1555 46880
rect 1611 46824 1679 46880
rect 1735 46824 1803 46880
rect 1859 46824 1927 46880
rect 1983 46824 2051 46880
rect 2107 46824 2117 46880
rect 305 46756 2117 46824
rect 305 46700 315 46756
rect 371 46700 439 46756
rect 495 46700 563 46756
rect 619 46700 687 46756
rect 743 46700 811 46756
rect 867 46700 935 46756
rect 991 46700 1059 46756
rect 1115 46700 1183 46756
rect 1239 46700 1307 46756
rect 1363 46700 1431 46756
rect 1487 46700 1555 46756
rect 1611 46700 1679 46756
rect 1735 46700 1803 46756
rect 1859 46700 1927 46756
rect 1983 46700 2051 46756
rect 2107 46700 2117 46756
rect 305 46632 2117 46700
rect 305 46576 315 46632
rect 371 46576 439 46632
rect 495 46576 563 46632
rect 619 46576 687 46632
rect 743 46576 811 46632
rect 867 46576 935 46632
rect 991 46576 1059 46632
rect 1115 46576 1183 46632
rect 1239 46576 1307 46632
rect 1363 46576 1431 46632
rect 1487 46576 1555 46632
rect 1611 46576 1679 46632
rect 1735 46576 1803 46632
rect 1859 46576 1927 46632
rect 1983 46576 2051 46632
rect 2107 46576 2117 46632
rect 305 46508 2117 46576
rect 305 46452 315 46508
rect 371 46452 439 46508
rect 495 46452 563 46508
rect 619 46452 687 46508
rect 743 46452 811 46508
rect 867 46452 935 46508
rect 991 46452 1059 46508
rect 1115 46452 1183 46508
rect 1239 46452 1307 46508
rect 1363 46452 1431 46508
rect 1487 46452 1555 46508
rect 1611 46452 1679 46508
rect 1735 46452 1803 46508
rect 1859 46452 1927 46508
rect 1983 46452 2051 46508
rect 2107 46452 2117 46508
rect 305 46442 2117 46452
rect 2798 47748 4734 47758
rect 2798 47692 2808 47748
rect 2864 47692 2932 47748
rect 2988 47692 3056 47748
rect 3112 47692 3180 47748
rect 3236 47692 3304 47748
rect 3360 47692 3428 47748
rect 3484 47692 3552 47748
rect 3608 47692 3676 47748
rect 3732 47692 3800 47748
rect 3856 47692 3924 47748
rect 3980 47692 4048 47748
rect 4104 47692 4172 47748
rect 4228 47692 4296 47748
rect 4352 47692 4420 47748
rect 4476 47692 4544 47748
rect 4600 47692 4668 47748
rect 4724 47692 4734 47748
rect 2798 47624 4734 47692
rect 2798 47568 2808 47624
rect 2864 47568 2932 47624
rect 2988 47568 3056 47624
rect 3112 47568 3180 47624
rect 3236 47568 3304 47624
rect 3360 47568 3428 47624
rect 3484 47568 3552 47624
rect 3608 47568 3676 47624
rect 3732 47568 3800 47624
rect 3856 47568 3924 47624
rect 3980 47568 4048 47624
rect 4104 47568 4172 47624
rect 4228 47568 4296 47624
rect 4352 47568 4420 47624
rect 4476 47568 4544 47624
rect 4600 47568 4668 47624
rect 4724 47568 4734 47624
rect 2798 47500 4734 47568
rect 2798 47444 2808 47500
rect 2864 47444 2932 47500
rect 2988 47444 3056 47500
rect 3112 47444 3180 47500
rect 3236 47444 3304 47500
rect 3360 47444 3428 47500
rect 3484 47444 3552 47500
rect 3608 47444 3676 47500
rect 3732 47444 3800 47500
rect 3856 47444 3924 47500
rect 3980 47444 4048 47500
rect 4104 47444 4172 47500
rect 4228 47444 4296 47500
rect 4352 47444 4420 47500
rect 4476 47444 4544 47500
rect 4600 47444 4668 47500
rect 4724 47444 4734 47500
rect 2798 47376 4734 47444
rect 2798 47320 2808 47376
rect 2864 47320 2932 47376
rect 2988 47320 3056 47376
rect 3112 47320 3180 47376
rect 3236 47320 3304 47376
rect 3360 47320 3428 47376
rect 3484 47320 3552 47376
rect 3608 47320 3676 47376
rect 3732 47320 3800 47376
rect 3856 47320 3924 47376
rect 3980 47320 4048 47376
rect 4104 47320 4172 47376
rect 4228 47320 4296 47376
rect 4352 47320 4420 47376
rect 4476 47320 4544 47376
rect 4600 47320 4668 47376
rect 4724 47320 4734 47376
rect 2798 47252 4734 47320
rect 2798 47196 2808 47252
rect 2864 47196 2932 47252
rect 2988 47196 3056 47252
rect 3112 47196 3180 47252
rect 3236 47196 3304 47252
rect 3360 47196 3428 47252
rect 3484 47196 3552 47252
rect 3608 47196 3676 47252
rect 3732 47196 3800 47252
rect 3856 47196 3924 47252
rect 3980 47196 4048 47252
rect 4104 47196 4172 47252
rect 4228 47196 4296 47252
rect 4352 47196 4420 47252
rect 4476 47196 4544 47252
rect 4600 47196 4668 47252
rect 4724 47196 4734 47252
rect 2798 47128 4734 47196
rect 2798 47072 2808 47128
rect 2864 47072 2932 47128
rect 2988 47072 3056 47128
rect 3112 47072 3180 47128
rect 3236 47072 3304 47128
rect 3360 47072 3428 47128
rect 3484 47072 3552 47128
rect 3608 47072 3676 47128
rect 3732 47072 3800 47128
rect 3856 47072 3924 47128
rect 3980 47072 4048 47128
rect 4104 47072 4172 47128
rect 4228 47072 4296 47128
rect 4352 47072 4420 47128
rect 4476 47072 4544 47128
rect 4600 47072 4668 47128
rect 4724 47072 4734 47128
rect 2798 47004 4734 47072
rect 2798 46948 2808 47004
rect 2864 46948 2932 47004
rect 2988 46948 3056 47004
rect 3112 46948 3180 47004
rect 3236 46948 3304 47004
rect 3360 46948 3428 47004
rect 3484 46948 3552 47004
rect 3608 46948 3676 47004
rect 3732 46948 3800 47004
rect 3856 46948 3924 47004
rect 3980 46948 4048 47004
rect 4104 46948 4172 47004
rect 4228 46948 4296 47004
rect 4352 46948 4420 47004
rect 4476 46948 4544 47004
rect 4600 46948 4668 47004
rect 4724 46948 4734 47004
rect 2798 46880 4734 46948
rect 2798 46824 2808 46880
rect 2864 46824 2932 46880
rect 2988 46824 3056 46880
rect 3112 46824 3180 46880
rect 3236 46824 3304 46880
rect 3360 46824 3428 46880
rect 3484 46824 3552 46880
rect 3608 46824 3676 46880
rect 3732 46824 3800 46880
rect 3856 46824 3924 46880
rect 3980 46824 4048 46880
rect 4104 46824 4172 46880
rect 4228 46824 4296 46880
rect 4352 46824 4420 46880
rect 4476 46824 4544 46880
rect 4600 46824 4668 46880
rect 4724 46824 4734 46880
rect 2798 46756 4734 46824
rect 2798 46700 2808 46756
rect 2864 46700 2932 46756
rect 2988 46700 3056 46756
rect 3112 46700 3180 46756
rect 3236 46700 3304 46756
rect 3360 46700 3428 46756
rect 3484 46700 3552 46756
rect 3608 46700 3676 46756
rect 3732 46700 3800 46756
rect 3856 46700 3924 46756
rect 3980 46700 4048 46756
rect 4104 46700 4172 46756
rect 4228 46700 4296 46756
rect 4352 46700 4420 46756
rect 4476 46700 4544 46756
rect 4600 46700 4668 46756
rect 4724 46700 4734 46756
rect 2798 46632 4734 46700
rect 2798 46576 2808 46632
rect 2864 46576 2932 46632
rect 2988 46576 3056 46632
rect 3112 46576 3180 46632
rect 3236 46576 3304 46632
rect 3360 46576 3428 46632
rect 3484 46576 3552 46632
rect 3608 46576 3676 46632
rect 3732 46576 3800 46632
rect 3856 46576 3924 46632
rect 3980 46576 4048 46632
rect 4104 46576 4172 46632
rect 4228 46576 4296 46632
rect 4352 46576 4420 46632
rect 4476 46576 4544 46632
rect 4600 46576 4668 46632
rect 4724 46576 4734 46632
rect 2798 46508 4734 46576
rect 2798 46452 2808 46508
rect 2864 46452 2932 46508
rect 2988 46452 3056 46508
rect 3112 46452 3180 46508
rect 3236 46452 3304 46508
rect 3360 46452 3428 46508
rect 3484 46452 3552 46508
rect 3608 46452 3676 46508
rect 3732 46452 3800 46508
rect 3856 46452 3924 46508
rect 3980 46452 4048 46508
rect 4104 46452 4172 46508
rect 4228 46452 4296 46508
rect 4352 46452 4420 46508
rect 4476 46452 4544 46508
rect 4600 46452 4668 46508
rect 4724 46452 4734 46508
rect 2798 46442 4734 46452
rect 5168 47748 7104 47758
rect 5168 47692 5178 47748
rect 5234 47692 5302 47748
rect 5358 47692 5426 47748
rect 5482 47692 5550 47748
rect 5606 47692 5674 47748
rect 5730 47692 5798 47748
rect 5854 47692 5922 47748
rect 5978 47692 6046 47748
rect 6102 47692 6170 47748
rect 6226 47692 6294 47748
rect 6350 47692 6418 47748
rect 6474 47692 6542 47748
rect 6598 47692 6666 47748
rect 6722 47692 6790 47748
rect 6846 47692 6914 47748
rect 6970 47692 7038 47748
rect 7094 47692 7104 47748
rect 5168 47624 7104 47692
rect 5168 47568 5178 47624
rect 5234 47568 5302 47624
rect 5358 47568 5426 47624
rect 5482 47568 5550 47624
rect 5606 47568 5674 47624
rect 5730 47568 5798 47624
rect 5854 47568 5922 47624
rect 5978 47568 6046 47624
rect 6102 47568 6170 47624
rect 6226 47568 6294 47624
rect 6350 47568 6418 47624
rect 6474 47568 6542 47624
rect 6598 47568 6666 47624
rect 6722 47568 6790 47624
rect 6846 47568 6914 47624
rect 6970 47568 7038 47624
rect 7094 47568 7104 47624
rect 5168 47500 7104 47568
rect 5168 47444 5178 47500
rect 5234 47444 5302 47500
rect 5358 47444 5426 47500
rect 5482 47444 5550 47500
rect 5606 47444 5674 47500
rect 5730 47444 5798 47500
rect 5854 47444 5922 47500
rect 5978 47444 6046 47500
rect 6102 47444 6170 47500
rect 6226 47444 6294 47500
rect 6350 47444 6418 47500
rect 6474 47444 6542 47500
rect 6598 47444 6666 47500
rect 6722 47444 6790 47500
rect 6846 47444 6914 47500
rect 6970 47444 7038 47500
rect 7094 47444 7104 47500
rect 5168 47376 7104 47444
rect 5168 47320 5178 47376
rect 5234 47320 5302 47376
rect 5358 47320 5426 47376
rect 5482 47320 5550 47376
rect 5606 47320 5674 47376
rect 5730 47320 5798 47376
rect 5854 47320 5922 47376
rect 5978 47320 6046 47376
rect 6102 47320 6170 47376
rect 6226 47320 6294 47376
rect 6350 47320 6418 47376
rect 6474 47320 6542 47376
rect 6598 47320 6666 47376
rect 6722 47320 6790 47376
rect 6846 47320 6914 47376
rect 6970 47320 7038 47376
rect 7094 47320 7104 47376
rect 5168 47252 7104 47320
rect 5168 47196 5178 47252
rect 5234 47196 5302 47252
rect 5358 47196 5426 47252
rect 5482 47196 5550 47252
rect 5606 47196 5674 47252
rect 5730 47196 5798 47252
rect 5854 47196 5922 47252
rect 5978 47196 6046 47252
rect 6102 47196 6170 47252
rect 6226 47196 6294 47252
rect 6350 47196 6418 47252
rect 6474 47196 6542 47252
rect 6598 47196 6666 47252
rect 6722 47196 6790 47252
rect 6846 47196 6914 47252
rect 6970 47196 7038 47252
rect 7094 47196 7104 47252
rect 5168 47128 7104 47196
rect 5168 47072 5178 47128
rect 5234 47072 5302 47128
rect 5358 47072 5426 47128
rect 5482 47072 5550 47128
rect 5606 47072 5674 47128
rect 5730 47072 5798 47128
rect 5854 47072 5922 47128
rect 5978 47072 6046 47128
rect 6102 47072 6170 47128
rect 6226 47072 6294 47128
rect 6350 47072 6418 47128
rect 6474 47072 6542 47128
rect 6598 47072 6666 47128
rect 6722 47072 6790 47128
rect 6846 47072 6914 47128
rect 6970 47072 7038 47128
rect 7094 47072 7104 47128
rect 5168 47004 7104 47072
rect 5168 46948 5178 47004
rect 5234 46948 5302 47004
rect 5358 46948 5426 47004
rect 5482 46948 5550 47004
rect 5606 46948 5674 47004
rect 5730 46948 5798 47004
rect 5854 46948 5922 47004
rect 5978 46948 6046 47004
rect 6102 46948 6170 47004
rect 6226 46948 6294 47004
rect 6350 46948 6418 47004
rect 6474 46948 6542 47004
rect 6598 46948 6666 47004
rect 6722 46948 6790 47004
rect 6846 46948 6914 47004
rect 6970 46948 7038 47004
rect 7094 46948 7104 47004
rect 5168 46880 7104 46948
rect 5168 46824 5178 46880
rect 5234 46824 5302 46880
rect 5358 46824 5426 46880
rect 5482 46824 5550 46880
rect 5606 46824 5674 46880
rect 5730 46824 5798 46880
rect 5854 46824 5922 46880
rect 5978 46824 6046 46880
rect 6102 46824 6170 46880
rect 6226 46824 6294 46880
rect 6350 46824 6418 46880
rect 6474 46824 6542 46880
rect 6598 46824 6666 46880
rect 6722 46824 6790 46880
rect 6846 46824 6914 46880
rect 6970 46824 7038 46880
rect 7094 46824 7104 46880
rect 5168 46756 7104 46824
rect 5168 46700 5178 46756
rect 5234 46700 5302 46756
rect 5358 46700 5426 46756
rect 5482 46700 5550 46756
rect 5606 46700 5674 46756
rect 5730 46700 5798 46756
rect 5854 46700 5922 46756
rect 5978 46700 6046 46756
rect 6102 46700 6170 46756
rect 6226 46700 6294 46756
rect 6350 46700 6418 46756
rect 6474 46700 6542 46756
rect 6598 46700 6666 46756
rect 6722 46700 6790 46756
rect 6846 46700 6914 46756
rect 6970 46700 7038 46756
rect 7094 46700 7104 46756
rect 5168 46632 7104 46700
rect 5168 46576 5178 46632
rect 5234 46576 5302 46632
rect 5358 46576 5426 46632
rect 5482 46576 5550 46632
rect 5606 46576 5674 46632
rect 5730 46576 5798 46632
rect 5854 46576 5922 46632
rect 5978 46576 6046 46632
rect 6102 46576 6170 46632
rect 6226 46576 6294 46632
rect 6350 46576 6418 46632
rect 6474 46576 6542 46632
rect 6598 46576 6666 46632
rect 6722 46576 6790 46632
rect 6846 46576 6914 46632
rect 6970 46576 7038 46632
rect 7094 46576 7104 46632
rect 5168 46508 7104 46576
rect 5168 46452 5178 46508
rect 5234 46452 5302 46508
rect 5358 46452 5426 46508
rect 5482 46452 5550 46508
rect 5606 46452 5674 46508
rect 5730 46452 5798 46508
rect 5854 46452 5922 46508
rect 5978 46452 6046 46508
rect 6102 46452 6170 46508
rect 6226 46452 6294 46508
rect 6350 46452 6418 46508
rect 6474 46452 6542 46508
rect 6598 46452 6666 46508
rect 6722 46452 6790 46508
rect 6846 46452 6914 46508
rect 6970 46452 7038 46508
rect 7094 46452 7104 46508
rect 5168 46442 7104 46452
rect 7874 47748 9810 47758
rect 7874 47692 7884 47748
rect 7940 47692 8008 47748
rect 8064 47692 8132 47748
rect 8188 47692 8256 47748
rect 8312 47692 8380 47748
rect 8436 47692 8504 47748
rect 8560 47692 8628 47748
rect 8684 47692 8752 47748
rect 8808 47692 8876 47748
rect 8932 47692 9000 47748
rect 9056 47692 9124 47748
rect 9180 47692 9248 47748
rect 9304 47692 9372 47748
rect 9428 47692 9496 47748
rect 9552 47692 9620 47748
rect 9676 47692 9744 47748
rect 9800 47692 9810 47748
rect 7874 47624 9810 47692
rect 7874 47568 7884 47624
rect 7940 47568 8008 47624
rect 8064 47568 8132 47624
rect 8188 47568 8256 47624
rect 8312 47568 8380 47624
rect 8436 47568 8504 47624
rect 8560 47568 8628 47624
rect 8684 47568 8752 47624
rect 8808 47568 8876 47624
rect 8932 47568 9000 47624
rect 9056 47568 9124 47624
rect 9180 47568 9248 47624
rect 9304 47568 9372 47624
rect 9428 47568 9496 47624
rect 9552 47568 9620 47624
rect 9676 47568 9744 47624
rect 9800 47568 9810 47624
rect 7874 47500 9810 47568
rect 7874 47444 7884 47500
rect 7940 47444 8008 47500
rect 8064 47444 8132 47500
rect 8188 47444 8256 47500
rect 8312 47444 8380 47500
rect 8436 47444 8504 47500
rect 8560 47444 8628 47500
rect 8684 47444 8752 47500
rect 8808 47444 8876 47500
rect 8932 47444 9000 47500
rect 9056 47444 9124 47500
rect 9180 47444 9248 47500
rect 9304 47444 9372 47500
rect 9428 47444 9496 47500
rect 9552 47444 9620 47500
rect 9676 47444 9744 47500
rect 9800 47444 9810 47500
rect 7874 47376 9810 47444
rect 7874 47320 7884 47376
rect 7940 47320 8008 47376
rect 8064 47320 8132 47376
rect 8188 47320 8256 47376
rect 8312 47320 8380 47376
rect 8436 47320 8504 47376
rect 8560 47320 8628 47376
rect 8684 47320 8752 47376
rect 8808 47320 8876 47376
rect 8932 47320 9000 47376
rect 9056 47320 9124 47376
rect 9180 47320 9248 47376
rect 9304 47320 9372 47376
rect 9428 47320 9496 47376
rect 9552 47320 9620 47376
rect 9676 47320 9744 47376
rect 9800 47320 9810 47376
rect 7874 47252 9810 47320
rect 7874 47196 7884 47252
rect 7940 47196 8008 47252
rect 8064 47196 8132 47252
rect 8188 47196 8256 47252
rect 8312 47196 8380 47252
rect 8436 47196 8504 47252
rect 8560 47196 8628 47252
rect 8684 47196 8752 47252
rect 8808 47196 8876 47252
rect 8932 47196 9000 47252
rect 9056 47196 9124 47252
rect 9180 47196 9248 47252
rect 9304 47196 9372 47252
rect 9428 47196 9496 47252
rect 9552 47196 9620 47252
rect 9676 47196 9744 47252
rect 9800 47196 9810 47252
rect 7874 47128 9810 47196
rect 7874 47072 7884 47128
rect 7940 47072 8008 47128
rect 8064 47072 8132 47128
rect 8188 47072 8256 47128
rect 8312 47072 8380 47128
rect 8436 47072 8504 47128
rect 8560 47072 8628 47128
rect 8684 47072 8752 47128
rect 8808 47072 8876 47128
rect 8932 47072 9000 47128
rect 9056 47072 9124 47128
rect 9180 47072 9248 47128
rect 9304 47072 9372 47128
rect 9428 47072 9496 47128
rect 9552 47072 9620 47128
rect 9676 47072 9744 47128
rect 9800 47072 9810 47128
rect 7874 47004 9810 47072
rect 7874 46948 7884 47004
rect 7940 46948 8008 47004
rect 8064 46948 8132 47004
rect 8188 46948 8256 47004
rect 8312 46948 8380 47004
rect 8436 46948 8504 47004
rect 8560 46948 8628 47004
rect 8684 46948 8752 47004
rect 8808 46948 8876 47004
rect 8932 46948 9000 47004
rect 9056 46948 9124 47004
rect 9180 46948 9248 47004
rect 9304 46948 9372 47004
rect 9428 46948 9496 47004
rect 9552 46948 9620 47004
rect 9676 46948 9744 47004
rect 9800 46948 9810 47004
rect 7874 46880 9810 46948
rect 7874 46824 7884 46880
rect 7940 46824 8008 46880
rect 8064 46824 8132 46880
rect 8188 46824 8256 46880
rect 8312 46824 8380 46880
rect 8436 46824 8504 46880
rect 8560 46824 8628 46880
rect 8684 46824 8752 46880
rect 8808 46824 8876 46880
rect 8932 46824 9000 46880
rect 9056 46824 9124 46880
rect 9180 46824 9248 46880
rect 9304 46824 9372 46880
rect 9428 46824 9496 46880
rect 9552 46824 9620 46880
rect 9676 46824 9744 46880
rect 9800 46824 9810 46880
rect 7874 46756 9810 46824
rect 7874 46700 7884 46756
rect 7940 46700 8008 46756
rect 8064 46700 8132 46756
rect 8188 46700 8256 46756
rect 8312 46700 8380 46756
rect 8436 46700 8504 46756
rect 8560 46700 8628 46756
rect 8684 46700 8752 46756
rect 8808 46700 8876 46756
rect 8932 46700 9000 46756
rect 9056 46700 9124 46756
rect 9180 46700 9248 46756
rect 9304 46700 9372 46756
rect 9428 46700 9496 46756
rect 9552 46700 9620 46756
rect 9676 46700 9744 46756
rect 9800 46700 9810 46756
rect 7874 46632 9810 46700
rect 7874 46576 7884 46632
rect 7940 46576 8008 46632
rect 8064 46576 8132 46632
rect 8188 46576 8256 46632
rect 8312 46576 8380 46632
rect 8436 46576 8504 46632
rect 8560 46576 8628 46632
rect 8684 46576 8752 46632
rect 8808 46576 8876 46632
rect 8932 46576 9000 46632
rect 9056 46576 9124 46632
rect 9180 46576 9248 46632
rect 9304 46576 9372 46632
rect 9428 46576 9496 46632
rect 9552 46576 9620 46632
rect 9676 46576 9744 46632
rect 9800 46576 9810 46632
rect 7874 46508 9810 46576
rect 7874 46452 7884 46508
rect 7940 46452 8008 46508
rect 8064 46452 8132 46508
rect 8188 46452 8256 46508
rect 8312 46452 8380 46508
rect 8436 46452 8504 46508
rect 8560 46452 8628 46508
rect 8684 46452 8752 46508
rect 8808 46452 8876 46508
rect 8932 46452 9000 46508
rect 9056 46452 9124 46508
rect 9180 46452 9248 46508
rect 9304 46452 9372 46508
rect 9428 46452 9496 46508
rect 9552 46452 9620 46508
rect 9676 46452 9744 46508
rect 9800 46452 9810 46508
rect 7874 46442 9810 46452
rect 10244 47748 12180 47758
rect 10244 47692 10254 47748
rect 10310 47692 10378 47748
rect 10434 47692 10502 47748
rect 10558 47692 10626 47748
rect 10682 47692 10750 47748
rect 10806 47692 10874 47748
rect 10930 47692 10998 47748
rect 11054 47692 11122 47748
rect 11178 47692 11246 47748
rect 11302 47692 11370 47748
rect 11426 47692 11494 47748
rect 11550 47692 11618 47748
rect 11674 47692 11742 47748
rect 11798 47692 11866 47748
rect 11922 47692 11990 47748
rect 12046 47692 12114 47748
rect 12170 47692 12180 47748
rect 10244 47624 12180 47692
rect 10244 47568 10254 47624
rect 10310 47568 10378 47624
rect 10434 47568 10502 47624
rect 10558 47568 10626 47624
rect 10682 47568 10750 47624
rect 10806 47568 10874 47624
rect 10930 47568 10998 47624
rect 11054 47568 11122 47624
rect 11178 47568 11246 47624
rect 11302 47568 11370 47624
rect 11426 47568 11494 47624
rect 11550 47568 11618 47624
rect 11674 47568 11742 47624
rect 11798 47568 11866 47624
rect 11922 47568 11990 47624
rect 12046 47568 12114 47624
rect 12170 47568 12180 47624
rect 10244 47500 12180 47568
rect 10244 47444 10254 47500
rect 10310 47444 10378 47500
rect 10434 47444 10502 47500
rect 10558 47444 10626 47500
rect 10682 47444 10750 47500
rect 10806 47444 10874 47500
rect 10930 47444 10998 47500
rect 11054 47444 11122 47500
rect 11178 47444 11246 47500
rect 11302 47444 11370 47500
rect 11426 47444 11494 47500
rect 11550 47444 11618 47500
rect 11674 47444 11742 47500
rect 11798 47444 11866 47500
rect 11922 47444 11990 47500
rect 12046 47444 12114 47500
rect 12170 47444 12180 47500
rect 10244 47376 12180 47444
rect 10244 47320 10254 47376
rect 10310 47320 10378 47376
rect 10434 47320 10502 47376
rect 10558 47320 10626 47376
rect 10682 47320 10750 47376
rect 10806 47320 10874 47376
rect 10930 47320 10998 47376
rect 11054 47320 11122 47376
rect 11178 47320 11246 47376
rect 11302 47320 11370 47376
rect 11426 47320 11494 47376
rect 11550 47320 11618 47376
rect 11674 47320 11742 47376
rect 11798 47320 11866 47376
rect 11922 47320 11990 47376
rect 12046 47320 12114 47376
rect 12170 47320 12180 47376
rect 10244 47252 12180 47320
rect 10244 47196 10254 47252
rect 10310 47196 10378 47252
rect 10434 47196 10502 47252
rect 10558 47196 10626 47252
rect 10682 47196 10750 47252
rect 10806 47196 10874 47252
rect 10930 47196 10998 47252
rect 11054 47196 11122 47252
rect 11178 47196 11246 47252
rect 11302 47196 11370 47252
rect 11426 47196 11494 47252
rect 11550 47196 11618 47252
rect 11674 47196 11742 47252
rect 11798 47196 11866 47252
rect 11922 47196 11990 47252
rect 12046 47196 12114 47252
rect 12170 47196 12180 47252
rect 10244 47128 12180 47196
rect 10244 47072 10254 47128
rect 10310 47072 10378 47128
rect 10434 47072 10502 47128
rect 10558 47072 10626 47128
rect 10682 47072 10750 47128
rect 10806 47072 10874 47128
rect 10930 47072 10998 47128
rect 11054 47072 11122 47128
rect 11178 47072 11246 47128
rect 11302 47072 11370 47128
rect 11426 47072 11494 47128
rect 11550 47072 11618 47128
rect 11674 47072 11742 47128
rect 11798 47072 11866 47128
rect 11922 47072 11990 47128
rect 12046 47072 12114 47128
rect 12170 47072 12180 47128
rect 10244 47004 12180 47072
rect 10244 46948 10254 47004
rect 10310 46948 10378 47004
rect 10434 46948 10502 47004
rect 10558 46948 10626 47004
rect 10682 46948 10750 47004
rect 10806 46948 10874 47004
rect 10930 46948 10998 47004
rect 11054 46948 11122 47004
rect 11178 46948 11246 47004
rect 11302 46948 11370 47004
rect 11426 46948 11494 47004
rect 11550 46948 11618 47004
rect 11674 46948 11742 47004
rect 11798 46948 11866 47004
rect 11922 46948 11990 47004
rect 12046 46948 12114 47004
rect 12170 46948 12180 47004
rect 10244 46880 12180 46948
rect 10244 46824 10254 46880
rect 10310 46824 10378 46880
rect 10434 46824 10502 46880
rect 10558 46824 10626 46880
rect 10682 46824 10750 46880
rect 10806 46824 10874 46880
rect 10930 46824 10998 46880
rect 11054 46824 11122 46880
rect 11178 46824 11246 46880
rect 11302 46824 11370 46880
rect 11426 46824 11494 46880
rect 11550 46824 11618 46880
rect 11674 46824 11742 46880
rect 11798 46824 11866 46880
rect 11922 46824 11990 46880
rect 12046 46824 12114 46880
rect 12170 46824 12180 46880
rect 10244 46756 12180 46824
rect 10244 46700 10254 46756
rect 10310 46700 10378 46756
rect 10434 46700 10502 46756
rect 10558 46700 10626 46756
rect 10682 46700 10750 46756
rect 10806 46700 10874 46756
rect 10930 46700 10998 46756
rect 11054 46700 11122 46756
rect 11178 46700 11246 46756
rect 11302 46700 11370 46756
rect 11426 46700 11494 46756
rect 11550 46700 11618 46756
rect 11674 46700 11742 46756
rect 11798 46700 11866 46756
rect 11922 46700 11990 46756
rect 12046 46700 12114 46756
rect 12170 46700 12180 46756
rect 10244 46632 12180 46700
rect 10244 46576 10254 46632
rect 10310 46576 10378 46632
rect 10434 46576 10502 46632
rect 10558 46576 10626 46632
rect 10682 46576 10750 46632
rect 10806 46576 10874 46632
rect 10930 46576 10998 46632
rect 11054 46576 11122 46632
rect 11178 46576 11246 46632
rect 11302 46576 11370 46632
rect 11426 46576 11494 46632
rect 11550 46576 11618 46632
rect 11674 46576 11742 46632
rect 11798 46576 11866 46632
rect 11922 46576 11990 46632
rect 12046 46576 12114 46632
rect 12170 46576 12180 46632
rect 10244 46508 12180 46576
rect 10244 46452 10254 46508
rect 10310 46452 10378 46508
rect 10434 46452 10502 46508
rect 10558 46452 10626 46508
rect 10682 46452 10750 46508
rect 10806 46452 10874 46508
rect 10930 46452 10998 46508
rect 11054 46452 11122 46508
rect 11178 46452 11246 46508
rect 11302 46452 11370 46508
rect 11426 46452 11494 46508
rect 11550 46452 11618 46508
rect 11674 46452 11742 46508
rect 11798 46452 11866 46508
rect 11922 46452 11990 46508
rect 12046 46452 12114 46508
rect 12170 46452 12180 46508
rect 10244 46442 12180 46452
rect 12861 47748 14673 47758
rect 12861 47692 12871 47748
rect 12927 47692 12995 47748
rect 13051 47692 13119 47748
rect 13175 47692 13243 47748
rect 13299 47692 13367 47748
rect 13423 47692 13491 47748
rect 13547 47692 13615 47748
rect 13671 47692 13739 47748
rect 13795 47692 13863 47748
rect 13919 47692 13987 47748
rect 14043 47692 14111 47748
rect 14167 47692 14235 47748
rect 14291 47692 14359 47748
rect 14415 47692 14483 47748
rect 14539 47692 14607 47748
rect 14663 47692 14673 47748
rect 12861 47624 14673 47692
rect 12861 47568 12871 47624
rect 12927 47568 12995 47624
rect 13051 47568 13119 47624
rect 13175 47568 13243 47624
rect 13299 47568 13367 47624
rect 13423 47568 13491 47624
rect 13547 47568 13615 47624
rect 13671 47568 13739 47624
rect 13795 47568 13863 47624
rect 13919 47568 13987 47624
rect 14043 47568 14111 47624
rect 14167 47568 14235 47624
rect 14291 47568 14359 47624
rect 14415 47568 14483 47624
rect 14539 47568 14607 47624
rect 14663 47568 14673 47624
rect 12861 47500 14673 47568
rect 12861 47444 12871 47500
rect 12927 47444 12995 47500
rect 13051 47444 13119 47500
rect 13175 47444 13243 47500
rect 13299 47444 13367 47500
rect 13423 47444 13491 47500
rect 13547 47444 13615 47500
rect 13671 47444 13739 47500
rect 13795 47444 13863 47500
rect 13919 47444 13987 47500
rect 14043 47444 14111 47500
rect 14167 47444 14235 47500
rect 14291 47444 14359 47500
rect 14415 47444 14483 47500
rect 14539 47444 14607 47500
rect 14663 47444 14673 47500
rect 12861 47376 14673 47444
rect 12861 47320 12871 47376
rect 12927 47320 12995 47376
rect 13051 47320 13119 47376
rect 13175 47320 13243 47376
rect 13299 47320 13367 47376
rect 13423 47320 13491 47376
rect 13547 47320 13615 47376
rect 13671 47320 13739 47376
rect 13795 47320 13863 47376
rect 13919 47320 13987 47376
rect 14043 47320 14111 47376
rect 14167 47320 14235 47376
rect 14291 47320 14359 47376
rect 14415 47320 14483 47376
rect 14539 47320 14607 47376
rect 14663 47320 14673 47376
rect 12861 47252 14673 47320
rect 12861 47196 12871 47252
rect 12927 47196 12995 47252
rect 13051 47196 13119 47252
rect 13175 47196 13243 47252
rect 13299 47196 13367 47252
rect 13423 47196 13491 47252
rect 13547 47196 13615 47252
rect 13671 47196 13739 47252
rect 13795 47196 13863 47252
rect 13919 47196 13987 47252
rect 14043 47196 14111 47252
rect 14167 47196 14235 47252
rect 14291 47196 14359 47252
rect 14415 47196 14483 47252
rect 14539 47196 14607 47252
rect 14663 47196 14673 47252
rect 12861 47128 14673 47196
rect 12861 47072 12871 47128
rect 12927 47072 12995 47128
rect 13051 47072 13119 47128
rect 13175 47072 13243 47128
rect 13299 47072 13367 47128
rect 13423 47072 13491 47128
rect 13547 47072 13615 47128
rect 13671 47072 13739 47128
rect 13795 47072 13863 47128
rect 13919 47072 13987 47128
rect 14043 47072 14111 47128
rect 14167 47072 14235 47128
rect 14291 47072 14359 47128
rect 14415 47072 14483 47128
rect 14539 47072 14607 47128
rect 14663 47072 14673 47128
rect 12861 47004 14673 47072
rect 12861 46948 12871 47004
rect 12927 46948 12995 47004
rect 13051 46948 13119 47004
rect 13175 46948 13243 47004
rect 13299 46948 13367 47004
rect 13423 46948 13491 47004
rect 13547 46948 13615 47004
rect 13671 46948 13739 47004
rect 13795 46948 13863 47004
rect 13919 46948 13987 47004
rect 14043 46948 14111 47004
rect 14167 46948 14235 47004
rect 14291 46948 14359 47004
rect 14415 46948 14483 47004
rect 14539 46948 14607 47004
rect 14663 46948 14673 47004
rect 12861 46880 14673 46948
rect 12861 46824 12871 46880
rect 12927 46824 12995 46880
rect 13051 46824 13119 46880
rect 13175 46824 13243 46880
rect 13299 46824 13367 46880
rect 13423 46824 13491 46880
rect 13547 46824 13615 46880
rect 13671 46824 13739 46880
rect 13795 46824 13863 46880
rect 13919 46824 13987 46880
rect 14043 46824 14111 46880
rect 14167 46824 14235 46880
rect 14291 46824 14359 46880
rect 14415 46824 14483 46880
rect 14539 46824 14607 46880
rect 14663 46824 14673 46880
rect 12861 46756 14673 46824
rect 12861 46700 12871 46756
rect 12927 46700 12995 46756
rect 13051 46700 13119 46756
rect 13175 46700 13243 46756
rect 13299 46700 13367 46756
rect 13423 46700 13491 46756
rect 13547 46700 13615 46756
rect 13671 46700 13739 46756
rect 13795 46700 13863 46756
rect 13919 46700 13987 46756
rect 14043 46700 14111 46756
rect 14167 46700 14235 46756
rect 14291 46700 14359 46756
rect 14415 46700 14483 46756
rect 14539 46700 14607 46756
rect 14663 46700 14673 46756
rect 12861 46632 14673 46700
rect 12861 46576 12871 46632
rect 12927 46576 12995 46632
rect 13051 46576 13119 46632
rect 13175 46576 13243 46632
rect 13299 46576 13367 46632
rect 13423 46576 13491 46632
rect 13547 46576 13615 46632
rect 13671 46576 13739 46632
rect 13795 46576 13863 46632
rect 13919 46576 13987 46632
rect 14043 46576 14111 46632
rect 14167 46576 14235 46632
rect 14291 46576 14359 46632
rect 14415 46576 14483 46632
rect 14539 46576 14607 46632
rect 14663 46576 14673 46632
rect 12861 46508 14673 46576
rect 12861 46452 12871 46508
rect 12927 46452 12995 46508
rect 13051 46452 13119 46508
rect 13175 46452 13243 46508
rect 13299 46452 13367 46508
rect 13423 46452 13491 46508
rect 13547 46452 13615 46508
rect 13671 46452 13739 46508
rect 13795 46452 13863 46508
rect 13919 46452 13987 46508
rect 14043 46452 14111 46508
rect 14167 46452 14235 46508
rect 14291 46452 14359 46508
rect 14415 46452 14483 46508
rect 14539 46452 14607 46508
rect 14663 46452 14673 46508
rect 12861 46442 14673 46452
rect 2481 46148 2681 46158
rect 2481 46092 2491 46148
rect 2547 46092 2615 46148
rect 2671 46092 2681 46148
rect 2481 46024 2681 46092
rect 2481 45968 2491 46024
rect 2547 45968 2615 46024
rect 2671 45968 2681 46024
rect 2481 45900 2681 45968
rect 2481 45844 2491 45900
rect 2547 45844 2615 45900
rect 2671 45844 2681 45900
rect 2481 45776 2681 45844
rect 2481 45720 2491 45776
rect 2547 45720 2615 45776
rect 2671 45720 2681 45776
rect 2481 45652 2681 45720
rect 2481 45596 2491 45652
rect 2547 45596 2615 45652
rect 2671 45596 2681 45652
rect 2481 45528 2681 45596
rect 2481 45472 2491 45528
rect 2547 45472 2615 45528
rect 2671 45472 2681 45528
rect 2481 45404 2681 45472
rect 2481 45348 2491 45404
rect 2547 45348 2615 45404
rect 2671 45348 2681 45404
rect 2481 45280 2681 45348
rect 2481 45224 2491 45280
rect 2547 45224 2615 45280
rect 2671 45224 2681 45280
rect 2481 45156 2681 45224
rect 2481 45100 2491 45156
rect 2547 45100 2615 45156
rect 2671 45100 2681 45156
rect 2481 45032 2681 45100
rect 2481 44976 2491 45032
rect 2547 44976 2615 45032
rect 2671 44976 2681 45032
rect 2481 44908 2681 44976
rect 2481 44852 2491 44908
rect 2547 44852 2615 44908
rect 2671 44852 2681 44908
rect 2481 44842 2681 44852
rect 4851 46148 5051 46158
rect 4851 46092 4861 46148
rect 4917 46092 4985 46148
rect 5041 46092 5051 46148
rect 4851 46024 5051 46092
rect 4851 45968 4861 46024
rect 4917 45968 4985 46024
rect 5041 45968 5051 46024
rect 4851 45900 5051 45968
rect 4851 45844 4861 45900
rect 4917 45844 4985 45900
rect 5041 45844 5051 45900
rect 4851 45776 5051 45844
rect 4851 45720 4861 45776
rect 4917 45720 4985 45776
rect 5041 45720 5051 45776
rect 4851 45652 5051 45720
rect 4851 45596 4861 45652
rect 4917 45596 4985 45652
rect 5041 45596 5051 45652
rect 4851 45528 5051 45596
rect 4851 45472 4861 45528
rect 4917 45472 4985 45528
rect 5041 45472 5051 45528
rect 4851 45404 5051 45472
rect 4851 45348 4861 45404
rect 4917 45348 4985 45404
rect 5041 45348 5051 45404
rect 4851 45280 5051 45348
rect 4851 45224 4861 45280
rect 4917 45224 4985 45280
rect 5041 45224 5051 45280
rect 4851 45156 5051 45224
rect 4851 45100 4861 45156
rect 4917 45100 4985 45156
rect 5041 45100 5051 45156
rect 4851 45032 5051 45100
rect 4851 44976 4861 45032
rect 4917 44976 4985 45032
rect 5041 44976 5051 45032
rect 4851 44908 5051 44976
rect 4851 44852 4861 44908
rect 4917 44852 4985 44908
rect 5041 44852 5051 44908
rect 4851 44842 5051 44852
rect 7265 46148 7713 46158
rect 7265 46092 7275 46148
rect 7331 46092 7399 46148
rect 7455 46092 7523 46148
rect 7579 46092 7647 46148
rect 7703 46092 7713 46148
rect 7265 46024 7713 46092
rect 7265 45968 7275 46024
rect 7331 45968 7399 46024
rect 7455 45968 7523 46024
rect 7579 45968 7647 46024
rect 7703 45968 7713 46024
rect 7265 45900 7713 45968
rect 7265 45844 7275 45900
rect 7331 45844 7399 45900
rect 7455 45844 7523 45900
rect 7579 45844 7647 45900
rect 7703 45844 7713 45900
rect 7265 45776 7713 45844
rect 7265 45720 7275 45776
rect 7331 45720 7399 45776
rect 7455 45720 7523 45776
rect 7579 45720 7647 45776
rect 7703 45720 7713 45776
rect 7265 45652 7713 45720
rect 7265 45596 7275 45652
rect 7331 45596 7399 45652
rect 7455 45596 7523 45652
rect 7579 45596 7647 45652
rect 7703 45596 7713 45652
rect 7265 45528 7713 45596
rect 7265 45472 7275 45528
rect 7331 45472 7399 45528
rect 7455 45472 7523 45528
rect 7579 45472 7647 45528
rect 7703 45472 7713 45528
rect 7265 45404 7713 45472
rect 7265 45348 7275 45404
rect 7331 45348 7399 45404
rect 7455 45348 7523 45404
rect 7579 45348 7647 45404
rect 7703 45348 7713 45404
rect 7265 45280 7713 45348
rect 7265 45224 7275 45280
rect 7331 45224 7399 45280
rect 7455 45224 7523 45280
rect 7579 45224 7647 45280
rect 7703 45224 7713 45280
rect 7265 45156 7713 45224
rect 7265 45100 7275 45156
rect 7331 45100 7399 45156
rect 7455 45100 7523 45156
rect 7579 45100 7647 45156
rect 7703 45100 7713 45156
rect 7265 45032 7713 45100
rect 7265 44976 7275 45032
rect 7331 44976 7399 45032
rect 7455 44976 7523 45032
rect 7579 44976 7647 45032
rect 7703 44976 7713 45032
rect 7265 44908 7713 44976
rect 7265 44852 7275 44908
rect 7331 44852 7399 44908
rect 7455 44852 7523 44908
rect 7579 44852 7647 44908
rect 7703 44852 7713 44908
rect 7265 44842 7713 44852
rect 9927 46148 10127 46158
rect 9927 46092 9937 46148
rect 9993 46092 10061 46148
rect 10117 46092 10127 46148
rect 9927 46024 10127 46092
rect 9927 45968 9937 46024
rect 9993 45968 10061 46024
rect 10117 45968 10127 46024
rect 9927 45900 10127 45968
rect 9927 45844 9937 45900
rect 9993 45844 10061 45900
rect 10117 45844 10127 45900
rect 9927 45776 10127 45844
rect 9927 45720 9937 45776
rect 9993 45720 10061 45776
rect 10117 45720 10127 45776
rect 9927 45652 10127 45720
rect 9927 45596 9937 45652
rect 9993 45596 10061 45652
rect 10117 45596 10127 45652
rect 9927 45528 10127 45596
rect 9927 45472 9937 45528
rect 9993 45472 10061 45528
rect 10117 45472 10127 45528
rect 9927 45404 10127 45472
rect 9927 45348 9937 45404
rect 9993 45348 10061 45404
rect 10117 45348 10127 45404
rect 9927 45280 10127 45348
rect 9927 45224 9937 45280
rect 9993 45224 10061 45280
rect 10117 45224 10127 45280
rect 9927 45156 10127 45224
rect 9927 45100 9937 45156
rect 9993 45100 10061 45156
rect 10117 45100 10127 45156
rect 9927 45032 10127 45100
rect 9927 44976 9937 45032
rect 9993 44976 10061 45032
rect 10117 44976 10127 45032
rect 9927 44908 10127 44976
rect 9927 44852 9937 44908
rect 9993 44852 10061 44908
rect 10117 44852 10127 44908
rect 9927 44842 10127 44852
rect 12297 46148 12497 46158
rect 12297 46092 12307 46148
rect 12363 46092 12431 46148
rect 12487 46092 12497 46148
rect 12297 46024 12497 46092
rect 12297 45968 12307 46024
rect 12363 45968 12431 46024
rect 12487 45968 12497 46024
rect 12297 45900 12497 45968
rect 12297 45844 12307 45900
rect 12363 45844 12431 45900
rect 12487 45844 12497 45900
rect 12297 45776 12497 45844
rect 12297 45720 12307 45776
rect 12363 45720 12431 45776
rect 12487 45720 12497 45776
rect 12297 45652 12497 45720
rect 12297 45596 12307 45652
rect 12363 45596 12431 45652
rect 12487 45596 12497 45652
rect 12297 45528 12497 45596
rect 12297 45472 12307 45528
rect 12363 45472 12431 45528
rect 12487 45472 12497 45528
rect 12297 45404 12497 45472
rect 12297 45348 12307 45404
rect 12363 45348 12431 45404
rect 12487 45348 12497 45404
rect 12297 45280 12497 45348
rect 12297 45224 12307 45280
rect 12363 45224 12431 45280
rect 12487 45224 12497 45280
rect 12297 45156 12497 45224
rect 12297 45100 12307 45156
rect 12363 45100 12431 45156
rect 12487 45100 12497 45156
rect 12297 45032 12497 45100
rect 12297 44976 12307 45032
rect 12363 44976 12431 45032
rect 12487 44976 12497 45032
rect 12297 44908 12497 44976
rect 12297 44852 12307 44908
rect 12363 44852 12431 44908
rect 12487 44852 12497 44908
rect 12297 44842 12497 44852
rect 305 44548 2117 44558
rect 305 44492 315 44548
rect 371 44492 439 44548
rect 495 44492 563 44548
rect 619 44492 687 44548
rect 743 44492 811 44548
rect 867 44492 935 44548
rect 991 44492 1059 44548
rect 1115 44492 1183 44548
rect 1239 44492 1307 44548
rect 1363 44492 1431 44548
rect 1487 44492 1555 44548
rect 1611 44492 1679 44548
rect 1735 44492 1803 44548
rect 1859 44492 1927 44548
rect 1983 44492 2051 44548
rect 2107 44492 2117 44548
rect 305 44424 2117 44492
rect 305 44368 315 44424
rect 371 44368 439 44424
rect 495 44368 563 44424
rect 619 44368 687 44424
rect 743 44368 811 44424
rect 867 44368 935 44424
rect 991 44368 1059 44424
rect 1115 44368 1183 44424
rect 1239 44368 1307 44424
rect 1363 44368 1431 44424
rect 1487 44368 1555 44424
rect 1611 44368 1679 44424
rect 1735 44368 1803 44424
rect 1859 44368 1927 44424
rect 1983 44368 2051 44424
rect 2107 44368 2117 44424
rect 305 44300 2117 44368
rect 305 44244 315 44300
rect 371 44244 439 44300
rect 495 44244 563 44300
rect 619 44244 687 44300
rect 743 44244 811 44300
rect 867 44244 935 44300
rect 991 44244 1059 44300
rect 1115 44244 1183 44300
rect 1239 44244 1307 44300
rect 1363 44244 1431 44300
rect 1487 44244 1555 44300
rect 1611 44244 1679 44300
rect 1735 44244 1803 44300
rect 1859 44244 1927 44300
rect 1983 44244 2051 44300
rect 2107 44244 2117 44300
rect 305 44176 2117 44244
rect 305 44120 315 44176
rect 371 44120 439 44176
rect 495 44120 563 44176
rect 619 44120 687 44176
rect 743 44120 811 44176
rect 867 44120 935 44176
rect 991 44120 1059 44176
rect 1115 44120 1183 44176
rect 1239 44120 1307 44176
rect 1363 44120 1431 44176
rect 1487 44120 1555 44176
rect 1611 44120 1679 44176
rect 1735 44120 1803 44176
rect 1859 44120 1927 44176
rect 1983 44120 2051 44176
rect 2107 44120 2117 44176
rect 305 44052 2117 44120
rect 305 43996 315 44052
rect 371 43996 439 44052
rect 495 43996 563 44052
rect 619 43996 687 44052
rect 743 43996 811 44052
rect 867 43996 935 44052
rect 991 43996 1059 44052
rect 1115 43996 1183 44052
rect 1239 43996 1307 44052
rect 1363 43996 1431 44052
rect 1487 43996 1555 44052
rect 1611 43996 1679 44052
rect 1735 43996 1803 44052
rect 1859 43996 1927 44052
rect 1983 43996 2051 44052
rect 2107 43996 2117 44052
rect 305 43928 2117 43996
rect 305 43872 315 43928
rect 371 43872 439 43928
rect 495 43872 563 43928
rect 619 43872 687 43928
rect 743 43872 811 43928
rect 867 43872 935 43928
rect 991 43872 1059 43928
rect 1115 43872 1183 43928
rect 1239 43872 1307 43928
rect 1363 43872 1431 43928
rect 1487 43872 1555 43928
rect 1611 43872 1679 43928
rect 1735 43872 1803 43928
rect 1859 43872 1927 43928
rect 1983 43872 2051 43928
rect 2107 43872 2117 43928
rect 305 43804 2117 43872
rect 305 43748 315 43804
rect 371 43748 439 43804
rect 495 43748 563 43804
rect 619 43748 687 43804
rect 743 43748 811 43804
rect 867 43748 935 43804
rect 991 43748 1059 43804
rect 1115 43748 1183 43804
rect 1239 43748 1307 43804
rect 1363 43748 1431 43804
rect 1487 43748 1555 43804
rect 1611 43748 1679 43804
rect 1735 43748 1803 43804
rect 1859 43748 1927 43804
rect 1983 43748 2051 43804
rect 2107 43748 2117 43804
rect 305 43680 2117 43748
rect 305 43624 315 43680
rect 371 43624 439 43680
rect 495 43624 563 43680
rect 619 43624 687 43680
rect 743 43624 811 43680
rect 867 43624 935 43680
rect 991 43624 1059 43680
rect 1115 43624 1183 43680
rect 1239 43624 1307 43680
rect 1363 43624 1431 43680
rect 1487 43624 1555 43680
rect 1611 43624 1679 43680
rect 1735 43624 1803 43680
rect 1859 43624 1927 43680
rect 1983 43624 2051 43680
rect 2107 43624 2117 43680
rect 305 43556 2117 43624
rect 305 43500 315 43556
rect 371 43500 439 43556
rect 495 43500 563 43556
rect 619 43500 687 43556
rect 743 43500 811 43556
rect 867 43500 935 43556
rect 991 43500 1059 43556
rect 1115 43500 1183 43556
rect 1239 43500 1307 43556
rect 1363 43500 1431 43556
rect 1487 43500 1555 43556
rect 1611 43500 1679 43556
rect 1735 43500 1803 43556
rect 1859 43500 1927 43556
rect 1983 43500 2051 43556
rect 2107 43500 2117 43556
rect 305 43432 2117 43500
rect 305 43376 315 43432
rect 371 43376 439 43432
rect 495 43376 563 43432
rect 619 43376 687 43432
rect 743 43376 811 43432
rect 867 43376 935 43432
rect 991 43376 1059 43432
rect 1115 43376 1183 43432
rect 1239 43376 1307 43432
rect 1363 43376 1431 43432
rect 1487 43376 1555 43432
rect 1611 43376 1679 43432
rect 1735 43376 1803 43432
rect 1859 43376 1927 43432
rect 1983 43376 2051 43432
rect 2107 43376 2117 43432
rect 305 43308 2117 43376
rect 305 43252 315 43308
rect 371 43252 439 43308
rect 495 43252 563 43308
rect 619 43252 687 43308
rect 743 43252 811 43308
rect 867 43252 935 43308
rect 991 43252 1059 43308
rect 1115 43252 1183 43308
rect 1239 43252 1307 43308
rect 1363 43252 1431 43308
rect 1487 43252 1555 43308
rect 1611 43252 1679 43308
rect 1735 43252 1803 43308
rect 1859 43252 1927 43308
rect 1983 43252 2051 43308
rect 2107 43252 2117 43308
rect 305 43242 2117 43252
rect 2798 44548 4734 44558
rect 2798 44492 2808 44548
rect 2864 44492 2932 44548
rect 2988 44492 3056 44548
rect 3112 44492 3180 44548
rect 3236 44492 3304 44548
rect 3360 44492 3428 44548
rect 3484 44492 3552 44548
rect 3608 44492 3676 44548
rect 3732 44492 3800 44548
rect 3856 44492 3924 44548
rect 3980 44492 4048 44548
rect 4104 44492 4172 44548
rect 4228 44492 4296 44548
rect 4352 44492 4420 44548
rect 4476 44492 4544 44548
rect 4600 44492 4668 44548
rect 4724 44492 4734 44548
rect 2798 44424 4734 44492
rect 2798 44368 2808 44424
rect 2864 44368 2932 44424
rect 2988 44368 3056 44424
rect 3112 44368 3180 44424
rect 3236 44368 3304 44424
rect 3360 44368 3428 44424
rect 3484 44368 3552 44424
rect 3608 44368 3676 44424
rect 3732 44368 3800 44424
rect 3856 44368 3924 44424
rect 3980 44368 4048 44424
rect 4104 44368 4172 44424
rect 4228 44368 4296 44424
rect 4352 44368 4420 44424
rect 4476 44368 4544 44424
rect 4600 44368 4668 44424
rect 4724 44368 4734 44424
rect 2798 44300 4734 44368
rect 2798 44244 2808 44300
rect 2864 44244 2932 44300
rect 2988 44244 3056 44300
rect 3112 44244 3180 44300
rect 3236 44244 3304 44300
rect 3360 44244 3428 44300
rect 3484 44244 3552 44300
rect 3608 44244 3676 44300
rect 3732 44244 3800 44300
rect 3856 44244 3924 44300
rect 3980 44244 4048 44300
rect 4104 44244 4172 44300
rect 4228 44244 4296 44300
rect 4352 44244 4420 44300
rect 4476 44244 4544 44300
rect 4600 44244 4668 44300
rect 4724 44244 4734 44300
rect 2798 44176 4734 44244
rect 2798 44120 2808 44176
rect 2864 44120 2932 44176
rect 2988 44120 3056 44176
rect 3112 44120 3180 44176
rect 3236 44120 3304 44176
rect 3360 44120 3428 44176
rect 3484 44120 3552 44176
rect 3608 44120 3676 44176
rect 3732 44120 3800 44176
rect 3856 44120 3924 44176
rect 3980 44120 4048 44176
rect 4104 44120 4172 44176
rect 4228 44120 4296 44176
rect 4352 44120 4420 44176
rect 4476 44120 4544 44176
rect 4600 44120 4668 44176
rect 4724 44120 4734 44176
rect 2798 44052 4734 44120
rect 2798 43996 2808 44052
rect 2864 43996 2932 44052
rect 2988 43996 3056 44052
rect 3112 43996 3180 44052
rect 3236 43996 3304 44052
rect 3360 43996 3428 44052
rect 3484 43996 3552 44052
rect 3608 43996 3676 44052
rect 3732 43996 3800 44052
rect 3856 43996 3924 44052
rect 3980 43996 4048 44052
rect 4104 43996 4172 44052
rect 4228 43996 4296 44052
rect 4352 43996 4420 44052
rect 4476 43996 4544 44052
rect 4600 43996 4668 44052
rect 4724 43996 4734 44052
rect 2798 43928 4734 43996
rect 2798 43872 2808 43928
rect 2864 43872 2932 43928
rect 2988 43872 3056 43928
rect 3112 43872 3180 43928
rect 3236 43872 3304 43928
rect 3360 43872 3428 43928
rect 3484 43872 3552 43928
rect 3608 43872 3676 43928
rect 3732 43872 3800 43928
rect 3856 43872 3924 43928
rect 3980 43872 4048 43928
rect 4104 43872 4172 43928
rect 4228 43872 4296 43928
rect 4352 43872 4420 43928
rect 4476 43872 4544 43928
rect 4600 43872 4668 43928
rect 4724 43872 4734 43928
rect 2798 43804 4734 43872
rect 2798 43748 2808 43804
rect 2864 43748 2932 43804
rect 2988 43748 3056 43804
rect 3112 43748 3180 43804
rect 3236 43748 3304 43804
rect 3360 43748 3428 43804
rect 3484 43748 3552 43804
rect 3608 43748 3676 43804
rect 3732 43748 3800 43804
rect 3856 43748 3924 43804
rect 3980 43748 4048 43804
rect 4104 43748 4172 43804
rect 4228 43748 4296 43804
rect 4352 43748 4420 43804
rect 4476 43748 4544 43804
rect 4600 43748 4668 43804
rect 4724 43748 4734 43804
rect 2798 43680 4734 43748
rect 2798 43624 2808 43680
rect 2864 43624 2932 43680
rect 2988 43624 3056 43680
rect 3112 43624 3180 43680
rect 3236 43624 3304 43680
rect 3360 43624 3428 43680
rect 3484 43624 3552 43680
rect 3608 43624 3676 43680
rect 3732 43624 3800 43680
rect 3856 43624 3924 43680
rect 3980 43624 4048 43680
rect 4104 43624 4172 43680
rect 4228 43624 4296 43680
rect 4352 43624 4420 43680
rect 4476 43624 4544 43680
rect 4600 43624 4668 43680
rect 4724 43624 4734 43680
rect 2798 43556 4734 43624
rect 2798 43500 2808 43556
rect 2864 43500 2932 43556
rect 2988 43500 3056 43556
rect 3112 43500 3180 43556
rect 3236 43500 3304 43556
rect 3360 43500 3428 43556
rect 3484 43500 3552 43556
rect 3608 43500 3676 43556
rect 3732 43500 3800 43556
rect 3856 43500 3924 43556
rect 3980 43500 4048 43556
rect 4104 43500 4172 43556
rect 4228 43500 4296 43556
rect 4352 43500 4420 43556
rect 4476 43500 4544 43556
rect 4600 43500 4668 43556
rect 4724 43500 4734 43556
rect 2798 43432 4734 43500
rect 2798 43376 2808 43432
rect 2864 43376 2932 43432
rect 2988 43376 3056 43432
rect 3112 43376 3180 43432
rect 3236 43376 3304 43432
rect 3360 43376 3428 43432
rect 3484 43376 3552 43432
rect 3608 43376 3676 43432
rect 3732 43376 3800 43432
rect 3856 43376 3924 43432
rect 3980 43376 4048 43432
rect 4104 43376 4172 43432
rect 4228 43376 4296 43432
rect 4352 43376 4420 43432
rect 4476 43376 4544 43432
rect 4600 43376 4668 43432
rect 4724 43376 4734 43432
rect 2798 43308 4734 43376
rect 2798 43252 2808 43308
rect 2864 43252 2932 43308
rect 2988 43252 3056 43308
rect 3112 43252 3180 43308
rect 3236 43252 3304 43308
rect 3360 43252 3428 43308
rect 3484 43252 3552 43308
rect 3608 43252 3676 43308
rect 3732 43252 3800 43308
rect 3856 43252 3924 43308
rect 3980 43252 4048 43308
rect 4104 43252 4172 43308
rect 4228 43252 4296 43308
rect 4352 43252 4420 43308
rect 4476 43252 4544 43308
rect 4600 43252 4668 43308
rect 4724 43252 4734 43308
rect 2798 43242 4734 43252
rect 5168 44548 7104 44558
rect 5168 44492 5178 44548
rect 5234 44492 5302 44548
rect 5358 44492 5426 44548
rect 5482 44492 5550 44548
rect 5606 44492 5674 44548
rect 5730 44492 5798 44548
rect 5854 44492 5922 44548
rect 5978 44492 6046 44548
rect 6102 44492 6170 44548
rect 6226 44492 6294 44548
rect 6350 44492 6418 44548
rect 6474 44492 6542 44548
rect 6598 44492 6666 44548
rect 6722 44492 6790 44548
rect 6846 44492 6914 44548
rect 6970 44492 7038 44548
rect 7094 44492 7104 44548
rect 5168 44424 7104 44492
rect 5168 44368 5178 44424
rect 5234 44368 5302 44424
rect 5358 44368 5426 44424
rect 5482 44368 5550 44424
rect 5606 44368 5674 44424
rect 5730 44368 5798 44424
rect 5854 44368 5922 44424
rect 5978 44368 6046 44424
rect 6102 44368 6170 44424
rect 6226 44368 6294 44424
rect 6350 44368 6418 44424
rect 6474 44368 6542 44424
rect 6598 44368 6666 44424
rect 6722 44368 6790 44424
rect 6846 44368 6914 44424
rect 6970 44368 7038 44424
rect 7094 44368 7104 44424
rect 5168 44300 7104 44368
rect 5168 44244 5178 44300
rect 5234 44244 5302 44300
rect 5358 44244 5426 44300
rect 5482 44244 5550 44300
rect 5606 44244 5674 44300
rect 5730 44244 5798 44300
rect 5854 44244 5922 44300
rect 5978 44244 6046 44300
rect 6102 44244 6170 44300
rect 6226 44244 6294 44300
rect 6350 44244 6418 44300
rect 6474 44244 6542 44300
rect 6598 44244 6666 44300
rect 6722 44244 6790 44300
rect 6846 44244 6914 44300
rect 6970 44244 7038 44300
rect 7094 44244 7104 44300
rect 5168 44176 7104 44244
rect 5168 44120 5178 44176
rect 5234 44120 5302 44176
rect 5358 44120 5426 44176
rect 5482 44120 5550 44176
rect 5606 44120 5674 44176
rect 5730 44120 5798 44176
rect 5854 44120 5922 44176
rect 5978 44120 6046 44176
rect 6102 44120 6170 44176
rect 6226 44120 6294 44176
rect 6350 44120 6418 44176
rect 6474 44120 6542 44176
rect 6598 44120 6666 44176
rect 6722 44120 6790 44176
rect 6846 44120 6914 44176
rect 6970 44120 7038 44176
rect 7094 44120 7104 44176
rect 5168 44052 7104 44120
rect 5168 43996 5178 44052
rect 5234 43996 5302 44052
rect 5358 43996 5426 44052
rect 5482 43996 5550 44052
rect 5606 43996 5674 44052
rect 5730 43996 5798 44052
rect 5854 43996 5922 44052
rect 5978 43996 6046 44052
rect 6102 43996 6170 44052
rect 6226 43996 6294 44052
rect 6350 43996 6418 44052
rect 6474 43996 6542 44052
rect 6598 43996 6666 44052
rect 6722 43996 6790 44052
rect 6846 43996 6914 44052
rect 6970 43996 7038 44052
rect 7094 43996 7104 44052
rect 5168 43928 7104 43996
rect 5168 43872 5178 43928
rect 5234 43872 5302 43928
rect 5358 43872 5426 43928
rect 5482 43872 5550 43928
rect 5606 43872 5674 43928
rect 5730 43872 5798 43928
rect 5854 43872 5922 43928
rect 5978 43872 6046 43928
rect 6102 43872 6170 43928
rect 6226 43872 6294 43928
rect 6350 43872 6418 43928
rect 6474 43872 6542 43928
rect 6598 43872 6666 43928
rect 6722 43872 6790 43928
rect 6846 43872 6914 43928
rect 6970 43872 7038 43928
rect 7094 43872 7104 43928
rect 5168 43804 7104 43872
rect 5168 43748 5178 43804
rect 5234 43748 5302 43804
rect 5358 43748 5426 43804
rect 5482 43748 5550 43804
rect 5606 43748 5674 43804
rect 5730 43748 5798 43804
rect 5854 43748 5922 43804
rect 5978 43748 6046 43804
rect 6102 43748 6170 43804
rect 6226 43748 6294 43804
rect 6350 43748 6418 43804
rect 6474 43748 6542 43804
rect 6598 43748 6666 43804
rect 6722 43748 6790 43804
rect 6846 43748 6914 43804
rect 6970 43748 7038 43804
rect 7094 43748 7104 43804
rect 5168 43680 7104 43748
rect 5168 43624 5178 43680
rect 5234 43624 5302 43680
rect 5358 43624 5426 43680
rect 5482 43624 5550 43680
rect 5606 43624 5674 43680
rect 5730 43624 5798 43680
rect 5854 43624 5922 43680
rect 5978 43624 6046 43680
rect 6102 43624 6170 43680
rect 6226 43624 6294 43680
rect 6350 43624 6418 43680
rect 6474 43624 6542 43680
rect 6598 43624 6666 43680
rect 6722 43624 6790 43680
rect 6846 43624 6914 43680
rect 6970 43624 7038 43680
rect 7094 43624 7104 43680
rect 5168 43556 7104 43624
rect 5168 43500 5178 43556
rect 5234 43500 5302 43556
rect 5358 43500 5426 43556
rect 5482 43500 5550 43556
rect 5606 43500 5674 43556
rect 5730 43500 5798 43556
rect 5854 43500 5922 43556
rect 5978 43500 6046 43556
rect 6102 43500 6170 43556
rect 6226 43500 6294 43556
rect 6350 43500 6418 43556
rect 6474 43500 6542 43556
rect 6598 43500 6666 43556
rect 6722 43500 6790 43556
rect 6846 43500 6914 43556
rect 6970 43500 7038 43556
rect 7094 43500 7104 43556
rect 5168 43432 7104 43500
rect 5168 43376 5178 43432
rect 5234 43376 5302 43432
rect 5358 43376 5426 43432
rect 5482 43376 5550 43432
rect 5606 43376 5674 43432
rect 5730 43376 5798 43432
rect 5854 43376 5922 43432
rect 5978 43376 6046 43432
rect 6102 43376 6170 43432
rect 6226 43376 6294 43432
rect 6350 43376 6418 43432
rect 6474 43376 6542 43432
rect 6598 43376 6666 43432
rect 6722 43376 6790 43432
rect 6846 43376 6914 43432
rect 6970 43376 7038 43432
rect 7094 43376 7104 43432
rect 5168 43308 7104 43376
rect 5168 43252 5178 43308
rect 5234 43252 5302 43308
rect 5358 43252 5426 43308
rect 5482 43252 5550 43308
rect 5606 43252 5674 43308
rect 5730 43252 5798 43308
rect 5854 43252 5922 43308
rect 5978 43252 6046 43308
rect 6102 43252 6170 43308
rect 6226 43252 6294 43308
rect 6350 43252 6418 43308
rect 6474 43252 6542 43308
rect 6598 43252 6666 43308
rect 6722 43252 6790 43308
rect 6846 43252 6914 43308
rect 6970 43252 7038 43308
rect 7094 43252 7104 43308
rect 5168 43242 7104 43252
rect 7874 44548 9810 44558
rect 7874 44492 7884 44548
rect 7940 44492 8008 44548
rect 8064 44492 8132 44548
rect 8188 44492 8256 44548
rect 8312 44492 8380 44548
rect 8436 44492 8504 44548
rect 8560 44492 8628 44548
rect 8684 44492 8752 44548
rect 8808 44492 8876 44548
rect 8932 44492 9000 44548
rect 9056 44492 9124 44548
rect 9180 44492 9248 44548
rect 9304 44492 9372 44548
rect 9428 44492 9496 44548
rect 9552 44492 9620 44548
rect 9676 44492 9744 44548
rect 9800 44492 9810 44548
rect 7874 44424 9810 44492
rect 7874 44368 7884 44424
rect 7940 44368 8008 44424
rect 8064 44368 8132 44424
rect 8188 44368 8256 44424
rect 8312 44368 8380 44424
rect 8436 44368 8504 44424
rect 8560 44368 8628 44424
rect 8684 44368 8752 44424
rect 8808 44368 8876 44424
rect 8932 44368 9000 44424
rect 9056 44368 9124 44424
rect 9180 44368 9248 44424
rect 9304 44368 9372 44424
rect 9428 44368 9496 44424
rect 9552 44368 9620 44424
rect 9676 44368 9744 44424
rect 9800 44368 9810 44424
rect 7874 44300 9810 44368
rect 7874 44244 7884 44300
rect 7940 44244 8008 44300
rect 8064 44244 8132 44300
rect 8188 44244 8256 44300
rect 8312 44244 8380 44300
rect 8436 44244 8504 44300
rect 8560 44244 8628 44300
rect 8684 44244 8752 44300
rect 8808 44244 8876 44300
rect 8932 44244 9000 44300
rect 9056 44244 9124 44300
rect 9180 44244 9248 44300
rect 9304 44244 9372 44300
rect 9428 44244 9496 44300
rect 9552 44244 9620 44300
rect 9676 44244 9744 44300
rect 9800 44244 9810 44300
rect 7874 44176 9810 44244
rect 7874 44120 7884 44176
rect 7940 44120 8008 44176
rect 8064 44120 8132 44176
rect 8188 44120 8256 44176
rect 8312 44120 8380 44176
rect 8436 44120 8504 44176
rect 8560 44120 8628 44176
rect 8684 44120 8752 44176
rect 8808 44120 8876 44176
rect 8932 44120 9000 44176
rect 9056 44120 9124 44176
rect 9180 44120 9248 44176
rect 9304 44120 9372 44176
rect 9428 44120 9496 44176
rect 9552 44120 9620 44176
rect 9676 44120 9744 44176
rect 9800 44120 9810 44176
rect 7874 44052 9810 44120
rect 7874 43996 7884 44052
rect 7940 43996 8008 44052
rect 8064 43996 8132 44052
rect 8188 43996 8256 44052
rect 8312 43996 8380 44052
rect 8436 43996 8504 44052
rect 8560 43996 8628 44052
rect 8684 43996 8752 44052
rect 8808 43996 8876 44052
rect 8932 43996 9000 44052
rect 9056 43996 9124 44052
rect 9180 43996 9248 44052
rect 9304 43996 9372 44052
rect 9428 43996 9496 44052
rect 9552 43996 9620 44052
rect 9676 43996 9744 44052
rect 9800 43996 9810 44052
rect 7874 43928 9810 43996
rect 7874 43872 7884 43928
rect 7940 43872 8008 43928
rect 8064 43872 8132 43928
rect 8188 43872 8256 43928
rect 8312 43872 8380 43928
rect 8436 43872 8504 43928
rect 8560 43872 8628 43928
rect 8684 43872 8752 43928
rect 8808 43872 8876 43928
rect 8932 43872 9000 43928
rect 9056 43872 9124 43928
rect 9180 43872 9248 43928
rect 9304 43872 9372 43928
rect 9428 43872 9496 43928
rect 9552 43872 9620 43928
rect 9676 43872 9744 43928
rect 9800 43872 9810 43928
rect 7874 43804 9810 43872
rect 7874 43748 7884 43804
rect 7940 43748 8008 43804
rect 8064 43748 8132 43804
rect 8188 43748 8256 43804
rect 8312 43748 8380 43804
rect 8436 43748 8504 43804
rect 8560 43748 8628 43804
rect 8684 43748 8752 43804
rect 8808 43748 8876 43804
rect 8932 43748 9000 43804
rect 9056 43748 9124 43804
rect 9180 43748 9248 43804
rect 9304 43748 9372 43804
rect 9428 43748 9496 43804
rect 9552 43748 9620 43804
rect 9676 43748 9744 43804
rect 9800 43748 9810 43804
rect 7874 43680 9810 43748
rect 7874 43624 7884 43680
rect 7940 43624 8008 43680
rect 8064 43624 8132 43680
rect 8188 43624 8256 43680
rect 8312 43624 8380 43680
rect 8436 43624 8504 43680
rect 8560 43624 8628 43680
rect 8684 43624 8752 43680
rect 8808 43624 8876 43680
rect 8932 43624 9000 43680
rect 9056 43624 9124 43680
rect 9180 43624 9248 43680
rect 9304 43624 9372 43680
rect 9428 43624 9496 43680
rect 9552 43624 9620 43680
rect 9676 43624 9744 43680
rect 9800 43624 9810 43680
rect 7874 43556 9810 43624
rect 7874 43500 7884 43556
rect 7940 43500 8008 43556
rect 8064 43500 8132 43556
rect 8188 43500 8256 43556
rect 8312 43500 8380 43556
rect 8436 43500 8504 43556
rect 8560 43500 8628 43556
rect 8684 43500 8752 43556
rect 8808 43500 8876 43556
rect 8932 43500 9000 43556
rect 9056 43500 9124 43556
rect 9180 43500 9248 43556
rect 9304 43500 9372 43556
rect 9428 43500 9496 43556
rect 9552 43500 9620 43556
rect 9676 43500 9744 43556
rect 9800 43500 9810 43556
rect 7874 43432 9810 43500
rect 7874 43376 7884 43432
rect 7940 43376 8008 43432
rect 8064 43376 8132 43432
rect 8188 43376 8256 43432
rect 8312 43376 8380 43432
rect 8436 43376 8504 43432
rect 8560 43376 8628 43432
rect 8684 43376 8752 43432
rect 8808 43376 8876 43432
rect 8932 43376 9000 43432
rect 9056 43376 9124 43432
rect 9180 43376 9248 43432
rect 9304 43376 9372 43432
rect 9428 43376 9496 43432
rect 9552 43376 9620 43432
rect 9676 43376 9744 43432
rect 9800 43376 9810 43432
rect 7874 43308 9810 43376
rect 7874 43252 7884 43308
rect 7940 43252 8008 43308
rect 8064 43252 8132 43308
rect 8188 43252 8256 43308
rect 8312 43252 8380 43308
rect 8436 43252 8504 43308
rect 8560 43252 8628 43308
rect 8684 43252 8752 43308
rect 8808 43252 8876 43308
rect 8932 43252 9000 43308
rect 9056 43252 9124 43308
rect 9180 43252 9248 43308
rect 9304 43252 9372 43308
rect 9428 43252 9496 43308
rect 9552 43252 9620 43308
rect 9676 43252 9744 43308
rect 9800 43252 9810 43308
rect 7874 43242 9810 43252
rect 10244 44548 12180 44558
rect 10244 44492 10254 44548
rect 10310 44492 10378 44548
rect 10434 44492 10502 44548
rect 10558 44492 10626 44548
rect 10682 44492 10750 44548
rect 10806 44492 10874 44548
rect 10930 44492 10998 44548
rect 11054 44492 11122 44548
rect 11178 44492 11246 44548
rect 11302 44492 11370 44548
rect 11426 44492 11494 44548
rect 11550 44492 11618 44548
rect 11674 44492 11742 44548
rect 11798 44492 11866 44548
rect 11922 44492 11990 44548
rect 12046 44492 12114 44548
rect 12170 44492 12180 44548
rect 10244 44424 12180 44492
rect 10244 44368 10254 44424
rect 10310 44368 10378 44424
rect 10434 44368 10502 44424
rect 10558 44368 10626 44424
rect 10682 44368 10750 44424
rect 10806 44368 10874 44424
rect 10930 44368 10998 44424
rect 11054 44368 11122 44424
rect 11178 44368 11246 44424
rect 11302 44368 11370 44424
rect 11426 44368 11494 44424
rect 11550 44368 11618 44424
rect 11674 44368 11742 44424
rect 11798 44368 11866 44424
rect 11922 44368 11990 44424
rect 12046 44368 12114 44424
rect 12170 44368 12180 44424
rect 10244 44300 12180 44368
rect 10244 44244 10254 44300
rect 10310 44244 10378 44300
rect 10434 44244 10502 44300
rect 10558 44244 10626 44300
rect 10682 44244 10750 44300
rect 10806 44244 10874 44300
rect 10930 44244 10998 44300
rect 11054 44244 11122 44300
rect 11178 44244 11246 44300
rect 11302 44244 11370 44300
rect 11426 44244 11494 44300
rect 11550 44244 11618 44300
rect 11674 44244 11742 44300
rect 11798 44244 11866 44300
rect 11922 44244 11990 44300
rect 12046 44244 12114 44300
rect 12170 44244 12180 44300
rect 10244 44176 12180 44244
rect 10244 44120 10254 44176
rect 10310 44120 10378 44176
rect 10434 44120 10502 44176
rect 10558 44120 10626 44176
rect 10682 44120 10750 44176
rect 10806 44120 10874 44176
rect 10930 44120 10998 44176
rect 11054 44120 11122 44176
rect 11178 44120 11246 44176
rect 11302 44120 11370 44176
rect 11426 44120 11494 44176
rect 11550 44120 11618 44176
rect 11674 44120 11742 44176
rect 11798 44120 11866 44176
rect 11922 44120 11990 44176
rect 12046 44120 12114 44176
rect 12170 44120 12180 44176
rect 10244 44052 12180 44120
rect 10244 43996 10254 44052
rect 10310 43996 10378 44052
rect 10434 43996 10502 44052
rect 10558 43996 10626 44052
rect 10682 43996 10750 44052
rect 10806 43996 10874 44052
rect 10930 43996 10998 44052
rect 11054 43996 11122 44052
rect 11178 43996 11246 44052
rect 11302 43996 11370 44052
rect 11426 43996 11494 44052
rect 11550 43996 11618 44052
rect 11674 43996 11742 44052
rect 11798 43996 11866 44052
rect 11922 43996 11990 44052
rect 12046 43996 12114 44052
rect 12170 43996 12180 44052
rect 10244 43928 12180 43996
rect 10244 43872 10254 43928
rect 10310 43872 10378 43928
rect 10434 43872 10502 43928
rect 10558 43872 10626 43928
rect 10682 43872 10750 43928
rect 10806 43872 10874 43928
rect 10930 43872 10998 43928
rect 11054 43872 11122 43928
rect 11178 43872 11246 43928
rect 11302 43872 11370 43928
rect 11426 43872 11494 43928
rect 11550 43872 11618 43928
rect 11674 43872 11742 43928
rect 11798 43872 11866 43928
rect 11922 43872 11990 43928
rect 12046 43872 12114 43928
rect 12170 43872 12180 43928
rect 10244 43804 12180 43872
rect 10244 43748 10254 43804
rect 10310 43748 10378 43804
rect 10434 43748 10502 43804
rect 10558 43748 10626 43804
rect 10682 43748 10750 43804
rect 10806 43748 10874 43804
rect 10930 43748 10998 43804
rect 11054 43748 11122 43804
rect 11178 43748 11246 43804
rect 11302 43748 11370 43804
rect 11426 43748 11494 43804
rect 11550 43748 11618 43804
rect 11674 43748 11742 43804
rect 11798 43748 11866 43804
rect 11922 43748 11990 43804
rect 12046 43748 12114 43804
rect 12170 43748 12180 43804
rect 10244 43680 12180 43748
rect 10244 43624 10254 43680
rect 10310 43624 10378 43680
rect 10434 43624 10502 43680
rect 10558 43624 10626 43680
rect 10682 43624 10750 43680
rect 10806 43624 10874 43680
rect 10930 43624 10998 43680
rect 11054 43624 11122 43680
rect 11178 43624 11246 43680
rect 11302 43624 11370 43680
rect 11426 43624 11494 43680
rect 11550 43624 11618 43680
rect 11674 43624 11742 43680
rect 11798 43624 11866 43680
rect 11922 43624 11990 43680
rect 12046 43624 12114 43680
rect 12170 43624 12180 43680
rect 10244 43556 12180 43624
rect 10244 43500 10254 43556
rect 10310 43500 10378 43556
rect 10434 43500 10502 43556
rect 10558 43500 10626 43556
rect 10682 43500 10750 43556
rect 10806 43500 10874 43556
rect 10930 43500 10998 43556
rect 11054 43500 11122 43556
rect 11178 43500 11246 43556
rect 11302 43500 11370 43556
rect 11426 43500 11494 43556
rect 11550 43500 11618 43556
rect 11674 43500 11742 43556
rect 11798 43500 11866 43556
rect 11922 43500 11990 43556
rect 12046 43500 12114 43556
rect 12170 43500 12180 43556
rect 10244 43432 12180 43500
rect 10244 43376 10254 43432
rect 10310 43376 10378 43432
rect 10434 43376 10502 43432
rect 10558 43376 10626 43432
rect 10682 43376 10750 43432
rect 10806 43376 10874 43432
rect 10930 43376 10998 43432
rect 11054 43376 11122 43432
rect 11178 43376 11246 43432
rect 11302 43376 11370 43432
rect 11426 43376 11494 43432
rect 11550 43376 11618 43432
rect 11674 43376 11742 43432
rect 11798 43376 11866 43432
rect 11922 43376 11990 43432
rect 12046 43376 12114 43432
rect 12170 43376 12180 43432
rect 10244 43308 12180 43376
rect 10244 43252 10254 43308
rect 10310 43252 10378 43308
rect 10434 43252 10502 43308
rect 10558 43252 10626 43308
rect 10682 43252 10750 43308
rect 10806 43252 10874 43308
rect 10930 43252 10998 43308
rect 11054 43252 11122 43308
rect 11178 43252 11246 43308
rect 11302 43252 11370 43308
rect 11426 43252 11494 43308
rect 11550 43252 11618 43308
rect 11674 43252 11742 43308
rect 11798 43252 11866 43308
rect 11922 43252 11990 43308
rect 12046 43252 12114 43308
rect 12170 43252 12180 43308
rect 10244 43242 12180 43252
rect 12861 44548 14673 44558
rect 12861 44492 12871 44548
rect 12927 44492 12995 44548
rect 13051 44492 13119 44548
rect 13175 44492 13243 44548
rect 13299 44492 13367 44548
rect 13423 44492 13491 44548
rect 13547 44492 13615 44548
rect 13671 44492 13739 44548
rect 13795 44492 13863 44548
rect 13919 44492 13987 44548
rect 14043 44492 14111 44548
rect 14167 44492 14235 44548
rect 14291 44492 14359 44548
rect 14415 44492 14483 44548
rect 14539 44492 14607 44548
rect 14663 44492 14673 44548
rect 12861 44424 14673 44492
rect 12861 44368 12871 44424
rect 12927 44368 12995 44424
rect 13051 44368 13119 44424
rect 13175 44368 13243 44424
rect 13299 44368 13367 44424
rect 13423 44368 13491 44424
rect 13547 44368 13615 44424
rect 13671 44368 13739 44424
rect 13795 44368 13863 44424
rect 13919 44368 13987 44424
rect 14043 44368 14111 44424
rect 14167 44368 14235 44424
rect 14291 44368 14359 44424
rect 14415 44368 14483 44424
rect 14539 44368 14607 44424
rect 14663 44368 14673 44424
rect 12861 44300 14673 44368
rect 12861 44244 12871 44300
rect 12927 44244 12995 44300
rect 13051 44244 13119 44300
rect 13175 44244 13243 44300
rect 13299 44244 13367 44300
rect 13423 44244 13491 44300
rect 13547 44244 13615 44300
rect 13671 44244 13739 44300
rect 13795 44244 13863 44300
rect 13919 44244 13987 44300
rect 14043 44244 14111 44300
rect 14167 44244 14235 44300
rect 14291 44244 14359 44300
rect 14415 44244 14483 44300
rect 14539 44244 14607 44300
rect 14663 44244 14673 44300
rect 12861 44176 14673 44244
rect 12861 44120 12871 44176
rect 12927 44120 12995 44176
rect 13051 44120 13119 44176
rect 13175 44120 13243 44176
rect 13299 44120 13367 44176
rect 13423 44120 13491 44176
rect 13547 44120 13615 44176
rect 13671 44120 13739 44176
rect 13795 44120 13863 44176
rect 13919 44120 13987 44176
rect 14043 44120 14111 44176
rect 14167 44120 14235 44176
rect 14291 44120 14359 44176
rect 14415 44120 14483 44176
rect 14539 44120 14607 44176
rect 14663 44120 14673 44176
rect 12861 44052 14673 44120
rect 12861 43996 12871 44052
rect 12927 43996 12995 44052
rect 13051 43996 13119 44052
rect 13175 43996 13243 44052
rect 13299 43996 13367 44052
rect 13423 43996 13491 44052
rect 13547 43996 13615 44052
rect 13671 43996 13739 44052
rect 13795 43996 13863 44052
rect 13919 43996 13987 44052
rect 14043 43996 14111 44052
rect 14167 43996 14235 44052
rect 14291 43996 14359 44052
rect 14415 43996 14483 44052
rect 14539 43996 14607 44052
rect 14663 43996 14673 44052
rect 12861 43928 14673 43996
rect 12861 43872 12871 43928
rect 12927 43872 12995 43928
rect 13051 43872 13119 43928
rect 13175 43872 13243 43928
rect 13299 43872 13367 43928
rect 13423 43872 13491 43928
rect 13547 43872 13615 43928
rect 13671 43872 13739 43928
rect 13795 43872 13863 43928
rect 13919 43872 13987 43928
rect 14043 43872 14111 43928
rect 14167 43872 14235 43928
rect 14291 43872 14359 43928
rect 14415 43872 14483 43928
rect 14539 43872 14607 43928
rect 14663 43872 14673 43928
rect 12861 43804 14673 43872
rect 12861 43748 12871 43804
rect 12927 43748 12995 43804
rect 13051 43748 13119 43804
rect 13175 43748 13243 43804
rect 13299 43748 13367 43804
rect 13423 43748 13491 43804
rect 13547 43748 13615 43804
rect 13671 43748 13739 43804
rect 13795 43748 13863 43804
rect 13919 43748 13987 43804
rect 14043 43748 14111 43804
rect 14167 43748 14235 43804
rect 14291 43748 14359 43804
rect 14415 43748 14483 43804
rect 14539 43748 14607 43804
rect 14663 43748 14673 43804
rect 12861 43680 14673 43748
rect 12861 43624 12871 43680
rect 12927 43624 12995 43680
rect 13051 43624 13119 43680
rect 13175 43624 13243 43680
rect 13299 43624 13367 43680
rect 13423 43624 13491 43680
rect 13547 43624 13615 43680
rect 13671 43624 13739 43680
rect 13795 43624 13863 43680
rect 13919 43624 13987 43680
rect 14043 43624 14111 43680
rect 14167 43624 14235 43680
rect 14291 43624 14359 43680
rect 14415 43624 14483 43680
rect 14539 43624 14607 43680
rect 14663 43624 14673 43680
rect 12861 43556 14673 43624
rect 12861 43500 12871 43556
rect 12927 43500 12995 43556
rect 13051 43500 13119 43556
rect 13175 43500 13243 43556
rect 13299 43500 13367 43556
rect 13423 43500 13491 43556
rect 13547 43500 13615 43556
rect 13671 43500 13739 43556
rect 13795 43500 13863 43556
rect 13919 43500 13987 43556
rect 14043 43500 14111 43556
rect 14167 43500 14235 43556
rect 14291 43500 14359 43556
rect 14415 43500 14483 43556
rect 14539 43500 14607 43556
rect 14663 43500 14673 43556
rect 12861 43432 14673 43500
rect 12861 43376 12871 43432
rect 12927 43376 12995 43432
rect 13051 43376 13119 43432
rect 13175 43376 13243 43432
rect 13299 43376 13367 43432
rect 13423 43376 13491 43432
rect 13547 43376 13615 43432
rect 13671 43376 13739 43432
rect 13795 43376 13863 43432
rect 13919 43376 13987 43432
rect 14043 43376 14111 43432
rect 14167 43376 14235 43432
rect 14291 43376 14359 43432
rect 14415 43376 14483 43432
rect 14539 43376 14607 43432
rect 14663 43376 14673 43432
rect 12861 43308 14673 43376
rect 12861 43252 12871 43308
rect 12927 43252 12995 43308
rect 13051 43252 13119 43308
rect 13175 43252 13243 43308
rect 13299 43252 13367 43308
rect 13423 43252 13491 43308
rect 13547 43252 13615 43308
rect 13671 43252 13739 43308
rect 13795 43252 13863 43308
rect 13919 43252 13987 43308
rect 14043 43252 14111 43308
rect 14167 43252 14235 43308
rect 14291 43252 14359 43308
rect 14415 43252 14483 43308
rect 14539 43252 14607 43308
rect 14663 43252 14673 43308
rect 12861 43242 14673 43252
rect 305 42948 2117 42958
rect 305 42892 315 42948
rect 371 42892 439 42948
rect 495 42892 563 42948
rect 619 42892 687 42948
rect 743 42892 811 42948
rect 867 42892 935 42948
rect 991 42892 1059 42948
rect 1115 42892 1183 42948
rect 1239 42892 1307 42948
rect 1363 42892 1431 42948
rect 1487 42892 1555 42948
rect 1611 42892 1679 42948
rect 1735 42892 1803 42948
rect 1859 42892 1927 42948
rect 1983 42892 2051 42948
rect 2107 42892 2117 42948
rect 305 42824 2117 42892
rect 305 42768 315 42824
rect 371 42768 439 42824
rect 495 42768 563 42824
rect 619 42768 687 42824
rect 743 42768 811 42824
rect 867 42768 935 42824
rect 991 42768 1059 42824
rect 1115 42768 1183 42824
rect 1239 42768 1307 42824
rect 1363 42768 1431 42824
rect 1487 42768 1555 42824
rect 1611 42768 1679 42824
rect 1735 42768 1803 42824
rect 1859 42768 1927 42824
rect 1983 42768 2051 42824
rect 2107 42768 2117 42824
rect 305 42700 2117 42768
rect 305 42644 315 42700
rect 371 42644 439 42700
rect 495 42644 563 42700
rect 619 42644 687 42700
rect 743 42644 811 42700
rect 867 42644 935 42700
rect 991 42644 1059 42700
rect 1115 42644 1183 42700
rect 1239 42644 1307 42700
rect 1363 42644 1431 42700
rect 1487 42644 1555 42700
rect 1611 42644 1679 42700
rect 1735 42644 1803 42700
rect 1859 42644 1927 42700
rect 1983 42644 2051 42700
rect 2107 42644 2117 42700
rect 305 42576 2117 42644
rect 305 42520 315 42576
rect 371 42520 439 42576
rect 495 42520 563 42576
rect 619 42520 687 42576
rect 743 42520 811 42576
rect 867 42520 935 42576
rect 991 42520 1059 42576
rect 1115 42520 1183 42576
rect 1239 42520 1307 42576
rect 1363 42520 1431 42576
rect 1487 42520 1555 42576
rect 1611 42520 1679 42576
rect 1735 42520 1803 42576
rect 1859 42520 1927 42576
rect 1983 42520 2051 42576
rect 2107 42520 2117 42576
rect 305 42452 2117 42520
rect 305 42396 315 42452
rect 371 42396 439 42452
rect 495 42396 563 42452
rect 619 42396 687 42452
rect 743 42396 811 42452
rect 867 42396 935 42452
rect 991 42396 1059 42452
rect 1115 42396 1183 42452
rect 1239 42396 1307 42452
rect 1363 42396 1431 42452
rect 1487 42396 1555 42452
rect 1611 42396 1679 42452
rect 1735 42396 1803 42452
rect 1859 42396 1927 42452
rect 1983 42396 2051 42452
rect 2107 42396 2117 42452
rect 305 42328 2117 42396
rect 305 42272 315 42328
rect 371 42272 439 42328
rect 495 42272 563 42328
rect 619 42272 687 42328
rect 743 42272 811 42328
rect 867 42272 935 42328
rect 991 42272 1059 42328
rect 1115 42272 1183 42328
rect 1239 42272 1307 42328
rect 1363 42272 1431 42328
rect 1487 42272 1555 42328
rect 1611 42272 1679 42328
rect 1735 42272 1803 42328
rect 1859 42272 1927 42328
rect 1983 42272 2051 42328
rect 2107 42272 2117 42328
rect 305 42204 2117 42272
rect 305 42148 315 42204
rect 371 42148 439 42204
rect 495 42148 563 42204
rect 619 42148 687 42204
rect 743 42148 811 42204
rect 867 42148 935 42204
rect 991 42148 1059 42204
rect 1115 42148 1183 42204
rect 1239 42148 1307 42204
rect 1363 42148 1431 42204
rect 1487 42148 1555 42204
rect 1611 42148 1679 42204
rect 1735 42148 1803 42204
rect 1859 42148 1927 42204
rect 1983 42148 2051 42204
rect 2107 42148 2117 42204
rect 305 42080 2117 42148
rect 305 42024 315 42080
rect 371 42024 439 42080
rect 495 42024 563 42080
rect 619 42024 687 42080
rect 743 42024 811 42080
rect 867 42024 935 42080
rect 991 42024 1059 42080
rect 1115 42024 1183 42080
rect 1239 42024 1307 42080
rect 1363 42024 1431 42080
rect 1487 42024 1555 42080
rect 1611 42024 1679 42080
rect 1735 42024 1803 42080
rect 1859 42024 1927 42080
rect 1983 42024 2051 42080
rect 2107 42024 2117 42080
rect 305 41956 2117 42024
rect 305 41900 315 41956
rect 371 41900 439 41956
rect 495 41900 563 41956
rect 619 41900 687 41956
rect 743 41900 811 41956
rect 867 41900 935 41956
rect 991 41900 1059 41956
rect 1115 41900 1183 41956
rect 1239 41900 1307 41956
rect 1363 41900 1431 41956
rect 1487 41900 1555 41956
rect 1611 41900 1679 41956
rect 1735 41900 1803 41956
rect 1859 41900 1927 41956
rect 1983 41900 2051 41956
rect 2107 41900 2117 41956
rect 305 41832 2117 41900
rect 305 41776 315 41832
rect 371 41776 439 41832
rect 495 41776 563 41832
rect 619 41776 687 41832
rect 743 41776 811 41832
rect 867 41776 935 41832
rect 991 41776 1059 41832
rect 1115 41776 1183 41832
rect 1239 41776 1307 41832
rect 1363 41776 1431 41832
rect 1487 41776 1555 41832
rect 1611 41776 1679 41832
rect 1735 41776 1803 41832
rect 1859 41776 1927 41832
rect 1983 41776 2051 41832
rect 2107 41776 2117 41832
rect 305 41708 2117 41776
rect 305 41652 315 41708
rect 371 41652 439 41708
rect 495 41652 563 41708
rect 619 41652 687 41708
rect 743 41652 811 41708
rect 867 41652 935 41708
rect 991 41652 1059 41708
rect 1115 41652 1183 41708
rect 1239 41652 1307 41708
rect 1363 41652 1431 41708
rect 1487 41652 1555 41708
rect 1611 41652 1679 41708
rect 1735 41652 1803 41708
rect 1859 41652 1927 41708
rect 1983 41652 2051 41708
rect 2107 41652 2117 41708
rect 305 41642 2117 41652
rect 2798 42948 4734 42958
rect 2798 42892 2808 42948
rect 2864 42892 2932 42948
rect 2988 42892 3056 42948
rect 3112 42892 3180 42948
rect 3236 42892 3304 42948
rect 3360 42892 3428 42948
rect 3484 42892 3552 42948
rect 3608 42892 3676 42948
rect 3732 42892 3800 42948
rect 3856 42892 3924 42948
rect 3980 42892 4048 42948
rect 4104 42892 4172 42948
rect 4228 42892 4296 42948
rect 4352 42892 4420 42948
rect 4476 42892 4544 42948
rect 4600 42892 4668 42948
rect 4724 42892 4734 42948
rect 2798 42824 4734 42892
rect 2798 42768 2808 42824
rect 2864 42768 2932 42824
rect 2988 42768 3056 42824
rect 3112 42768 3180 42824
rect 3236 42768 3304 42824
rect 3360 42768 3428 42824
rect 3484 42768 3552 42824
rect 3608 42768 3676 42824
rect 3732 42768 3800 42824
rect 3856 42768 3924 42824
rect 3980 42768 4048 42824
rect 4104 42768 4172 42824
rect 4228 42768 4296 42824
rect 4352 42768 4420 42824
rect 4476 42768 4544 42824
rect 4600 42768 4668 42824
rect 4724 42768 4734 42824
rect 2798 42700 4734 42768
rect 2798 42644 2808 42700
rect 2864 42644 2932 42700
rect 2988 42644 3056 42700
rect 3112 42644 3180 42700
rect 3236 42644 3304 42700
rect 3360 42644 3428 42700
rect 3484 42644 3552 42700
rect 3608 42644 3676 42700
rect 3732 42644 3800 42700
rect 3856 42644 3924 42700
rect 3980 42644 4048 42700
rect 4104 42644 4172 42700
rect 4228 42644 4296 42700
rect 4352 42644 4420 42700
rect 4476 42644 4544 42700
rect 4600 42644 4668 42700
rect 4724 42644 4734 42700
rect 2798 42576 4734 42644
rect 2798 42520 2808 42576
rect 2864 42520 2932 42576
rect 2988 42520 3056 42576
rect 3112 42520 3180 42576
rect 3236 42520 3304 42576
rect 3360 42520 3428 42576
rect 3484 42520 3552 42576
rect 3608 42520 3676 42576
rect 3732 42520 3800 42576
rect 3856 42520 3924 42576
rect 3980 42520 4048 42576
rect 4104 42520 4172 42576
rect 4228 42520 4296 42576
rect 4352 42520 4420 42576
rect 4476 42520 4544 42576
rect 4600 42520 4668 42576
rect 4724 42520 4734 42576
rect 2798 42452 4734 42520
rect 2798 42396 2808 42452
rect 2864 42396 2932 42452
rect 2988 42396 3056 42452
rect 3112 42396 3180 42452
rect 3236 42396 3304 42452
rect 3360 42396 3428 42452
rect 3484 42396 3552 42452
rect 3608 42396 3676 42452
rect 3732 42396 3800 42452
rect 3856 42396 3924 42452
rect 3980 42396 4048 42452
rect 4104 42396 4172 42452
rect 4228 42396 4296 42452
rect 4352 42396 4420 42452
rect 4476 42396 4544 42452
rect 4600 42396 4668 42452
rect 4724 42396 4734 42452
rect 2798 42328 4734 42396
rect 2798 42272 2808 42328
rect 2864 42272 2932 42328
rect 2988 42272 3056 42328
rect 3112 42272 3180 42328
rect 3236 42272 3304 42328
rect 3360 42272 3428 42328
rect 3484 42272 3552 42328
rect 3608 42272 3676 42328
rect 3732 42272 3800 42328
rect 3856 42272 3924 42328
rect 3980 42272 4048 42328
rect 4104 42272 4172 42328
rect 4228 42272 4296 42328
rect 4352 42272 4420 42328
rect 4476 42272 4544 42328
rect 4600 42272 4668 42328
rect 4724 42272 4734 42328
rect 2798 42204 4734 42272
rect 2798 42148 2808 42204
rect 2864 42148 2932 42204
rect 2988 42148 3056 42204
rect 3112 42148 3180 42204
rect 3236 42148 3304 42204
rect 3360 42148 3428 42204
rect 3484 42148 3552 42204
rect 3608 42148 3676 42204
rect 3732 42148 3800 42204
rect 3856 42148 3924 42204
rect 3980 42148 4048 42204
rect 4104 42148 4172 42204
rect 4228 42148 4296 42204
rect 4352 42148 4420 42204
rect 4476 42148 4544 42204
rect 4600 42148 4668 42204
rect 4724 42148 4734 42204
rect 2798 42080 4734 42148
rect 2798 42024 2808 42080
rect 2864 42024 2932 42080
rect 2988 42024 3056 42080
rect 3112 42024 3180 42080
rect 3236 42024 3304 42080
rect 3360 42024 3428 42080
rect 3484 42024 3552 42080
rect 3608 42024 3676 42080
rect 3732 42024 3800 42080
rect 3856 42024 3924 42080
rect 3980 42024 4048 42080
rect 4104 42024 4172 42080
rect 4228 42024 4296 42080
rect 4352 42024 4420 42080
rect 4476 42024 4544 42080
rect 4600 42024 4668 42080
rect 4724 42024 4734 42080
rect 2798 41956 4734 42024
rect 2798 41900 2808 41956
rect 2864 41900 2932 41956
rect 2988 41900 3056 41956
rect 3112 41900 3180 41956
rect 3236 41900 3304 41956
rect 3360 41900 3428 41956
rect 3484 41900 3552 41956
rect 3608 41900 3676 41956
rect 3732 41900 3800 41956
rect 3856 41900 3924 41956
rect 3980 41900 4048 41956
rect 4104 41900 4172 41956
rect 4228 41900 4296 41956
rect 4352 41900 4420 41956
rect 4476 41900 4544 41956
rect 4600 41900 4668 41956
rect 4724 41900 4734 41956
rect 2798 41832 4734 41900
rect 2798 41776 2808 41832
rect 2864 41776 2932 41832
rect 2988 41776 3056 41832
rect 3112 41776 3180 41832
rect 3236 41776 3304 41832
rect 3360 41776 3428 41832
rect 3484 41776 3552 41832
rect 3608 41776 3676 41832
rect 3732 41776 3800 41832
rect 3856 41776 3924 41832
rect 3980 41776 4048 41832
rect 4104 41776 4172 41832
rect 4228 41776 4296 41832
rect 4352 41776 4420 41832
rect 4476 41776 4544 41832
rect 4600 41776 4668 41832
rect 4724 41776 4734 41832
rect 2798 41708 4734 41776
rect 2798 41652 2808 41708
rect 2864 41652 2932 41708
rect 2988 41652 3056 41708
rect 3112 41652 3180 41708
rect 3236 41652 3304 41708
rect 3360 41652 3428 41708
rect 3484 41652 3552 41708
rect 3608 41652 3676 41708
rect 3732 41652 3800 41708
rect 3856 41652 3924 41708
rect 3980 41652 4048 41708
rect 4104 41652 4172 41708
rect 4228 41652 4296 41708
rect 4352 41652 4420 41708
rect 4476 41652 4544 41708
rect 4600 41652 4668 41708
rect 4724 41652 4734 41708
rect 2798 41642 4734 41652
rect 5168 42948 7104 42958
rect 5168 42892 5178 42948
rect 5234 42892 5302 42948
rect 5358 42892 5426 42948
rect 5482 42892 5550 42948
rect 5606 42892 5674 42948
rect 5730 42892 5798 42948
rect 5854 42892 5922 42948
rect 5978 42892 6046 42948
rect 6102 42892 6170 42948
rect 6226 42892 6294 42948
rect 6350 42892 6418 42948
rect 6474 42892 6542 42948
rect 6598 42892 6666 42948
rect 6722 42892 6790 42948
rect 6846 42892 6914 42948
rect 6970 42892 7038 42948
rect 7094 42892 7104 42948
rect 5168 42824 7104 42892
rect 5168 42768 5178 42824
rect 5234 42768 5302 42824
rect 5358 42768 5426 42824
rect 5482 42768 5550 42824
rect 5606 42768 5674 42824
rect 5730 42768 5798 42824
rect 5854 42768 5922 42824
rect 5978 42768 6046 42824
rect 6102 42768 6170 42824
rect 6226 42768 6294 42824
rect 6350 42768 6418 42824
rect 6474 42768 6542 42824
rect 6598 42768 6666 42824
rect 6722 42768 6790 42824
rect 6846 42768 6914 42824
rect 6970 42768 7038 42824
rect 7094 42768 7104 42824
rect 5168 42700 7104 42768
rect 5168 42644 5178 42700
rect 5234 42644 5302 42700
rect 5358 42644 5426 42700
rect 5482 42644 5550 42700
rect 5606 42644 5674 42700
rect 5730 42644 5798 42700
rect 5854 42644 5922 42700
rect 5978 42644 6046 42700
rect 6102 42644 6170 42700
rect 6226 42644 6294 42700
rect 6350 42644 6418 42700
rect 6474 42644 6542 42700
rect 6598 42644 6666 42700
rect 6722 42644 6790 42700
rect 6846 42644 6914 42700
rect 6970 42644 7038 42700
rect 7094 42644 7104 42700
rect 5168 42576 7104 42644
rect 5168 42520 5178 42576
rect 5234 42520 5302 42576
rect 5358 42520 5426 42576
rect 5482 42520 5550 42576
rect 5606 42520 5674 42576
rect 5730 42520 5798 42576
rect 5854 42520 5922 42576
rect 5978 42520 6046 42576
rect 6102 42520 6170 42576
rect 6226 42520 6294 42576
rect 6350 42520 6418 42576
rect 6474 42520 6542 42576
rect 6598 42520 6666 42576
rect 6722 42520 6790 42576
rect 6846 42520 6914 42576
rect 6970 42520 7038 42576
rect 7094 42520 7104 42576
rect 5168 42452 7104 42520
rect 5168 42396 5178 42452
rect 5234 42396 5302 42452
rect 5358 42396 5426 42452
rect 5482 42396 5550 42452
rect 5606 42396 5674 42452
rect 5730 42396 5798 42452
rect 5854 42396 5922 42452
rect 5978 42396 6046 42452
rect 6102 42396 6170 42452
rect 6226 42396 6294 42452
rect 6350 42396 6418 42452
rect 6474 42396 6542 42452
rect 6598 42396 6666 42452
rect 6722 42396 6790 42452
rect 6846 42396 6914 42452
rect 6970 42396 7038 42452
rect 7094 42396 7104 42452
rect 5168 42328 7104 42396
rect 5168 42272 5178 42328
rect 5234 42272 5302 42328
rect 5358 42272 5426 42328
rect 5482 42272 5550 42328
rect 5606 42272 5674 42328
rect 5730 42272 5798 42328
rect 5854 42272 5922 42328
rect 5978 42272 6046 42328
rect 6102 42272 6170 42328
rect 6226 42272 6294 42328
rect 6350 42272 6418 42328
rect 6474 42272 6542 42328
rect 6598 42272 6666 42328
rect 6722 42272 6790 42328
rect 6846 42272 6914 42328
rect 6970 42272 7038 42328
rect 7094 42272 7104 42328
rect 5168 42204 7104 42272
rect 5168 42148 5178 42204
rect 5234 42148 5302 42204
rect 5358 42148 5426 42204
rect 5482 42148 5550 42204
rect 5606 42148 5674 42204
rect 5730 42148 5798 42204
rect 5854 42148 5922 42204
rect 5978 42148 6046 42204
rect 6102 42148 6170 42204
rect 6226 42148 6294 42204
rect 6350 42148 6418 42204
rect 6474 42148 6542 42204
rect 6598 42148 6666 42204
rect 6722 42148 6790 42204
rect 6846 42148 6914 42204
rect 6970 42148 7038 42204
rect 7094 42148 7104 42204
rect 5168 42080 7104 42148
rect 5168 42024 5178 42080
rect 5234 42024 5302 42080
rect 5358 42024 5426 42080
rect 5482 42024 5550 42080
rect 5606 42024 5674 42080
rect 5730 42024 5798 42080
rect 5854 42024 5922 42080
rect 5978 42024 6046 42080
rect 6102 42024 6170 42080
rect 6226 42024 6294 42080
rect 6350 42024 6418 42080
rect 6474 42024 6542 42080
rect 6598 42024 6666 42080
rect 6722 42024 6790 42080
rect 6846 42024 6914 42080
rect 6970 42024 7038 42080
rect 7094 42024 7104 42080
rect 5168 41956 7104 42024
rect 5168 41900 5178 41956
rect 5234 41900 5302 41956
rect 5358 41900 5426 41956
rect 5482 41900 5550 41956
rect 5606 41900 5674 41956
rect 5730 41900 5798 41956
rect 5854 41900 5922 41956
rect 5978 41900 6046 41956
rect 6102 41900 6170 41956
rect 6226 41900 6294 41956
rect 6350 41900 6418 41956
rect 6474 41900 6542 41956
rect 6598 41900 6666 41956
rect 6722 41900 6790 41956
rect 6846 41900 6914 41956
rect 6970 41900 7038 41956
rect 7094 41900 7104 41956
rect 5168 41832 7104 41900
rect 5168 41776 5178 41832
rect 5234 41776 5302 41832
rect 5358 41776 5426 41832
rect 5482 41776 5550 41832
rect 5606 41776 5674 41832
rect 5730 41776 5798 41832
rect 5854 41776 5922 41832
rect 5978 41776 6046 41832
rect 6102 41776 6170 41832
rect 6226 41776 6294 41832
rect 6350 41776 6418 41832
rect 6474 41776 6542 41832
rect 6598 41776 6666 41832
rect 6722 41776 6790 41832
rect 6846 41776 6914 41832
rect 6970 41776 7038 41832
rect 7094 41776 7104 41832
rect 5168 41708 7104 41776
rect 5168 41652 5178 41708
rect 5234 41652 5302 41708
rect 5358 41652 5426 41708
rect 5482 41652 5550 41708
rect 5606 41652 5674 41708
rect 5730 41652 5798 41708
rect 5854 41652 5922 41708
rect 5978 41652 6046 41708
rect 6102 41652 6170 41708
rect 6226 41652 6294 41708
rect 6350 41652 6418 41708
rect 6474 41652 6542 41708
rect 6598 41652 6666 41708
rect 6722 41652 6790 41708
rect 6846 41652 6914 41708
rect 6970 41652 7038 41708
rect 7094 41652 7104 41708
rect 5168 41642 7104 41652
rect 7874 42948 9810 42958
rect 7874 42892 7884 42948
rect 7940 42892 8008 42948
rect 8064 42892 8132 42948
rect 8188 42892 8256 42948
rect 8312 42892 8380 42948
rect 8436 42892 8504 42948
rect 8560 42892 8628 42948
rect 8684 42892 8752 42948
rect 8808 42892 8876 42948
rect 8932 42892 9000 42948
rect 9056 42892 9124 42948
rect 9180 42892 9248 42948
rect 9304 42892 9372 42948
rect 9428 42892 9496 42948
rect 9552 42892 9620 42948
rect 9676 42892 9744 42948
rect 9800 42892 9810 42948
rect 7874 42824 9810 42892
rect 7874 42768 7884 42824
rect 7940 42768 8008 42824
rect 8064 42768 8132 42824
rect 8188 42768 8256 42824
rect 8312 42768 8380 42824
rect 8436 42768 8504 42824
rect 8560 42768 8628 42824
rect 8684 42768 8752 42824
rect 8808 42768 8876 42824
rect 8932 42768 9000 42824
rect 9056 42768 9124 42824
rect 9180 42768 9248 42824
rect 9304 42768 9372 42824
rect 9428 42768 9496 42824
rect 9552 42768 9620 42824
rect 9676 42768 9744 42824
rect 9800 42768 9810 42824
rect 7874 42700 9810 42768
rect 7874 42644 7884 42700
rect 7940 42644 8008 42700
rect 8064 42644 8132 42700
rect 8188 42644 8256 42700
rect 8312 42644 8380 42700
rect 8436 42644 8504 42700
rect 8560 42644 8628 42700
rect 8684 42644 8752 42700
rect 8808 42644 8876 42700
rect 8932 42644 9000 42700
rect 9056 42644 9124 42700
rect 9180 42644 9248 42700
rect 9304 42644 9372 42700
rect 9428 42644 9496 42700
rect 9552 42644 9620 42700
rect 9676 42644 9744 42700
rect 9800 42644 9810 42700
rect 7874 42576 9810 42644
rect 7874 42520 7884 42576
rect 7940 42520 8008 42576
rect 8064 42520 8132 42576
rect 8188 42520 8256 42576
rect 8312 42520 8380 42576
rect 8436 42520 8504 42576
rect 8560 42520 8628 42576
rect 8684 42520 8752 42576
rect 8808 42520 8876 42576
rect 8932 42520 9000 42576
rect 9056 42520 9124 42576
rect 9180 42520 9248 42576
rect 9304 42520 9372 42576
rect 9428 42520 9496 42576
rect 9552 42520 9620 42576
rect 9676 42520 9744 42576
rect 9800 42520 9810 42576
rect 7874 42452 9810 42520
rect 7874 42396 7884 42452
rect 7940 42396 8008 42452
rect 8064 42396 8132 42452
rect 8188 42396 8256 42452
rect 8312 42396 8380 42452
rect 8436 42396 8504 42452
rect 8560 42396 8628 42452
rect 8684 42396 8752 42452
rect 8808 42396 8876 42452
rect 8932 42396 9000 42452
rect 9056 42396 9124 42452
rect 9180 42396 9248 42452
rect 9304 42396 9372 42452
rect 9428 42396 9496 42452
rect 9552 42396 9620 42452
rect 9676 42396 9744 42452
rect 9800 42396 9810 42452
rect 7874 42328 9810 42396
rect 7874 42272 7884 42328
rect 7940 42272 8008 42328
rect 8064 42272 8132 42328
rect 8188 42272 8256 42328
rect 8312 42272 8380 42328
rect 8436 42272 8504 42328
rect 8560 42272 8628 42328
rect 8684 42272 8752 42328
rect 8808 42272 8876 42328
rect 8932 42272 9000 42328
rect 9056 42272 9124 42328
rect 9180 42272 9248 42328
rect 9304 42272 9372 42328
rect 9428 42272 9496 42328
rect 9552 42272 9620 42328
rect 9676 42272 9744 42328
rect 9800 42272 9810 42328
rect 7874 42204 9810 42272
rect 7874 42148 7884 42204
rect 7940 42148 8008 42204
rect 8064 42148 8132 42204
rect 8188 42148 8256 42204
rect 8312 42148 8380 42204
rect 8436 42148 8504 42204
rect 8560 42148 8628 42204
rect 8684 42148 8752 42204
rect 8808 42148 8876 42204
rect 8932 42148 9000 42204
rect 9056 42148 9124 42204
rect 9180 42148 9248 42204
rect 9304 42148 9372 42204
rect 9428 42148 9496 42204
rect 9552 42148 9620 42204
rect 9676 42148 9744 42204
rect 9800 42148 9810 42204
rect 7874 42080 9810 42148
rect 7874 42024 7884 42080
rect 7940 42024 8008 42080
rect 8064 42024 8132 42080
rect 8188 42024 8256 42080
rect 8312 42024 8380 42080
rect 8436 42024 8504 42080
rect 8560 42024 8628 42080
rect 8684 42024 8752 42080
rect 8808 42024 8876 42080
rect 8932 42024 9000 42080
rect 9056 42024 9124 42080
rect 9180 42024 9248 42080
rect 9304 42024 9372 42080
rect 9428 42024 9496 42080
rect 9552 42024 9620 42080
rect 9676 42024 9744 42080
rect 9800 42024 9810 42080
rect 7874 41956 9810 42024
rect 7874 41900 7884 41956
rect 7940 41900 8008 41956
rect 8064 41900 8132 41956
rect 8188 41900 8256 41956
rect 8312 41900 8380 41956
rect 8436 41900 8504 41956
rect 8560 41900 8628 41956
rect 8684 41900 8752 41956
rect 8808 41900 8876 41956
rect 8932 41900 9000 41956
rect 9056 41900 9124 41956
rect 9180 41900 9248 41956
rect 9304 41900 9372 41956
rect 9428 41900 9496 41956
rect 9552 41900 9620 41956
rect 9676 41900 9744 41956
rect 9800 41900 9810 41956
rect 7874 41832 9810 41900
rect 7874 41776 7884 41832
rect 7940 41776 8008 41832
rect 8064 41776 8132 41832
rect 8188 41776 8256 41832
rect 8312 41776 8380 41832
rect 8436 41776 8504 41832
rect 8560 41776 8628 41832
rect 8684 41776 8752 41832
rect 8808 41776 8876 41832
rect 8932 41776 9000 41832
rect 9056 41776 9124 41832
rect 9180 41776 9248 41832
rect 9304 41776 9372 41832
rect 9428 41776 9496 41832
rect 9552 41776 9620 41832
rect 9676 41776 9744 41832
rect 9800 41776 9810 41832
rect 7874 41708 9810 41776
rect 7874 41652 7884 41708
rect 7940 41652 8008 41708
rect 8064 41652 8132 41708
rect 8188 41652 8256 41708
rect 8312 41652 8380 41708
rect 8436 41652 8504 41708
rect 8560 41652 8628 41708
rect 8684 41652 8752 41708
rect 8808 41652 8876 41708
rect 8932 41652 9000 41708
rect 9056 41652 9124 41708
rect 9180 41652 9248 41708
rect 9304 41652 9372 41708
rect 9428 41652 9496 41708
rect 9552 41652 9620 41708
rect 9676 41652 9744 41708
rect 9800 41652 9810 41708
rect 7874 41642 9810 41652
rect 10244 42948 12180 42958
rect 10244 42892 10254 42948
rect 10310 42892 10378 42948
rect 10434 42892 10502 42948
rect 10558 42892 10626 42948
rect 10682 42892 10750 42948
rect 10806 42892 10874 42948
rect 10930 42892 10998 42948
rect 11054 42892 11122 42948
rect 11178 42892 11246 42948
rect 11302 42892 11370 42948
rect 11426 42892 11494 42948
rect 11550 42892 11618 42948
rect 11674 42892 11742 42948
rect 11798 42892 11866 42948
rect 11922 42892 11990 42948
rect 12046 42892 12114 42948
rect 12170 42892 12180 42948
rect 10244 42824 12180 42892
rect 10244 42768 10254 42824
rect 10310 42768 10378 42824
rect 10434 42768 10502 42824
rect 10558 42768 10626 42824
rect 10682 42768 10750 42824
rect 10806 42768 10874 42824
rect 10930 42768 10998 42824
rect 11054 42768 11122 42824
rect 11178 42768 11246 42824
rect 11302 42768 11370 42824
rect 11426 42768 11494 42824
rect 11550 42768 11618 42824
rect 11674 42768 11742 42824
rect 11798 42768 11866 42824
rect 11922 42768 11990 42824
rect 12046 42768 12114 42824
rect 12170 42768 12180 42824
rect 10244 42700 12180 42768
rect 10244 42644 10254 42700
rect 10310 42644 10378 42700
rect 10434 42644 10502 42700
rect 10558 42644 10626 42700
rect 10682 42644 10750 42700
rect 10806 42644 10874 42700
rect 10930 42644 10998 42700
rect 11054 42644 11122 42700
rect 11178 42644 11246 42700
rect 11302 42644 11370 42700
rect 11426 42644 11494 42700
rect 11550 42644 11618 42700
rect 11674 42644 11742 42700
rect 11798 42644 11866 42700
rect 11922 42644 11990 42700
rect 12046 42644 12114 42700
rect 12170 42644 12180 42700
rect 10244 42576 12180 42644
rect 10244 42520 10254 42576
rect 10310 42520 10378 42576
rect 10434 42520 10502 42576
rect 10558 42520 10626 42576
rect 10682 42520 10750 42576
rect 10806 42520 10874 42576
rect 10930 42520 10998 42576
rect 11054 42520 11122 42576
rect 11178 42520 11246 42576
rect 11302 42520 11370 42576
rect 11426 42520 11494 42576
rect 11550 42520 11618 42576
rect 11674 42520 11742 42576
rect 11798 42520 11866 42576
rect 11922 42520 11990 42576
rect 12046 42520 12114 42576
rect 12170 42520 12180 42576
rect 10244 42452 12180 42520
rect 10244 42396 10254 42452
rect 10310 42396 10378 42452
rect 10434 42396 10502 42452
rect 10558 42396 10626 42452
rect 10682 42396 10750 42452
rect 10806 42396 10874 42452
rect 10930 42396 10998 42452
rect 11054 42396 11122 42452
rect 11178 42396 11246 42452
rect 11302 42396 11370 42452
rect 11426 42396 11494 42452
rect 11550 42396 11618 42452
rect 11674 42396 11742 42452
rect 11798 42396 11866 42452
rect 11922 42396 11990 42452
rect 12046 42396 12114 42452
rect 12170 42396 12180 42452
rect 10244 42328 12180 42396
rect 10244 42272 10254 42328
rect 10310 42272 10378 42328
rect 10434 42272 10502 42328
rect 10558 42272 10626 42328
rect 10682 42272 10750 42328
rect 10806 42272 10874 42328
rect 10930 42272 10998 42328
rect 11054 42272 11122 42328
rect 11178 42272 11246 42328
rect 11302 42272 11370 42328
rect 11426 42272 11494 42328
rect 11550 42272 11618 42328
rect 11674 42272 11742 42328
rect 11798 42272 11866 42328
rect 11922 42272 11990 42328
rect 12046 42272 12114 42328
rect 12170 42272 12180 42328
rect 10244 42204 12180 42272
rect 10244 42148 10254 42204
rect 10310 42148 10378 42204
rect 10434 42148 10502 42204
rect 10558 42148 10626 42204
rect 10682 42148 10750 42204
rect 10806 42148 10874 42204
rect 10930 42148 10998 42204
rect 11054 42148 11122 42204
rect 11178 42148 11246 42204
rect 11302 42148 11370 42204
rect 11426 42148 11494 42204
rect 11550 42148 11618 42204
rect 11674 42148 11742 42204
rect 11798 42148 11866 42204
rect 11922 42148 11990 42204
rect 12046 42148 12114 42204
rect 12170 42148 12180 42204
rect 10244 42080 12180 42148
rect 10244 42024 10254 42080
rect 10310 42024 10378 42080
rect 10434 42024 10502 42080
rect 10558 42024 10626 42080
rect 10682 42024 10750 42080
rect 10806 42024 10874 42080
rect 10930 42024 10998 42080
rect 11054 42024 11122 42080
rect 11178 42024 11246 42080
rect 11302 42024 11370 42080
rect 11426 42024 11494 42080
rect 11550 42024 11618 42080
rect 11674 42024 11742 42080
rect 11798 42024 11866 42080
rect 11922 42024 11990 42080
rect 12046 42024 12114 42080
rect 12170 42024 12180 42080
rect 10244 41956 12180 42024
rect 10244 41900 10254 41956
rect 10310 41900 10378 41956
rect 10434 41900 10502 41956
rect 10558 41900 10626 41956
rect 10682 41900 10750 41956
rect 10806 41900 10874 41956
rect 10930 41900 10998 41956
rect 11054 41900 11122 41956
rect 11178 41900 11246 41956
rect 11302 41900 11370 41956
rect 11426 41900 11494 41956
rect 11550 41900 11618 41956
rect 11674 41900 11742 41956
rect 11798 41900 11866 41956
rect 11922 41900 11990 41956
rect 12046 41900 12114 41956
rect 12170 41900 12180 41956
rect 10244 41832 12180 41900
rect 10244 41776 10254 41832
rect 10310 41776 10378 41832
rect 10434 41776 10502 41832
rect 10558 41776 10626 41832
rect 10682 41776 10750 41832
rect 10806 41776 10874 41832
rect 10930 41776 10998 41832
rect 11054 41776 11122 41832
rect 11178 41776 11246 41832
rect 11302 41776 11370 41832
rect 11426 41776 11494 41832
rect 11550 41776 11618 41832
rect 11674 41776 11742 41832
rect 11798 41776 11866 41832
rect 11922 41776 11990 41832
rect 12046 41776 12114 41832
rect 12170 41776 12180 41832
rect 10244 41708 12180 41776
rect 10244 41652 10254 41708
rect 10310 41652 10378 41708
rect 10434 41652 10502 41708
rect 10558 41652 10626 41708
rect 10682 41652 10750 41708
rect 10806 41652 10874 41708
rect 10930 41652 10998 41708
rect 11054 41652 11122 41708
rect 11178 41652 11246 41708
rect 11302 41652 11370 41708
rect 11426 41652 11494 41708
rect 11550 41652 11618 41708
rect 11674 41652 11742 41708
rect 11798 41652 11866 41708
rect 11922 41652 11990 41708
rect 12046 41652 12114 41708
rect 12170 41652 12180 41708
rect 10244 41642 12180 41652
rect 12861 42948 14673 42958
rect 12861 42892 12871 42948
rect 12927 42892 12995 42948
rect 13051 42892 13119 42948
rect 13175 42892 13243 42948
rect 13299 42892 13367 42948
rect 13423 42892 13491 42948
rect 13547 42892 13615 42948
rect 13671 42892 13739 42948
rect 13795 42892 13863 42948
rect 13919 42892 13987 42948
rect 14043 42892 14111 42948
rect 14167 42892 14235 42948
rect 14291 42892 14359 42948
rect 14415 42892 14483 42948
rect 14539 42892 14607 42948
rect 14663 42892 14673 42948
rect 12861 42824 14673 42892
rect 12861 42768 12871 42824
rect 12927 42768 12995 42824
rect 13051 42768 13119 42824
rect 13175 42768 13243 42824
rect 13299 42768 13367 42824
rect 13423 42768 13491 42824
rect 13547 42768 13615 42824
rect 13671 42768 13739 42824
rect 13795 42768 13863 42824
rect 13919 42768 13987 42824
rect 14043 42768 14111 42824
rect 14167 42768 14235 42824
rect 14291 42768 14359 42824
rect 14415 42768 14483 42824
rect 14539 42768 14607 42824
rect 14663 42768 14673 42824
rect 12861 42700 14673 42768
rect 12861 42644 12871 42700
rect 12927 42644 12995 42700
rect 13051 42644 13119 42700
rect 13175 42644 13243 42700
rect 13299 42644 13367 42700
rect 13423 42644 13491 42700
rect 13547 42644 13615 42700
rect 13671 42644 13739 42700
rect 13795 42644 13863 42700
rect 13919 42644 13987 42700
rect 14043 42644 14111 42700
rect 14167 42644 14235 42700
rect 14291 42644 14359 42700
rect 14415 42644 14483 42700
rect 14539 42644 14607 42700
rect 14663 42644 14673 42700
rect 12861 42576 14673 42644
rect 12861 42520 12871 42576
rect 12927 42520 12995 42576
rect 13051 42520 13119 42576
rect 13175 42520 13243 42576
rect 13299 42520 13367 42576
rect 13423 42520 13491 42576
rect 13547 42520 13615 42576
rect 13671 42520 13739 42576
rect 13795 42520 13863 42576
rect 13919 42520 13987 42576
rect 14043 42520 14111 42576
rect 14167 42520 14235 42576
rect 14291 42520 14359 42576
rect 14415 42520 14483 42576
rect 14539 42520 14607 42576
rect 14663 42520 14673 42576
rect 12861 42452 14673 42520
rect 12861 42396 12871 42452
rect 12927 42396 12995 42452
rect 13051 42396 13119 42452
rect 13175 42396 13243 42452
rect 13299 42396 13367 42452
rect 13423 42396 13491 42452
rect 13547 42396 13615 42452
rect 13671 42396 13739 42452
rect 13795 42396 13863 42452
rect 13919 42396 13987 42452
rect 14043 42396 14111 42452
rect 14167 42396 14235 42452
rect 14291 42396 14359 42452
rect 14415 42396 14483 42452
rect 14539 42396 14607 42452
rect 14663 42396 14673 42452
rect 12861 42328 14673 42396
rect 12861 42272 12871 42328
rect 12927 42272 12995 42328
rect 13051 42272 13119 42328
rect 13175 42272 13243 42328
rect 13299 42272 13367 42328
rect 13423 42272 13491 42328
rect 13547 42272 13615 42328
rect 13671 42272 13739 42328
rect 13795 42272 13863 42328
rect 13919 42272 13987 42328
rect 14043 42272 14111 42328
rect 14167 42272 14235 42328
rect 14291 42272 14359 42328
rect 14415 42272 14483 42328
rect 14539 42272 14607 42328
rect 14663 42272 14673 42328
rect 12861 42204 14673 42272
rect 12861 42148 12871 42204
rect 12927 42148 12995 42204
rect 13051 42148 13119 42204
rect 13175 42148 13243 42204
rect 13299 42148 13367 42204
rect 13423 42148 13491 42204
rect 13547 42148 13615 42204
rect 13671 42148 13739 42204
rect 13795 42148 13863 42204
rect 13919 42148 13987 42204
rect 14043 42148 14111 42204
rect 14167 42148 14235 42204
rect 14291 42148 14359 42204
rect 14415 42148 14483 42204
rect 14539 42148 14607 42204
rect 14663 42148 14673 42204
rect 12861 42080 14673 42148
rect 12861 42024 12871 42080
rect 12927 42024 12995 42080
rect 13051 42024 13119 42080
rect 13175 42024 13243 42080
rect 13299 42024 13367 42080
rect 13423 42024 13491 42080
rect 13547 42024 13615 42080
rect 13671 42024 13739 42080
rect 13795 42024 13863 42080
rect 13919 42024 13987 42080
rect 14043 42024 14111 42080
rect 14167 42024 14235 42080
rect 14291 42024 14359 42080
rect 14415 42024 14483 42080
rect 14539 42024 14607 42080
rect 14663 42024 14673 42080
rect 12861 41956 14673 42024
rect 12861 41900 12871 41956
rect 12927 41900 12995 41956
rect 13051 41900 13119 41956
rect 13175 41900 13243 41956
rect 13299 41900 13367 41956
rect 13423 41900 13491 41956
rect 13547 41900 13615 41956
rect 13671 41900 13739 41956
rect 13795 41900 13863 41956
rect 13919 41900 13987 41956
rect 14043 41900 14111 41956
rect 14167 41900 14235 41956
rect 14291 41900 14359 41956
rect 14415 41900 14483 41956
rect 14539 41900 14607 41956
rect 14663 41900 14673 41956
rect 12861 41832 14673 41900
rect 12861 41776 12871 41832
rect 12927 41776 12995 41832
rect 13051 41776 13119 41832
rect 13175 41776 13243 41832
rect 13299 41776 13367 41832
rect 13423 41776 13491 41832
rect 13547 41776 13615 41832
rect 13671 41776 13739 41832
rect 13795 41776 13863 41832
rect 13919 41776 13987 41832
rect 14043 41776 14111 41832
rect 14167 41776 14235 41832
rect 14291 41776 14359 41832
rect 14415 41776 14483 41832
rect 14539 41776 14607 41832
rect 14663 41776 14673 41832
rect 12861 41708 14673 41776
rect 12861 41652 12871 41708
rect 12927 41652 12995 41708
rect 13051 41652 13119 41708
rect 13175 41652 13243 41708
rect 13299 41652 13367 41708
rect 13423 41652 13491 41708
rect 13547 41652 13615 41708
rect 13671 41652 13739 41708
rect 13795 41652 13863 41708
rect 13919 41652 13987 41708
rect 14043 41652 14111 41708
rect 14167 41652 14235 41708
rect 14291 41652 14359 41708
rect 14415 41652 14483 41708
rect 14539 41652 14607 41708
rect 14663 41652 14673 41708
rect 12861 41642 14673 41652
rect 305 41348 2117 41358
rect 305 41292 315 41348
rect 371 41292 439 41348
rect 495 41292 563 41348
rect 619 41292 687 41348
rect 743 41292 811 41348
rect 867 41292 935 41348
rect 991 41292 1059 41348
rect 1115 41292 1183 41348
rect 1239 41292 1307 41348
rect 1363 41292 1431 41348
rect 1487 41292 1555 41348
rect 1611 41292 1679 41348
rect 1735 41292 1803 41348
rect 1859 41292 1927 41348
rect 1983 41292 2051 41348
rect 2107 41292 2117 41348
rect 305 41224 2117 41292
rect 305 41168 315 41224
rect 371 41168 439 41224
rect 495 41168 563 41224
rect 619 41168 687 41224
rect 743 41168 811 41224
rect 867 41168 935 41224
rect 991 41168 1059 41224
rect 1115 41168 1183 41224
rect 1239 41168 1307 41224
rect 1363 41168 1431 41224
rect 1487 41168 1555 41224
rect 1611 41168 1679 41224
rect 1735 41168 1803 41224
rect 1859 41168 1927 41224
rect 1983 41168 2051 41224
rect 2107 41168 2117 41224
rect 305 41100 2117 41168
rect 305 41044 315 41100
rect 371 41044 439 41100
rect 495 41044 563 41100
rect 619 41044 687 41100
rect 743 41044 811 41100
rect 867 41044 935 41100
rect 991 41044 1059 41100
rect 1115 41044 1183 41100
rect 1239 41044 1307 41100
rect 1363 41044 1431 41100
rect 1487 41044 1555 41100
rect 1611 41044 1679 41100
rect 1735 41044 1803 41100
rect 1859 41044 1927 41100
rect 1983 41044 2051 41100
rect 2107 41044 2117 41100
rect 305 40976 2117 41044
rect 305 40920 315 40976
rect 371 40920 439 40976
rect 495 40920 563 40976
rect 619 40920 687 40976
rect 743 40920 811 40976
rect 867 40920 935 40976
rect 991 40920 1059 40976
rect 1115 40920 1183 40976
rect 1239 40920 1307 40976
rect 1363 40920 1431 40976
rect 1487 40920 1555 40976
rect 1611 40920 1679 40976
rect 1735 40920 1803 40976
rect 1859 40920 1927 40976
rect 1983 40920 2051 40976
rect 2107 40920 2117 40976
rect 305 40852 2117 40920
rect 305 40796 315 40852
rect 371 40796 439 40852
rect 495 40796 563 40852
rect 619 40796 687 40852
rect 743 40796 811 40852
rect 867 40796 935 40852
rect 991 40796 1059 40852
rect 1115 40796 1183 40852
rect 1239 40796 1307 40852
rect 1363 40796 1431 40852
rect 1487 40796 1555 40852
rect 1611 40796 1679 40852
rect 1735 40796 1803 40852
rect 1859 40796 1927 40852
rect 1983 40796 2051 40852
rect 2107 40796 2117 40852
rect 305 40728 2117 40796
rect 305 40672 315 40728
rect 371 40672 439 40728
rect 495 40672 563 40728
rect 619 40672 687 40728
rect 743 40672 811 40728
rect 867 40672 935 40728
rect 991 40672 1059 40728
rect 1115 40672 1183 40728
rect 1239 40672 1307 40728
rect 1363 40672 1431 40728
rect 1487 40672 1555 40728
rect 1611 40672 1679 40728
rect 1735 40672 1803 40728
rect 1859 40672 1927 40728
rect 1983 40672 2051 40728
rect 2107 40672 2117 40728
rect 305 40604 2117 40672
rect 305 40548 315 40604
rect 371 40548 439 40604
rect 495 40548 563 40604
rect 619 40548 687 40604
rect 743 40548 811 40604
rect 867 40548 935 40604
rect 991 40548 1059 40604
rect 1115 40548 1183 40604
rect 1239 40548 1307 40604
rect 1363 40548 1431 40604
rect 1487 40548 1555 40604
rect 1611 40548 1679 40604
rect 1735 40548 1803 40604
rect 1859 40548 1927 40604
rect 1983 40548 2051 40604
rect 2107 40548 2117 40604
rect 305 40480 2117 40548
rect 305 40424 315 40480
rect 371 40424 439 40480
rect 495 40424 563 40480
rect 619 40424 687 40480
rect 743 40424 811 40480
rect 867 40424 935 40480
rect 991 40424 1059 40480
rect 1115 40424 1183 40480
rect 1239 40424 1307 40480
rect 1363 40424 1431 40480
rect 1487 40424 1555 40480
rect 1611 40424 1679 40480
rect 1735 40424 1803 40480
rect 1859 40424 1927 40480
rect 1983 40424 2051 40480
rect 2107 40424 2117 40480
rect 305 40356 2117 40424
rect 305 40300 315 40356
rect 371 40300 439 40356
rect 495 40300 563 40356
rect 619 40300 687 40356
rect 743 40300 811 40356
rect 867 40300 935 40356
rect 991 40300 1059 40356
rect 1115 40300 1183 40356
rect 1239 40300 1307 40356
rect 1363 40300 1431 40356
rect 1487 40300 1555 40356
rect 1611 40300 1679 40356
rect 1735 40300 1803 40356
rect 1859 40300 1927 40356
rect 1983 40300 2051 40356
rect 2107 40300 2117 40356
rect 305 40232 2117 40300
rect 305 40176 315 40232
rect 371 40176 439 40232
rect 495 40176 563 40232
rect 619 40176 687 40232
rect 743 40176 811 40232
rect 867 40176 935 40232
rect 991 40176 1059 40232
rect 1115 40176 1183 40232
rect 1239 40176 1307 40232
rect 1363 40176 1431 40232
rect 1487 40176 1555 40232
rect 1611 40176 1679 40232
rect 1735 40176 1803 40232
rect 1859 40176 1927 40232
rect 1983 40176 2051 40232
rect 2107 40176 2117 40232
rect 305 40108 2117 40176
rect 305 40052 315 40108
rect 371 40052 439 40108
rect 495 40052 563 40108
rect 619 40052 687 40108
rect 743 40052 811 40108
rect 867 40052 935 40108
rect 991 40052 1059 40108
rect 1115 40052 1183 40108
rect 1239 40052 1307 40108
rect 1363 40052 1431 40108
rect 1487 40052 1555 40108
rect 1611 40052 1679 40108
rect 1735 40052 1803 40108
rect 1859 40052 1927 40108
rect 1983 40052 2051 40108
rect 2107 40052 2117 40108
rect 305 40042 2117 40052
rect 2798 41348 4734 41358
rect 2798 41292 2808 41348
rect 2864 41292 2932 41348
rect 2988 41292 3056 41348
rect 3112 41292 3180 41348
rect 3236 41292 3304 41348
rect 3360 41292 3428 41348
rect 3484 41292 3552 41348
rect 3608 41292 3676 41348
rect 3732 41292 3800 41348
rect 3856 41292 3924 41348
rect 3980 41292 4048 41348
rect 4104 41292 4172 41348
rect 4228 41292 4296 41348
rect 4352 41292 4420 41348
rect 4476 41292 4544 41348
rect 4600 41292 4668 41348
rect 4724 41292 4734 41348
rect 2798 41224 4734 41292
rect 2798 41168 2808 41224
rect 2864 41168 2932 41224
rect 2988 41168 3056 41224
rect 3112 41168 3180 41224
rect 3236 41168 3304 41224
rect 3360 41168 3428 41224
rect 3484 41168 3552 41224
rect 3608 41168 3676 41224
rect 3732 41168 3800 41224
rect 3856 41168 3924 41224
rect 3980 41168 4048 41224
rect 4104 41168 4172 41224
rect 4228 41168 4296 41224
rect 4352 41168 4420 41224
rect 4476 41168 4544 41224
rect 4600 41168 4668 41224
rect 4724 41168 4734 41224
rect 2798 41100 4734 41168
rect 2798 41044 2808 41100
rect 2864 41044 2932 41100
rect 2988 41044 3056 41100
rect 3112 41044 3180 41100
rect 3236 41044 3304 41100
rect 3360 41044 3428 41100
rect 3484 41044 3552 41100
rect 3608 41044 3676 41100
rect 3732 41044 3800 41100
rect 3856 41044 3924 41100
rect 3980 41044 4048 41100
rect 4104 41044 4172 41100
rect 4228 41044 4296 41100
rect 4352 41044 4420 41100
rect 4476 41044 4544 41100
rect 4600 41044 4668 41100
rect 4724 41044 4734 41100
rect 2798 40976 4734 41044
rect 2798 40920 2808 40976
rect 2864 40920 2932 40976
rect 2988 40920 3056 40976
rect 3112 40920 3180 40976
rect 3236 40920 3304 40976
rect 3360 40920 3428 40976
rect 3484 40920 3552 40976
rect 3608 40920 3676 40976
rect 3732 40920 3800 40976
rect 3856 40920 3924 40976
rect 3980 40920 4048 40976
rect 4104 40920 4172 40976
rect 4228 40920 4296 40976
rect 4352 40920 4420 40976
rect 4476 40920 4544 40976
rect 4600 40920 4668 40976
rect 4724 40920 4734 40976
rect 2798 40852 4734 40920
rect 2798 40796 2808 40852
rect 2864 40796 2932 40852
rect 2988 40796 3056 40852
rect 3112 40796 3180 40852
rect 3236 40796 3304 40852
rect 3360 40796 3428 40852
rect 3484 40796 3552 40852
rect 3608 40796 3676 40852
rect 3732 40796 3800 40852
rect 3856 40796 3924 40852
rect 3980 40796 4048 40852
rect 4104 40796 4172 40852
rect 4228 40796 4296 40852
rect 4352 40796 4420 40852
rect 4476 40796 4544 40852
rect 4600 40796 4668 40852
rect 4724 40796 4734 40852
rect 2798 40728 4734 40796
rect 2798 40672 2808 40728
rect 2864 40672 2932 40728
rect 2988 40672 3056 40728
rect 3112 40672 3180 40728
rect 3236 40672 3304 40728
rect 3360 40672 3428 40728
rect 3484 40672 3552 40728
rect 3608 40672 3676 40728
rect 3732 40672 3800 40728
rect 3856 40672 3924 40728
rect 3980 40672 4048 40728
rect 4104 40672 4172 40728
rect 4228 40672 4296 40728
rect 4352 40672 4420 40728
rect 4476 40672 4544 40728
rect 4600 40672 4668 40728
rect 4724 40672 4734 40728
rect 2798 40604 4734 40672
rect 2798 40548 2808 40604
rect 2864 40548 2932 40604
rect 2988 40548 3056 40604
rect 3112 40548 3180 40604
rect 3236 40548 3304 40604
rect 3360 40548 3428 40604
rect 3484 40548 3552 40604
rect 3608 40548 3676 40604
rect 3732 40548 3800 40604
rect 3856 40548 3924 40604
rect 3980 40548 4048 40604
rect 4104 40548 4172 40604
rect 4228 40548 4296 40604
rect 4352 40548 4420 40604
rect 4476 40548 4544 40604
rect 4600 40548 4668 40604
rect 4724 40548 4734 40604
rect 2798 40480 4734 40548
rect 2798 40424 2808 40480
rect 2864 40424 2932 40480
rect 2988 40424 3056 40480
rect 3112 40424 3180 40480
rect 3236 40424 3304 40480
rect 3360 40424 3428 40480
rect 3484 40424 3552 40480
rect 3608 40424 3676 40480
rect 3732 40424 3800 40480
rect 3856 40424 3924 40480
rect 3980 40424 4048 40480
rect 4104 40424 4172 40480
rect 4228 40424 4296 40480
rect 4352 40424 4420 40480
rect 4476 40424 4544 40480
rect 4600 40424 4668 40480
rect 4724 40424 4734 40480
rect 2798 40356 4734 40424
rect 2798 40300 2808 40356
rect 2864 40300 2932 40356
rect 2988 40300 3056 40356
rect 3112 40300 3180 40356
rect 3236 40300 3304 40356
rect 3360 40300 3428 40356
rect 3484 40300 3552 40356
rect 3608 40300 3676 40356
rect 3732 40300 3800 40356
rect 3856 40300 3924 40356
rect 3980 40300 4048 40356
rect 4104 40300 4172 40356
rect 4228 40300 4296 40356
rect 4352 40300 4420 40356
rect 4476 40300 4544 40356
rect 4600 40300 4668 40356
rect 4724 40300 4734 40356
rect 2798 40232 4734 40300
rect 2798 40176 2808 40232
rect 2864 40176 2932 40232
rect 2988 40176 3056 40232
rect 3112 40176 3180 40232
rect 3236 40176 3304 40232
rect 3360 40176 3428 40232
rect 3484 40176 3552 40232
rect 3608 40176 3676 40232
rect 3732 40176 3800 40232
rect 3856 40176 3924 40232
rect 3980 40176 4048 40232
rect 4104 40176 4172 40232
rect 4228 40176 4296 40232
rect 4352 40176 4420 40232
rect 4476 40176 4544 40232
rect 4600 40176 4668 40232
rect 4724 40176 4734 40232
rect 2798 40108 4734 40176
rect 2798 40052 2808 40108
rect 2864 40052 2932 40108
rect 2988 40052 3056 40108
rect 3112 40052 3180 40108
rect 3236 40052 3304 40108
rect 3360 40052 3428 40108
rect 3484 40052 3552 40108
rect 3608 40052 3676 40108
rect 3732 40052 3800 40108
rect 3856 40052 3924 40108
rect 3980 40052 4048 40108
rect 4104 40052 4172 40108
rect 4228 40052 4296 40108
rect 4352 40052 4420 40108
rect 4476 40052 4544 40108
rect 4600 40052 4668 40108
rect 4724 40052 4734 40108
rect 2798 40042 4734 40052
rect 5168 41348 7104 41358
rect 5168 41292 5178 41348
rect 5234 41292 5302 41348
rect 5358 41292 5426 41348
rect 5482 41292 5550 41348
rect 5606 41292 5674 41348
rect 5730 41292 5798 41348
rect 5854 41292 5922 41348
rect 5978 41292 6046 41348
rect 6102 41292 6170 41348
rect 6226 41292 6294 41348
rect 6350 41292 6418 41348
rect 6474 41292 6542 41348
rect 6598 41292 6666 41348
rect 6722 41292 6790 41348
rect 6846 41292 6914 41348
rect 6970 41292 7038 41348
rect 7094 41292 7104 41348
rect 5168 41224 7104 41292
rect 5168 41168 5178 41224
rect 5234 41168 5302 41224
rect 5358 41168 5426 41224
rect 5482 41168 5550 41224
rect 5606 41168 5674 41224
rect 5730 41168 5798 41224
rect 5854 41168 5922 41224
rect 5978 41168 6046 41224
rect 6102 41168 6170 41224
rect 6226 41168 6294 41224
rect 6350 41168 6418 41224
rect 6474 41168 6542 41224
rect 6598 41168 6666 41224
rect 6722 41168 6790 41224
rect 6846 41168 6914 41224
rect 6970 41168 7038 41224
rect 7094 41168 7104 41224
rect 5168 41100 7104 41168
rect 5168 41044 5178 41100
rect 5234 41044 5302 41100
rect 5358 41044 5426 41100
rect 5482 41044 5550 41100
rect 5606 41044 5674 41100
rect 5730 41044 5798 41100
rect 5854 41044 5922 41100
rect 5978 41044 6046 41100
rect 6102 41044 6170 41100
rect 6226 41044 6294 41100
rect 6350 41044 6418 41100
rect 6474 41044 6542 41100
rect 6598 41044 6666 41100
rect 6722 41044 6790 41100
rect 6846 41044 6914 41100
rect 6970 41044 7038 41100
rect 7094 41044 7104 41100
rect 5168 40976 7104 41044
rect 5168 40920 5178 40976
rect 5234 40920 5302 40976
rect 5358 40920 5426 40976
rect 5482 40920 5550 40976
rect 5606 40920 5674 40976
rect 5730 40920 5798 40976
rect 5854 40920 5922 40976
rect 5978 40920 6046 40976
rect 6102 40920 6170 40976
rect 6226 40920 6294 40976
rect 6350 40920 6418 40976
rect 6474 40920 6542 40976
rect 6598 40920 6666 40976
rect 6722 40920 6790 40976
rect 6846 40920 6914 40976
rect 6970 40920 7038 40976
rect 7094 40920 7104 40976
rect 5168 40852 7104 40920
rect 5168 40796 5178 40852
rect 5234 40796 5302 40852
rect 5358 40796 5426 40852
rect 5482 40796 5550 40852
rect 5606 40796 5674 40852
rect 5730 40796 5798 40852
rect 5854 40796 5922 40852
rect 5978 40796 6046 40852
rect 6102 40796 6170 40852
rect 6226 40796 6294 40852
rect 6350 40796 6418 40852
rect 6474 40796 6542 40852
rect 6598 40796 6666 40852
rect 6722 40796 6790 40852
rect 6846 40796 6914 40852
rect 6970 40796 7038 40852
rect 7094 40796 7104 40852
rect 5168 40728 7104 40796
rect 5168 40672 5178 40728
rect 5234 40672 5302 40728
rect 5358 40672 5426 40728
rect 5482 40672 5550 40728
rect 5606 40672 5674 40728
rect 5730 40672 5798 40728
rect 5854 40672 5922 40728
rect 5978 40672 6046 40728
rect 6102 40672 6170 40728
rect 6226 40672 6294 40728
rect 6350 40672 6418 40728
rect 6474 40672 6542 40728
rect 6598 40672 6666 40728
rect 6722 40672 6790 40728
rect 6846 40672 6914 40728
rect 6970 40672 7038 40728
rect 7094 40672 7104 40728
rect 5168 40604 7104 40672
rect 5168 40548 5178 40604
rect 5234 40548 5302 40604
rect 5358 40548 5426 40604
rect 5482 40548 5550 40604
rect 5606 40548 5674 40604
rect 5730 40548 5798 40604
rect 5854 40548 5922 40604
rect 5978 40548 6046 40604
rect 6102 40548 6170 40604
rect 6226 40548 6294 40604
rect 6350 40548 6418 40604
rect 6474 40548 6542 40604
rect 6598 40548 6666 40604
rect 6722 40548 6790 40604
rect 6846 40548 6914 40604
rect 6970 40548 7038 40604
rect 7094 40548 7104 40604
rect 5168 40480 7104 40548
rect 5168 40424 5178 40480
rect 5234 40424 5302 40480
rect 5358 40424 5426 40480
rect 5482 40424 5550 40480
rect 5606 40424 5674 40480
rect 5730 40424 5798 40480
rect 5854 40424 5922 40480
rect 5978 40424 6046 40480
rect 6102 40424 6170 40480
rect 6226 40424 6294 40480
rect 6350 40424 6418 40480
rect 6474 40424 6542 40480
rect 6598 40424 6666 40480
rect 6722 40424 6790 40480
rect 6846 40424 6914 40480
rect 6970 40424 7038 40480
rect 7094 40424 7104 40480
rect 5168 40356 7104 40424
rect 5168 40300 5178 40356
rect 5234 40300 5302 40356
rect 5358 40300 5426 40356
rect 5482 40300 5550 40356
rect 5606 40300 5674 40356
rect 5730 40300 5798 40356
rect 5854 40300 5922 40356
rect 5978 40300 6046 40356
rect 6102 40300 6170 40356
rect 6226 40300 6294 40356
rect 6350 40300 6418 40356
rect 6474 40300 6542 40356
rect 6598 40300 6666 40356
rect 6722 40300 6790 40356
rect 6846 40300 6914 40356
rect 6970 40300 7038 40356
rect 7094 40300 7104 40356
rect 5168 40232 7104 40300
rect 5168 40176 5178 40232
rect 5234 40176 5302 40232
rect 5358 40176 5426 40232
rect 5482 40176 5550 40232
rect 5606 40176 5674 40232
rect 5730 40176 5798 40232
rect 5854 40176 5922 40232
rect 5978 40176 6046 40232
rect 6102 40176 6170 40232
rect 6226 40176 6294 40232
rect 6350 40176 6418 40232
rect 6474 40176 6542 40232
rect 6598 40176 6666 40232
rect 6722 40176 6790 40232
rect 6846 40176 6914 40232
rect 6970 40176 7038 40232
rect 7094 40176 7104 40232
rect 5168 40108 7104 40176
rect 5168 40052 5178 40108
rect 5234 40052 5302 40108
rect 5358 40052 5426 40108
rect 5482 40052 5550 40108
rect 5606 40052 5674 40108
rect 5730 40052 5798 40108
rect 5854 40052 5922 40108
rect 5978 40052 6046 40108
rect 6102 40052 6170 40108
rect 6226 40052 6294 40108
rect 6350 40052 6418 40108
rect 6474 40052 6542 40108
rect 6598 40052 6666 40108
rect 6722 40052 6790 40108
rect 6846 40052 6914 40108
rect 6970 40052 7038 40108
rect 7094 40052 7104 40108
rect 5168 40042 7104 40052
rect 7874 41348 9810 41358
rect 7874 41292 7884 41348
rect 7940 41292 8008 41348
rect 8064 41292 8132 41348
rect 8188 41292 8256 41348
rect 8312 41292 8380 41348
rect 8436 41292 8504 41348
rect 8560 41292 8628 41348
rect 8684 41292 8752 41348
rect 8808 41292 8876 41348
rect 8932 41292 9000 41348
rect 9056 41292 9124 41348
rect 9180 41292 9248 41348
rect 9304 41292 9372 41348
rect 9428 41292 9496 41348
rect 9552 41292 9620 41348
rect 9676 41292 9744 41348
rect 9800 41292 9810 41348
rect 7874 41224 9810 41292
rect 7874 41168 7884 41224
rect 7940 41168 8008 41224
rect 8064 41168 8132 41224
rect 8188 41168 8256 41224
rect 8312 41168 8380 41224
rect 8436 41168 8504 41224
rect 8560 41168 8628 41224
rect 8684 41168 8752 41224
rect 8808 41168 8876 41224
rect 8932 41168 9000 41224
rect 9056 41168 9124 41224
rect 9180 41168 9248 41224
rect 9304 41168 9372 41224
rect 9428 41168 9496 41224
rect 9552 41168 9620 41224
rect 9676 41168 9744 41224
rect 9800 41168 9810 41224
rect 7874 41100 9810 41168
rect 7874 41044 7884 41100
rect 7940 41044 8008 41100
rect 8064 41044 8132 41100
rect 8188 41044 8256 41100
rect 8312 41044 8380 41100
rect 8436 41044 8504 41100
rect 8560 41044 8628 41100
rect 8684 41044 8752 41100
rect 8808 41044 8876 41100
rect 8932 41044 9000 41100
rect 9056 41044 9124 41100
rect 9180 41044 9248 41100
rect 9304 41044 9372 41100
rect 9428 41044 9496 41100
rect 9552 41044 9620 41100
rect 9676 41044 9744 41100
rect 9800 41044 9810 41100
rect 7874 40976 9810 41044
rect 7874 40920 7884 40976
rect 7940 40920 8008 40976
rect 8064 40920 8132 40976
rect 8188 40920 8256 40976
rect 8312 40920 8380 40976
rect 8436 40920 8504 40976
rect 8560 40920 8628 40976
rect 8684 40920 8752 40976
rect 8808 40920 8876 40976
rect 8932 40920 9000 40976
rect 9056 40920 9124 40976
rect 9180 40920 9248 40976
rect 9304 40920 9372 40976
rect 9428 40920 9496 40976
rect 9552 40920 9620 40976
rect 9676 40920 9744 40976
rect 9800 40920 9810 40976
rect 7874 40852 9810 40920
rect 7874 40796 7884 40852
rect 7940 40796 8008 40852
rect 8064 40796 8132 40852
rect 8188 40796 8256 40852
rect 8312 40796 8380 40852
rect 8436 40796 8504 40852
rect 8560 40796 8628 40852
rect 8684 40796 8752 40852
rect 8808 40796 8876 40852
rect 8932 40796 9000 40852
rect 9056 40796 9124 40852
rect 9180 40796 9248 40852
rect 9304 40796 9372 40852
rect 9428 40796 9496 40852
rect 9552 40796 9620 40852
rect 9676 40796 9744 40852
rect 9800 40796 9810 40852
rect 7874 40728 9810 40796
rect 7874 40672 7884 40728
rect 7940 40672 8008 40728
rect 8064 40672 8132 40728
rect 8188 40672 8256 40728
rect 8312 40672 8380 40728
rect 8436 40672 8504 40728
rect 8560 40672 8628 40728
rect 8684 40672 8752 40728
rect 8808 40672 8876 40728
rect 8932 40672 9000 40728
rect 9056 40672 9124 40728
rect 9180 40672 9248 40728
rect 9304 40672 9372 40728
rect 9428 40672 9496 40728
rect 9552 40672 9620 40728
rect 9676 40672 9744 40728
rect 9800 40672 9810 40728
rect 7874 40604 9810 40672
rect 7874 40548 7884 40604
rect 7940 40548 8008 40604
rect 8064 40548 8132 40604
rect 8188 40548 8256 40604
rect 8312 40548 8380 40604
rect 8436 40548 8504 40604
rect 8560 40548 8628 40604
rect 8684 40548 8752 40604
rect 8808 40548 8876 40604
rect 8932 40548 9000 40604
rect 9056 40548 9124 40604
rect 9180 40548 9248 40604
rect 9304 40548 9372 40604
rect 9428 40548 9496 40604
rect 9552 40548 9620 40604
rect 9676 40548 9744 40604
rect 9800 40548 9810 40604
rect 7874 40480 9810 40548
rect 7874 40424 7884 40480
rect 7940 40424 8008 40480
rect 8064 40424 8132 40480
rect 8188 40424 8256 40480
rect 8312 40424 8380 40480
rect 8436 40424 8504 40480
rect 8560 40424 8628 40480
rect 8684 40424 8752 40480
rect 8808 40424 8876 40480
rect 8932 40424 9000 40480
rect 9056 40424 9124 40480
rect 9180 40424 9248 40480
rect 9304 40424 9372 40480
rect 9428 40424 9496 40480
rect 9552 40424 9620 40480
rect 9676 40424 9744 40480
rect 9800 40424 9810 40480
rect 7874 40356 9810 40424
rect 7874 40300 7884 40356
rect 7940 40300 8008 40356
rect 8064 40300 8132 40356
rect 8188 40300 8256 40356
rect 8312 40300 8380 40356
rect 8436 40300 8504 40356
rect 8560 40300 8628 40356
rect 8684 40300 8752 40356
rect 8808 40300 8876 40356
rect 8932 40300 9000 40356
rect 9056 40300 9124 40356
rect 9180 40300 9248 40356
rect 9304 40300 9372 40356
rect 9428 40300 9496 40356
rect 9552 40300 9620 40356
rect 9676 40300 9744 40356
rect 9800 40300 9810 40356
rect 7874 40232 9810 40300
rect 7874 40176 7884 40232
rect 7940 40176 8008 40232
rect 8064 40176 8132 40232
rect 8188 40176 8256 40232
rect 8312 40176 8380 40232
rect 8436 40176 8504 40232
rect 8560 40176 8628 40232
rect 8684 40176 8752 40232
rect 8808 40176 8876 40232
rect 8932 40176 9000 40232
rect 9056 40176 9124 40232
rect 9180 40176 9248 40232
rect 9304 40176 9372 40232
rect 9428 40176 9496 40232
rect 9552 40176 9620 40232
rect 9676 40176 9744 40232
rect 9800 40176 9810 40232
rect 7874 40108 9810 40176
rect 7874 40052 7884 40108
rect 7940 40052 8008 40108
rect 8064 40052 8132 40108
rect 8188 40052 8256 40108
rect 8312 40052 8380 40108
rect 8436 40052 8504 40108
rect 8560 40052 8628 40108
rect 8684 40052 8752 40108
rect 8808 40052 8876 40108
rect 8932 40052 9000 40108
rect 9056 40052 9124 40108
rect 9180 40052 9248 40108
rect 9304 40052 9372 40108
rect 9428 40052 9496 40108
rect 9552 40052 9620 40108
rect 9676 40052 9744 40108
rect 9800 40052 9810 40108
rect 7874 40042 9810 40052
rect 10244 41348 12180 41358
rect 10244 41292 10254 41348
rect 10310 41292 10378 41348
rect 10434 41292 10502 41348
rect 10558 41292 10626 41348
rect 10682 41292 10750 41348
rect 10806 41292 10874 41348
rect 10930 41292 10998 41348
rect 11054 41292 11122 41348
rect 11178 41292 11246 41348
rect 11302 41292 11370 41348
rect 11426 41292 11494 41348
rect 11550 41292 11618 41348
rect 11674 41292 11742 41348
rect 11798 41292 11866 41348
rect 11922 41292 11990 41348
rect 12046 41292 12114 41348
rect 12170 41292 12180 41348
rect 10244 41224 12180 41292
rect 10244 41168 10254 41224
rect 10310 41168 10378 41224
rect 10434 41168 10502 41224
rect 10558 41168 10626 41224
rect 10682 41168 10750 41224
rect 10806 41168 10874 41224
rect 10930 41168 10998 41224
rect 11054 41168 11122 41224
rect 11178 41168 11246 41224
rect 11302 41168 11370 41224
rect 11426 41168 11494 41224
rect 11550 41168 11618 41224
rect 11674 41168 11742 41224
rect 11798 41168 11866 41224
rect 11922 41168 11990 41224
rect 12046 41168 12114 41224
rect 12170 41168 12180 41224
rect 10244 41100 12180 41168
rect 10244 41044 10254 41100
rect 10310 41044 10378 41100
rect 10434 41044 10502 41100
rect 10558 41044 10626 41100
rect 10682 41044 10750 41100
rect 10806 41044 10874 41100
rect 10930 41044 10998 41100
rect 11054 41044 11122 41100
rect 11178 41044 11246 41100
rect 11302 41044 11370 41100
rect 11426 41044 11494 41100
rect 11550 41044 11618 41100
rect 11674 41044 11742 41100
rect 11798 41044 11866 41100
rect 11922 41044 11990 41100
rect 12046 41044 12114 41100
rect 12170 41044 12180 41100
rect 10244 40976 12180 41044
rect 10244 40920 10254 40976
rect 10310 40920 10378 40976
rect 10434 40920 10502 40976
rect 10558 40920 10626 40976
rect 10682 40920 10750 40976
rect 10806 40920 10874 40976
rect 10930 40920 10998 40976
rect 11054 40920 11122 40976
rect 11178 40920 11246 40976
rect 11302 40920 11370 40976
rect 11426 40920 11494 40976
rect 11550 40920 11618 40976
rect 11674 40920 11742 40976
rect 11798 40920 11866 40976
rect 11922 40920 11990 40976
rect 12046 40920 12114 40976
rect 12170 40920 12180 40976
rect 10244 40852 12180 40920
rect 10244 40796 10254 40852
rect 10310 40796 10378 40852
rect 10434 40796 10502 40852
rect 10558 40796 10626 40852
rect 10682 40796 10750 40852
rect 10806 40796 10874 40852
rect 10930 40796 10998 40852
rect 11054 40796 11122 40852
rect 11178 40796 11246 40852
rect 11302 40796 11370 40852
rect 11426 40796 11494 40852
rect 11550 40796 11618 40852
rect 11674 40796 11742 40852
rect 11798 40796 11866 40852
rect 11922 40796 11990 40852
rect 12046 40796 12114 40852
rect 12170 40796 12180 40852
rect 10244 40728 12180 40796
rect 10244 40672 10254 40728
rect 10310 40672 10378 40728
rect 10434 40672 10502 40728
rect 10558 40672 10626 40728
rect 10682 40672 10750 40728
rect 10806 40672 10874 40728
rect 10930 40672 10998 40728
rect 11054 40672 11122 40728
rect 11178 40672 11246 40728
rect 11302 40672 11370 40728
rect 11426 40672 11494 40728
rect 11550 40672 11618 40728
rect 11674 40672 11742 40728
rect 11798 40672 11866 40728
rect 11922 40672 11990 40728
rect 12046 40672 12114 40728
rect 12170 40672 12180 40728
rect 10244 40604 12180 40672
rect 10244 40548 10254 40604
rect 10310 40548 10378 40604
rect 10434 40548 10502 40604
rect 10558 40548 10626 40604
rect 10682 40548 10750 40604
rect 10806 40548 10874 40604
rect 10930 40548 10998 40604
rect 11054 40548 11122 40604
rect 11178 40548 11246 40604
rect 11302 40548 11370 40604
rect 11426 40548 11494 40604
rect 11550 40548 11618 40604
rect 11674 40548 11742 40604
rect 11798 40548 11866 40604
rect 11922 40548 11990 40604
rect 12046 40548 12114 40604
rect 12170 40548 12180 40604
rect 10244 40480 12180 40548
rect 10244 40424 10254 40480
rect 10310 40424 10378 40480
rect 10434 40424 10502 40480
rect 10558 40424 10626 40480
rect 10682 40424 10750 40480
rect 10806 40424 10874 40480
rect 10930 40424 10998 40480
rect 11054 40424 11122 40480
rect 11178 40424 11246 40480
rect 11302 40424 11370 40480
rect 11426 40424 11494 40480
rect 11550 40424 11618 40480
rect 11674 40424 11742 40480
rect 11798 40424 11866 40480
rect 11922 40424 11990 40480
rect 12046 40424 12114 40480
rect 12170 40424 12180 40480
rect 10244 40356 12180 40424
rect 10244 40300 10254 40356
rect 10310 40300 10378 40356
rect 10434 40300 10502 40356
rect 10558 40300 10626 40356
rect 10682 40300 10750 40356
rect 10806 40300 10874 40356
rect 10930 40300 10998 40356
rect 11054 40300 11122 40356
rect 11178 40300 11246 40356
rect 11302 40300 11370 40356
rect 11426 40300 11494 40356
rect 11550 40300 11618 40356
rect 11674 40300 11742 40356
rect 11798 40300 11866 40356
rect 11922 40300 11990 40356
rect 12046 40300 12114 40356
rect 12170 40300 12180 40356
rect 10244 40232 12180 40300
rect 10244 40176 10254 40232
rect 10310 40176 10378 40232
rect 10434 40176 10502 40232
rect 10558 40176 10626 40232
rect 10682 40176 10750 40232
rect 10806 40176 10874 40232
rect 10930 40176 10998 40232
rect 11054 40176 11122 40232
rect 11178 40176 11246 40232
rect 11302 40176 11370 40232
rect 11426 40176 11494 40232
rect 11550 40176 11618 40232
rect 11674 40176 11742 40232
rect 11798 40176 11866 40232
rect 11922 40176 11990 40232
rect 12046 40176 12114 40232
rect 12170 40176 12180 40232
rect 10244 40108 12180 40176
rect 10244 40052 10254 40108
rect 10310 40052 10378 40108
rect 10434 40052 10502 40108
rect 10558 40052 10626 40108
rect 10682 40052 10750 40108
rect 10806 40052 10874 40108
rect 10930 40052 10998 40108
rect 11054 40052 11122 40108
rect 11178 40052 11246 40108
rect 11302 40052 11370 40108
rect 11426 40052 11494 40108
rect 11550 40052 11618 40108
rect 11674 40052 11742 40108
rect 11798 40052 11866 40108
rect 11922 40052 11990 40108
rect 12046 40052 12114 40108
rect 12170 40052 12180 40108
rect 10244 40042 12180 40052
rect 12861 41348 14673 41358
rect 12861 41292 12871 41348
rect 12927 41292 12995 41348
rect 13051 41292 13119 41348
rect 13175 41292 13243 41348
rect 13299 41292 13367 41348
rect 13423 41292 13491 41348
rect 13547 41292 13615 41348
rect 13671 41292 13739 41348
rect 13795 41292 13863 41348
rect 13919 41292 13987 41348
rect 14043 41292 14111 41348
rect 14167 41292 14235 41348
rect 14291 41292 14359 41348
rect 14415 41292 14483 41348
rect 14539 41292 14607 41348
rect 14663 41292 14673 41348
rect 12861 41224 14673 41292
rect 12861 41168 12871 41224
rect 12927 41168 12995 41224
rect 13051 41168 13119 41224
rect 13175 41168 13243 41224
rect 13299 41168 13367 41224
rect 13423 41168 13491 41224
rect 13547 41168 13615 41224
rect 13671 41168 13739 41224
rect 13795 41168 13863 41224
rect 13919 41168 13987 41224
rect 14043 41168 14111 41224
rect 14167 41168 14235 41224
rect 14291 41168 14359 41224
rect 14415 41168 14483 41224
rect 14539 41168 14607 41224
rect 14663 41168 14673 41224
rect 12861 41100 14673 41168
rect 12861 41044 12871 41100
rect 12927 41044 12995 41100
rect 13051 41044 13119 41100
rect 13175 41044 13243 41100
rect 13299 41044 13367 41100
rect 13423 41044 13491 41100
rect 13547 41044 13615 41100
rect 13671 41044 13739 41100
rect 13795 41044 13863 41100
rect 13919 41044 13987 41100
rect 14043 41044 14111 41100
rect 14167 41044 14235 41100
rect 14291 41044 14359 41100
rect 14415 41044 14483 41100
rect 14539 41044 14607 41100
rect 14663 41044 14673 41100
rect 12861 40976 14673 41044
rect 12861 40920 12871 40976
rect 12927 40920 12995 40976
rect 13051 40920 13119 40976
rect 13175 40920 13243 40976
rect 13299 40920 13367 40976
rect 13423 40920 13491 40976
rect 13547 40920 13615 40976
rect 13671 40920 13739 40976
rect 13795 40920 13863 40976
rect 13919 40920 13987 40976
rect 14043 40920 14111 40976
rect 14167 40920 14235 40976
rect 14291 40920 14359 40976
rect 14415 40920 14483 40976
rect 14539 40920 14607 40976
rect 14663 40920 14673 40976
rect 12861 40852 14673 40920
rect 12861 40796 12871 40852
rect 12927 40796 12995 40852
rect 13051 40796 13119 40852
rect 13175 40796 13243 40852
rect 13299 40796 13367 40852
rect 13423 40796 13491 40852
rect 13547 40796 13615 40852
rect 13671 40796 13739 40852
rect 13795 40796 13863 40852
rect 13919 40796 13987 40852
rect 14043 40796 14111 40852
rect 14167 40796 14235 40852
rect 14291 40796 14359 40852
rect 14415 40796 14483 40852
rect 14539 40796 14607 40852
rect 14663 40796 14673 40852
rect 12861 40728 14673 40796
rect 12861 40672 12871 40728
rect 12927 40672 12995 40728
rect 13051 40672 13119 40728
rect 13175 40672 13243 40728
rect 13299 40672 13367 40728
rect 13423 40672 13491 40728
rect 13547 40672 13615 40728
rect 13671 40672 13739 40728
rect 13795 40672 13863 40728
rect 13919 40672 13987 40728
rect 14043 40672 14111 40728
rect 14167 40672 14235 40728
rect 14291 40672 14359 40728
rect 14415 40672 14483 40728
rect 14539 40672 14607 40728
rect 14663 40672 14673 40728
rect 12861 40604 14673 40672
rect 12861 40548 12871 40604
rect 12927 40548 12995 40604
rect 13051 40548 13119 40604
rect 13175 40548 13243 40604
rect 13299 40548 13367 40604
rect 13423 40548 13491 40604
rect 13547 40548 13615 40604
rect 13671 40548 13739 40604
rect 13795 40548 13863 40604
rect 13919 40548 13987 40604
rect 14043 40548 14111 40604
rect 14167 40548 14235 40604
rect 14291 40548 14359 40604
rect 14415 40548 14483 40604
rect 14539 40548 14607 40604
rect 14663 40548 14673 40604
rect 12861 40480 14673 40548
rect 12861 40424 12871 40480
rect 12927 40424 12995 40480
rect 13051 40424 13119 40480
rect 13175 40424 13243 40480
rect 13299 40424 13367 40480
rect 13423 40424 13491 40480
rect 13547 40424 13615 40480
rect 13671 40424 13739 40480
rect 13795 40424 13863 40480
rect 13919 40424 13987 40480
rect 14043 40424 14111 40480
rect 14167 40424 14235 40480
rect 14291 40424 14359 40480
rect 14415 40424 14483 40480
rect 14539 40424 14607 40480
rect 14663 40424 14673 40480
rect 12861 40356 14673 40424
rect 12861 40300 12871 40356
rect 12927 40300 12995 40356
rect 13051 40300 13119 40356
rect 13175 40300 13243 40356
rect 13299 40300 13367 40356
rect 13423 40300 13491 40356
rect 13547 40300 13615 40356
rect 13671 40300 13739 40356
rect 13795 40300 13863 40356
rect 13919 40300 13987 40356
rect 14043 40300 14111 40356
rect 14167 40300 14235 40356
rect 14291 40300 14359 40356
rect 14415 40300 14483 40356
rect 14539 40300 14607 40356
rect 14663 40300 14673 40356
rect 12861 40232 14673 40300
rect 12861 40176 12871 40232
rect 12927 40176 12995 40232
rect 13051 40176 13119 40232
rect 13175 40176 13243 40232
rect 13299 40176 13367 40232
rect 13423 40176 13491 40232
rect 13547 40176 13615 40232
rect 13671 40176 13739 40232
rect 13795 40176 13863 40232
rect 13919 40176 13987 40232
rect 14043 40176 14111 40232
rect 14167 40176 14235 40232
rect 14291 40176 14359 40232
rect 14415 40176 14483 40232
rect 14539 40176 14607 40232
rect 14663 40176 14673 40232
rect 12861 40108 14673 40176
rect 12861 40052 12871 40108
rect 12927 40052 12995 40108
rect 13051 40052 13119 40108
rect 13175 40052 13243 40108
rect 13299 40052 13367 40108
rect 13423 40052 13491 40108
rect 13547 40052 13615 40108
rect 13671 40052 13739 40108
rect 13795 40052 13863 40108
rect 13919 40052 13987 40108
rect 14043 40052 14111 40108
rect 14167 40052 14235 40108
rect 14291 40052 14359 40108
rect 14415 40052 14483 40108
rect 14539 40052 14607 40108
rect 14663 40052 14673 40108
rect 12861 40042 14673 40052
rect 305 39748 2117 39758
rect 305 39692 315 39748
rect 371 39692 439 39748
rect 495 39692 563 39748
rect 619 39692 687 39748
rect 743 39692 811 39748
rect 867 39692 935 39748
rect 991 39692 1059 39748
rect 1115 39692 1183 39748
rect 1239 39692 1307 39748
rect 1363 39692 1431 39748
rect 1487 39692 1555 39748
rect 1611 39692 1679 39748
rect 1735 39692 1803 39748
rect 1859 39692 1927 39748
rect 1983 39692 2051 39748
rect 2107 39692 2117 39748
rect 305 39624 2117 39692
rect 305 39568 315 39624
rect 371 39568 439 39624
rect 495 39568 563 39624
rect 619 39568 687 39624
rect 743 39568 811 39624
rect 867 39568 935 39624
rect 991 39568 1059 39624
rect 1115 39568 1183 39624
rect 1239 39568 1307 39624
rect 1363 39568 1431 39624
rect 1487 39568 1555 39624
rect 1611 39568 1679 39624
rect 1735 39568 1803 39624
rect 1859 39568 1927 39624
rect 1983 39568 2051 39624
rect 2107 39568 2117 39624
rect 305 39500 2117 39568
rect 305 39444 315 39500
rect 371 39444 439 39500
rect 495 39444 563 39500
rect 619 39444 687 39500
rect 743 39444 811 39500
rect 867 39444 935 39500
rect 991 39444 1059 39500
rect 1115 39444 1183 39500
rect 1239 39444 1307 39500
rect 1363 39444 1431 39500
rect 1487 39444 1555 39500
rect 1611 39444 1679 39500
rect 1735 39444 1803 39500
rect 1859 39444 1927 39500
rect 1983 39444 2051 39500
rect 2107 39444 2117 39500
rect 305 39376 2117 39444
rect 305 39320 315 39376
rect 371 39320 439 39376
rect 495 39320 563 39376
rect 619 39320 687 39376
rect 743 39320 811 39376
rect 867 39320 935 39376
rect 991 39320 1059 39376
rect 1115 39320 1183 39376
rect 1239 39320 1307 39376
rect 1363 39320 1431 39376
rect 1487 39320 1555 39376
rect 1611 39320 1679 39376
rect 1735 39320 1803 39376
rect 1859 39320 1927 39376
rect 1983 39320 2051 39376
rect 2107 39320 2117 39376
rect 305 39252 2117 39320
rect 305 39196 315 39252
rect 371 39196 439 39252
rect 495 39196 563 39252
rect 619 39196 687 39252
rect 743 39196 811 39252
rect 867 39196 935 39252
rect 991 39196 1059 39252
rect 1115 39196 1183 39252
rect 1239 39196 1307 39252
rect 1363 39196 1431 39252
rect 1487 39196 1555 39252
rect 1611 39196 1679 39252
rect 1735 39196 1803 39252
rect 1859 39196 1927 39252
rect 1983 39196 2051 39252
rect 2107 39196 2117 39252
rect 305 39128 2117 39196
rect 305 39072 315 39128
rect 371 39072 439 39128
rect 495 39072 563 39128
rect 619 39072 687 39128
rect 743 39072 811 39128
rect 867 39072 935 39128
rect 991 39072 1059 39128
rect 1115 39072 1183 39128
rect 1239 39072 1307 39128
rect 1363 39072 1431 39128
rect 1487 39072 1555 39128
rect 1611 39072 1679 39128
rect 1735 39072 1803 39128
rect 1859 39072 1927 39128
rect 1983 39072 2051 39128
rect 2107 39072 2117 39128
rect 305 39004 2117 39072
rect 305 38948 315 39004
rect 371 38948 439 39004
rect 495 38948 563 39004
rect 619 38948 687 39004
rect 743 38948 811 39004
rect 867 38948 935 39004
rect 991 38948 1059 39004
rect 1115 38948 1183 39004
rect 1239 38948 1307 39004
rect 1363 38948 1431 39004
rect 1487 38948 1555 39004
rect 1611 38948 1679 39004
rect 1735 38948 1803 39004
rect 1859 38948 1927 39004
rect 1983 38948 2051 39004
rect 2107 38948 2117 39004
rect 305 38880 2117 38948
rect 305 38824 315 38880
rect 371 38824 439 38880
rect 495 38824 563 38880
rect 619 38824 687 38880
rect 743 38824 811 38880
rect 867 38824 935 38880
rect 991 38824 1059 38880
rect 1115 38824 1183 38880
rect 1239 38824 1307 38880
rect 1363 38824 1431 38880
rect 1487 38824 1555 38880
rect 1611 38824 1679 38880
rect 1735 38824 1803 38880
rect 1859 38824 1927 38880
rect 1983 38824 2051 38880
rect 2107 38824 2117 38880
rect 305 38756 2117 38824
rect 305 38700 315 38756
rect 371 38700 439 38756
rect 495 38700 563 38756
rect 619 38700 687 38756
rect 743 38700 811 38756
rect 867 38700 935 38756
rect 991 38700 1059 38756
rect 1115 38700 1183 38756
rect 1239 38700 1307 38756
rect 1363 38700 1431 38756
rect 1487 38700 1555 38756
rect 1611 38700 1679 38756
rect 1735 38700 1803 38756
rect 1859 38700 1927 38756
rect 1983 38700 2051 38756
rect 2107 38700 2117 38756
rect 305 38632 2117 38700
rect 305 38576 315 38632
rect 371 38576 439 38632
rect 495 38576 563 38632
rect 619 38576 687 38632
rect 743 38576 811 38632
rect 867 38576 935 38632
rect 991 38576 1059 38632
rect 1115 38576 1183 38632
rect 1239 38576 1307 38632
rect 1363 38576 1431 38632
rect 1487 38576 1555 38632
rect 1611 38576 1679 38632
rect 1735 38576 1803 38632
rect 1859 38576 1927 38632
rect 1983 38576 2051 38632
rect 2107 38576 2117 38632
rect 305 38508 2117 38576
rect 305 38452 315 38508
rect 371 38452 439 38508
rect 495 38452 563 38508
rect 619 38452 687 38508
rect 743 38452 811 38508
rect 867 38452 935 38508
rect 991 38452 1059 38508
rect 1115 38452 1183 38508
rect 1239 38452 1307 38508
rect 1363 38452 1431 38508
rect 1487 38452 1555 38508
rect 1611 38452 1679 38508
rect 1735 38452 1803 38508
rect 1859 38452 1927 38508
rect 1983 38452 2051 38508
rect 2107 38452 2117 38508
rect 305 38442 2117 38452
rect 2798 39748 4734 39758
rect 2798 39692 2808 39748
rect 2864 39692 2932 39748
rect 2988 39692 3056 39748
rect 3112 39692 3180 39748
rect 3236 39692 3304 39748
rect 3360 39692 3428 39748
rect 3484 39692 3552 39748
rect 3608 39692 3676 39748
rect 3732 39692 3800 39748
rect 3856 39692 3924 39748
rect 3980 39692 4048 39748
rect 4104 39692 4172 39748
rect 4228 39692 4296 39748
rect 4352 39692 4420 39748
rect 4476 39692 4544 39748
rect 4600 39692 4668 39748
rect 4724 39692 4734 39748
rect 2798 39624 4734 39692
rect 2798 39568 2808 39624
rect 2864 39568 2932 39624
rect 2988 39568 3056 39624
rect 3112 39568 3180 39624
rect 3236 39568 3304 39624
rect 3360 39568 3428 39624
rect 3484 39568 3552 39624
rect 3608 39568 3676 39624
rect 3732 39568 3800 39624
rect 3856 39568 3924 39624
rect 3980 39568 4048 39624
rect 4104 39568 4172 39624
rect 4228 39568 4296 39624
rect 4352 39568 4420 39624
rect 4476 39568 4544 39624
rect 4600 39568 4668 39624
rect 4724 39568 4734 39624
rect 2798 39500 4734 39568
rect 2798 39444 2808 39500
rect 2864 39444 2932 39500
rect 2988 39444 3056 39500
rect 3112 39444 3180 39500
rect 3236 39444 3304 39500
rect 3360 39444 3428 39500
rect 3484 39444 3552 39500
rect 3608 39444 3676 39500
rect 3732 39444 3800 39500
rect 3856 39444 3924 39500
rect 3980 39444 4048 39500
rect 4104 39444 4172 39500
rect 4228 39444 4296 39500
rect 4352 39444 4420 39500
rect 4476 39444 4544 39500
rect 4600 39444 4668 39500
rect 4724 39444 4734 39500
rect 2798 39376 4734 39444
rect 2798 39320 2808 39376
rect 2864 39320 2932 39376
rect 2988 39320 3056 39376
rect 3112 39320 3180 39376
rect 3236 39320 3304 39376
rect 3360 39320 3428 39376
rect 3484 39320 3552 39376
rect 3608 39320 3676 39376
rect 3732 39320 3800 39376
rect 3856 39320 3924 39376
rect 3980 39320 4048 39376
rect 4104 39320 4172 39376
rect 4228 39320 4296 39376
rect 4352 39320 4420 39376
rect 4476 39320 4544 39376
rect 4600 39320 4668 39376
rect 4724 39320 4734 39376
rect 2798 39252 4734 39320
rect 2798 39196 2808 39252
rect 2864 39196 2932 39252
rect 2988 39196 3056 39252
rect 3112 39196 3180 39252
rect 3236 39196 3304 39252
rect 3360 39196 3428 39252
rect 3484 39196 3552 39252
rect 3608 39196 3676 39252
rect 3732 39196 3800 39252
rect 3856 39196 3924 39252
rect 3980 39196 4048 39252
rect 4104 39196 4172 39252
rect 4228 39196 4296 39252
rect 4352 39196 4420 39252
rect 4476 39196 4544 39252
rect 4600 39196 4668 39252
rect 4724 39196 4734 39252
rect 2798 39128 4734 39196
rect 2798 39072 2808 39128
rect 2864 39072 2932 39128
rect 2988 39072 3056 39128
rect 3112 39072 3180 39128
rect 3236 39072 3304 39128
rect 3360 39072 3428 39128
rect 3484 39072 3552 39128
rect 3608 39072 3676 39128
rect 3732 39072 3800 39128
rect 3856 39072 3924 39128
rect 3980 39072 4048 39128
rect 4104 39072 4172 39128
rect 4228 39072 4296 39128
rect 4352 39072 4420 39128
rect 4476 39072 4544 39128
rect 4600 39072 4668 39128
rect 4724 39072 4734 39128
rect 2798 39004 4734 39072
rect 2798 38948 2808 39004
rect 2864 38948 2932 39004
rect 2988 38948 3056 39004
rect 3112 38948 3180 39004
rect 3236 38948 3304 39004
rect 3360 38948 3428 39004
rect 3484 38948 3552 39004
rect 3608 38948 3676 39004
rect 3732 38948 3800 39004
rect 3856 38948 3924 39004
rect 3980 38948 4048 39004
rect 4104 38948 4172 39004
rect 4228 38948 4296 39004
rect 4352 38948 4420 39004
rect 4476 38948 4544 39004
rect 4600 38948 4668 39004
rect 4724 38948 4734 39004
rect 2798 38880 4734 38948
rect 2798 38824 2808 38880
rect 2864 38824 2932 38880
rect 2988 38824 3056 38880
rect 3112 38824 3180 38880
rect 3236 38824 3304 38880
rect 3360 38824 3428 38880
rect 3484 38824 3552 38880
rect 3608 38824 3676 38880
rect 3732 38824 3800 38880
rect 3856 38824 3924 38880
rect 3980 38824 4048 38880
rect 4104 38824 4172 38880
rect 4228 38824 4296 38880
rect 4352 38824 4420 38880
rect 4476 38824 4544 38880
rect 4600 38824 4668 38880
rect 4724 38824 4734 38880
rect 2798 38756 4734 38824
rect 2798 38700 2808 38756
rect 2864 38700 2932 38756
rect 2988 38700 3056 38756
rect 3112 38700 3180 38756
rect 3236 38700 3304 38756
rect 3360 38700 3428 38756
rect 3484 38700 3552 38756
rect 3608 38700 3676 38756
rect 3732 38700 3800 38756
rect 3856 38700 3924 38756
rect 3980 38700 4048 38756
rect 4104 38700 4172 38756
rect 4228 38700 4296 38756
rect 4352 38700 4420 38756
rect 4476 38700 4544 38756
rect 4600 38700 4668 38756
rect 4724 38700 4734 38756
rect 2798 38632 4734 38700
rect 2798 38576 2808 38632
rect 2864 38576 2932 38632
rect 2988 38576 3056 38632
rect 3112 38576 3180 38632
rect 3236 38576 3304 38632
rect 3360 38576 3428 38632
rect 3484 38576 3552 38632
rect 3608 38576 3676 38632
rect 3732 38576 3800 38632
rect 3856 38576 3924 38632
rect 3980 38576 4048 38632
rect 4104 38576 4172 38632
rect 4228 38576 4296 38632
rect 4352 38576 4420 38632
rect 4476 38576 4544 38632
rect 4600 38576 4668 38632
rect 4724 38576 4734 38632
rect 2798 38508 4734 38576
rect 2798 38452 2808 38508
rect 2864 38452 2932 38508
rect 2988 38452 3056 38508
rect 3112 38452 3180 38508
rect 3236 38452 3304 38508
rect 3360 38452 3428 38508
rect 3484 38452 3552 38508
rect 3608 38452 3676 38508
rect 3732 38452 3800 38508
rect 3856 38452 3924 38508
rect 3980 38452 4048 38508
rect 4104 38452 4172 38508
rect 4228 38452 4296 38508
rect 4352 38452 4420 38508
rect 4476 38452 4544 38508
rect 4600 38452 4668 38508
rect 4724 38452 4734 38508
rect 2798 38442 4734 38452
rect 5168 39748 7104 39758
rect 5168 39692 5178 39748
rect 5234 39692 5302 39748
rect 5358 39692 5426 39748
rect 5482 39692 5550 39748
rect 5606 39692 5674 39748
rect 5730 39692 5798 39748
rect 5854 39692 5922 39748
rect 5978 39692 6046 39748
rect 6102 39692 6170 39748
rect 6226 39692 6294 39748
rect 6350 39692 6418 39748
rect 6474 39692 6542 39748
rect 6598 39692 6666 39748
rect 6722 39692 6790 39748
rect 6846 39692 6914 39748
rect 6970 39692 7038 39748
rect 7094 39692 7104 39748
rect 5168 39624 7104 39692
rect 5168 39568 5178 39624
rect 5234 39568 5302 39624
rect 5358 39568 5426 39624
rect 5482 39568 5550 39624
rect 5606 39568 5674 39624
rect 5730 39568 5798 39624
rect 5854 39568 5922 39624
rect 5978 39568 6046 39624
rect 6102 39568 6170 39624
rect 6226 39568 6294 39624
rect 6350 39568 6418 39624
rect 6474 39568 6542 39624
rect 6598 39568 6666 39624
rect 6722 39568 6790 39624
rect 6846 39568 6914 39624
rect 6970 39568 7038 39624
rect 7094 39568 7104 39624
rect 5168 39500 7104 39568
rect 5168 39444 5178 39500
rect 5234 39444 5302 39500
rect 5358 39444 5426 39500
rect 5482 39444 5550 39500
rect 5606 39444 5674 39500
rect 5730 39444 5798 39500
rect 5854 39444 5922 39500
rect 5978 39444 6046 39500
rect 6102 39444 6170 39500
rect 6226 39444 6294 39500
rect 6350 39444 6418 39500
rect 6474 39444 6542 39500
rect 6598 39444 6666 39500
rect 6722 39444 6790 39500
rect 6846 39444 6914 39500
rect 6970 39444 7038 39500
rect 7094 39444 7104 39500
rect 5168 39376 7104 39444
rect 5168 39320 5178 39376
rect 5234 39320 5302 39376
rect 5358 39320 5426 39376
rect 5482 39320 5550 39376
rect 5606 39320 5674 39376
rect 5730 39320 5798 39376
rect 5854 39320 5922 39376
rect 5978 39320 6046 39376
rect 6102 39320 6170 39376
rect 6226 39320 6294 39376
rect 6350 39320 6418 39376
rect 6474 39320 6542 39376
rect 6598 39320 6666 39376
rect 6722 39320 6790 39376
rect 6846 39320 6914 39376
rect 6970 39320 7038 39376
rect 7094 39320 7104 39376
rect 5168 39252 7104 39320
rect 5168 39196 5178 39252
rect 5234 39196 5302 39252
rect 5358 39196 5426 39252
rect 5482 39196 5550 39252
rect 5606 39196 5674 39252
rect 5730 39196 5798 39252
rect 5854 39196 5922 39252
rect 5978 39196 6046 39252
rect 6102 39196 6170 39252
rect 6226 39196 6294 39252
rect 6350 39196 6418 39252
rect 6474 39196 6542 39252
rect 6598 39196 6666 39252
rect 6722 39196 6790 39252
rect 6846 39196 6914 39252
rect 6970 39196 7038 39252
rect 7094 39196 7104 39252
rect 5168 39128 7104 39196
rect 5168 39072 5178 39128
rect 5234 39072 5302 39128
rect 5358 39072 5426 39128
rect 5482 39072 5550 39128
rect 5606 39072 5674 39128
rect 5730 39072 5798 39128
rect 5854 39072 5922 39128
rect 5978 39072 6046 39128
rect 6102 39072 6170 39128
rect 6226 39072 6294 39128
rect 6350 39072 6418 39128
rect 6474 39072 6542 39128
rect 6598 39072 6666 39128
rect 6722 39072 6790 39128
rect 6846 39072 6914 39128
rect 6970 39072 7038 39128
rect 7094 39072 7104 39128
rect 5168 39004 7104 39072
rect 5168 38948 5178 39004
rect 5234 38948 5302 39004
rect 5358 38948 5426 39004
rect 5482 38948 5550 39004
rect 5606 38948 5674 39004
rect 5730 38948 5798 39004
rect 5854 38948 5922 39004
rect 5978 38948 6046 39004
rect 6102 38948 6170 39004
rect 6226 38948 6294 39004
rect 6350 38948 6418 39004
rect 6474 38948 6542 39004
rect 6598 38948 6666 39004
rect 6722 38948 6790 39004
rect 6846 38948 6914 39004
rect 6970 38948 7038 39004
rect 7094 38948 7104 39004
rect 5168 38880 7104 38948
rect 5168 38824 5178 38880
rect 5234 38824 5302 38880
rect 5358 38824 5426 38880
rect 5482 38824 5550 38880
rect 5606 38824 5674 38880
rect 5730 38824 5798 38880
rect 5854 38824 5922 38880
rect 5978 38824 6046 38880
rect 6102 38824 6170 38880
rect 6226 38824 6294 38880
rect 6350 38824 6418 38880
rect 6474 38824 6542 38880
rect 6598 38824 6666 38880
rect 6722 38824 6790 38880
rect 6846 38824 6914 38880
rect 6970 38824 7038 38880
rect 7094 38824 7104 38880
rect 5168 38756 7104 38824
rect 5168 38700 5178 38756
rect 5234 38700 5302 38756
rect 5358 38700 5426 38756
rect 5482 38700 5550 38756
rect 5606 38700 5674 38756
rect 5730 38700 5798 38756
rect 5854 38700 5922 38756
rect 5978 38700 6046 38756
rect 6102 38700 6170 38756
rect 6226 38700 6294 38756
rect 6350 38700 6418 38756
rect 6474 38700 6542 38756
rect 6598 38700 6666 38756
rect 6722 38700 6790 38756
rect 6846 38700 6914 38756
rect 6970 38700 7038 38756
rect 7094 38700 7104 38756
rect 5168 38632 7104 38700
rect 5168 38576 5178 38632
rect 5234 38576 5302 38632
rect 5358 38576 5426 38632
rect 5482 38576 5550 38632
rect 5606 38576 5674 38632
rect 5730 38576 5798 38632
rect 5854 38576 5922 38632
rect 5978 38576 6046 38632
rect 6102 38576 6170 38632
rect 6226 38576 6294 38632
rect 6350 38576 6418 38632
rect 6474 38576 6542 38632
rect 6598 38576 6666 38632
rect 6722 38576 6790 38632
rect 6846 38576 6914 38632
rect 6970 38576 7038 38632
rect 7094 38576 7104 38632
rect 5168 38508 7104 38576
rect 5168 38452 5178 38508
rect 5234 38452 5302 38508
rect 5358 38452 5426 38508
rect 5482 38452 5550 38508
rect 5606 38452 5674 38508
rect 5730 38452 5798 38508
rect 5854 38452 5922 38508
rect 5978 38452 6046 38508
rect 6102 38452 6170 38508
rect 6226 38452 6294 38508
rect 6350 38452 6418 38508
rect 6474 38452 6542 38508
rect 6598 38452 6666 38508
rect 6722 38452 6790 38508
rect 6846 38452 6914 38508
rect 6970 38452 7038 38508
rect 7094 38452 7104 38508
rect 5168 38442 7104 38452
rect 7874 39748 9810 39758
rect 7874 39692 7884 39748
rect 7940 39692 8008 39748
rect 8064 39692 8132 39748
rect 8188 39692 8256 39748
rect 8312 39692 8380 39748
rect 8436 39692 8504 39748
rect 8560 39692 8628 39748
rect 8684 39692 8752 39748
rect 8808 39692 8876 39748
rect 8932 39692 9000 39748
rect 9056 39692 9124 39748
rect 9180 39692 9248 39748
rect 9304 39692 9372 39748
rect 9428 39692 9496 39748
rect 9552 39692 9620 39748
rect 9676 39692 9744 39748
rect 9800 39692 9810 39748
rect 7874 39624 9810 39692
rect 7874 39568 7884 39624
rect 7940 39568 8008 39624
rect 8064 39568 8132 39624
rect 8188 39568 8256 39624
rect 8312 39568 8380 39624
rect 8436 39568 8504 39624
rect 8560 39568 8628 39624
rect 8684 39568 8752 39624
rect 8808 39568 8876 39624
rect 8932 39568 9000 39624
rect 9056 39568 9124 39624
rect 9180 39568 9248 39624
rect 9304 39568 9372 39624
rect 9428 39568 9496 39624
rect 9552 39568 9620 39624
rect 9676 39568 9744 39624
rect 9800 39568 9810 39624
rect 7874 39500 9810 39568
rect 7874 39444 7884 39500
rect 7940 39444 8008 39500
rect 8064 39444 8132 39500
rect 8188 39444 8256 39500
rect 8312 39444 8380 39500
rect 8436 39444 8504 39500
rect 8560 39444 8628 39500
rect 8684 39444 8752 39500
rect 8808 39444 8876 39500
rect 8932 39444 9000 39500
rect 9056 39444 9124 39500
rect 9180 39444 9248 39500
rect 9304 39444 9372 39500
rect 9428 39444 9496 39500
rect 9552 39444 9620 39500
rect 9676 39444 9744 39500
rect 9800 39444 9810 39500
rect 7874 39376 9810 39444
rect 7874 39320 7884 39376
rect 7940 39320 8008 39376
rect 8064 39320 8132 39376
rect 8188 39320 8256 39376
rect 8312 39320 8380 39376
rect 8436 39320 8504 39376
rect 8560 39320 8628 39376
rect 8684 39320 8752 39376
rect 8808 39320 8876 39376
rect 8932 39320 9000 39376
rect 9056 39320 9124 39376
rect 9180 39320 9248 39376
rect 9304 39320 9372 39376
rect 9428 39320 9496 39376
rect 9552 39320 9620 39376
rect 9676 39320 9744 39376
rect 9800 39320 9810 39376
rect 7874 39252 9810 39320
rect 7874 39196 7884 39252
rect 7940 39196 8008 39252
rect 8064 39196 8132 39252
rect 8188 39196 8256 39252
rect 8312 39196 8380 39252
rect 8436 39196 8504 39252
rect 8560 39196 8628 39252
rect 8684 39196 8752 39252
rect 8808 39196 8876 39252
rect 8932 39196 9000 39252
rect 9056 39196 9124 39252
rect 9180 39196 9248 39252
rect 9304 39196 9372 39252
rect 9428 39196 9496 39252
rect 9552 39196 9620 39252
rect 9676 39196 9744 39252
rect 9800 39196 9810 39252
rect 7874 39128 9810 39196
rect 7874 39072 7884 39128
rect 7940 39072 8008 39128
rect 8064 39072 8132 39128
rect 8188 39072 8256 39128
rect 8312 39072 8380 39128
rect 8436 39072 8504 39128
rect 8560 39072 8628 39128
rect 8684 39072 8752 39128
rect 8808 39072 8876 39128
rect 8932 39072 9000 39128
rect 9056 39072 9124 39128
rect 9180 39072 9248 39128
rect 9304 39072 9372 39128
rect 9428 39072 9496 39128
rect 9552 39072 9620 39128
rect 9676 39072 9744 39128
rect 9800 39072 9810 39128
rect 7874 39004 9810 39072
rect 7874 38948 7884 39004
rect 7940 38948 8008 39004
rect 8064 38948 8132 39004
rect 8188 38948 8256 39004
rect 8312 38948 8380 39004
rect 8436 38948 8504 39004
rect 8560 38948 8628 39004
rect 8684 38948 8752 39004
rect 8808 38948 8876 39004
rect 8932 38948 9000 39004
rect 9056 38948 9124 39004
rect 9180 38948 9248 39004
rect 9304 38948 9372 39004
rect 9428 38948 9496 39004
rect 9552 38948 9620 39004
rect 9676 38948 9744 39004
rect 9800 38948 9810 39004
rect 7874 38880 9810 38948
rect 7874 38824 7884 38880
rect 7940 38824 8008 38880
rect 8064 38824 8132 38880
rect 8188 38824 8256 38880
rect 8312 38824 8380 38880
rect 8436 38824 8504 38880
rect 8560 38824 8628 38880
rect 8684 38824 8752 38880
rect 8808 38824 8876 38880
rect 8932 38824 9000 38880
rect 9056 38824 9124 38880
rect 9180 38824 9248 38880
rect 9304 38824 9372 38880
rect 9428 38824 9496 38880
rect 9552 38824 9620 38880
rect 9676 38824 9744 38880
rect 9800 38824 9810 38880
rect 7874 38756 9810 38824
rect 7874 38700 7884 38756
rect 7940 38700 8008 38756
rect 8064 38700 8132 38756
rect 8188 38700 8256 38756
rect 8312 38700 8380 38756
rect 8436 38700 8504 38756
rect 8560 38700 8628 38756
rect 8684 38700 8752 38756
rect 8808 38700 8876 38756
rect 8932 38700 9000 38756
rect 9056 38700 9124 38756
rect 9180 38700 9248 38756
rect 9304 38700 9372 38756
rect 9428 38700 9496 38756
rect 9552 38700 9620 38756
rect 9676 38700 9744 38756
rect 9800 38700 9810 38756
rect 7874 38632 9810 38700
rect 7874 38576 7884 38632
rect 7940 38576 8008 38632
rect 8064 38576 8132 38632
rect 8188 38576 8256 38632
rect 8312 38576 8380 38632
rect 8436 38576 8504 38632
rect 8560 38576 8628 38632
rect 8684 38576 8752 38632
rect 8808 38576 8876 38632
rect 8932 38576 9000 38632
rect 9056 38576 9124 38632
rect 9180 38576 9248 38632
rect 9304 38576 9372 38632
rect 9428 38576 9496 38632
rect 9552 38576 9620 38632
rect 9676 38576 9744 38632
rect 9800 38576 9810 38632
rect 7874 38508 9810 38576
rect 7874 38452 7884 38508
rect 7940 38452 8008 38508
rect 8064 38452 8132 38508
rect 8188 38452 8256 38508
rect 8312 38452 8380 38508
rect 8436 38452 8504 38508
rect 8560 38452 8628 38508
rect 8684 38452 8752 38508
rect 8808 38452 8876 38508
rect 8932 38452 9000 38508
rect 9056 38452 9124 38508
rect 9180 38452 9248 38508
rect 9304 38452 9372 38508
rect 9428 38452 9496 38508
rect 9552 38452 9620 38508
rect 9676 38452 9744 38508
rect 9800 38452 9810 38508
rect 7874 38442 9810 38452
rect 10244 39748 12180 39758
rect 10244 39692 10254 39748
rect 10310 39692 10378 39748
rect 10434 39692 10502 39748
rect 10558 39692 10626 39748
rect 10682 39692 10750 39748
rect 10806 39692 10874 39748
rect 10930 39692 10998 39748
rect 11054 39692 11122 39748
rect 11178 39692 11246 39748
rect 11302 39692 11370 39748
rect 11426 39692 11494 39748
rect 11550 39692 11618 39748
rect 11674 39692 11742 39748
rect 11798 39692 11866 39748
rect 11922 39692 11990 39748
rect 12046 39692 12114 39748
rect 12170 39692 12180 39748
rect 10244 39624 12180 39692
rect 10244 39568 10254 39624
rect 10310 39568 10378 39624
rect 10434 39568 10502 39624
rect 10558 39568 10626 39624
rect 10682 39568 10750 39624
rect 10806 39568 10874 39624
rect 10930 39568 10998 39624
rect 11054 39568 11122 39624
rect 11178 39568 11246 39624
rect 11302 39568 11370 39624
rect 11426 39568 11494 39624
rect 11550 39568 11618 39624
rect 11674 39568 11742 39624
rect 11798 39568 11866 39624
rect 11922 39568 11990 39624
rect 12046 39568 12114 39624
rect 12170 39568 12180 39624
rect 10244 39500 12180 39568
rect 10244 39444 10254 39500
rect 10310 39444 10378 39500
rect 10434 39444 10502 39500
rect 10558 39444 10626 39500
rect 10682 39444 10750 39500
rect 10806 39444 10874 39500
rect 10930 39444 10998 39500
rect 11054 39444 11122 39500
rect 11178 39444 11246 39500
rect 11302 39444 11370 39500
rect 11426 39444 11494 39500
rect 11550 39444 11618 39500
rect 11674 39444 11742 39500
rect 11798 39444 11866 39500
rect 11922 39444 11990 39500
rect 12046 39444 12114 39500
rect 12170 39444 12180 39500
rect 10244 39376 12180 39444
rect 10244 39320 10254 39376
rect 10310 39320 10378 39376
rect 10434 39320 10502 39376
rect 10558 39320 10626 39376
rect 10682 39320 10750 39376
rect 10806 39320 10874 39376
rect 10930 39320 10998 39376
rect 11054 39320 11122 39376
rect 11178 39320 11246 39376
rect 11302 39320 11370 39376
rect 11426 39320 11494 39376
rect 11550 39320 11618 39376
rect 11674 39320 11742 39376
rect 11798 39320 11866 39376
rect 11922 39320 11990 39376
rect 12046 39320 12114 39376
rect 12170 39320 12180 39376
rect 10244 39252 12180 39320
rect 10244 39196 10254 39252
rect 10310 39196 10378 39252
rect 10434 39196 10502 39252
rect 10558 39196 10626 39252
rect 10682 39196 10750 39252
rect 10806 39196 10874 39252
rect 10930 39196 10998 39252
rect 11054 39196 11122 39252
rect 11178 39196 11246 39252
rect 11302 39196 11370 39252
rect 11426 39196 11494 39252
rect 11550 39196 11618 39252
rect 11674 39196 11742 39252
rect 11798 39196 11866 39252
rect 11922 39196 11990 39252
rect 12046 39196 12114 39252
rect 12170 39196 12180 39252
rect 10244 39128 12180 39196
rect 10244 39072 10254 39128
rect 10310 39072 10378 39128
rect 10434 39072 10502 39128
rect 10558 39072 10626 39128
rect 10682 39072 10750 39128
rect 10806 39072 10874 39128
rect 10930 39072 10998 39128
rect 11054 39072 11122 39128
rect 11178 39072 11246 39128
rect 11302 39072 11370 39128
rect 11426 39072 11494 39128
rect 11550 39072 11618 39128
rect 11674 39072 11742 39128
rect 11798 39072 11866 39128
rect 11922 39072 11990 39128
rect 12046 39072 12114 39128
rect 12170 39072 12180 39128
rect 10244 39004 12180 39072
rect 10244 38948 10254 39004
rect 10310 38948 10378 39004
rect 10434 38948 10502 39004
rect 10558 38948 10626 39004
rect 10682 38948 10750 39004
rect 10806 38948 10874 39004
rect 10930 38948 10998 39004
rect 11054 38948 11122 39004
rect 11178 38948 11246 39004
rect 11302 38948 11370 39004
rect 11426 38948 11494 39004
rect 11550 38948 11618 39004
rect 11674 38948 11742 39004
rect 11798 38948 11866 39004
rect 11922 38948 11990 39004
rect 12046 38948 12114 39004
rect 12170 38948 12180 39004
rect 10244 38880 12180 38948
rect 10244 38824 10254 38880
rect 10310 38824 10378 38880
rect 10434 38824 10502 38880
rect 10558 38824 10626 38880
rect 10682 38824 10750 38880
rect 10806 38824 10874 38880
rect 10930 38824 10998 38880
rect 11054 38824 11122 38880
rect 11178 38824 11246 38880
rect 11302 38824 11370 38880
rect 11426 38824 11494 38880
rect 11550 38824 11618 38880
rect 11674 38824 11742 38880
rect 11798 38824 11866 38880
rect 11922 38824 11990 38880
rect 12046 38824 12114 38880
rect 12170 38824 12180 38880
rect 10244 38756 12180 38824
rect 10244 38700 10254 38756
rect 10310 38700 10378 38756
rect 10434 38700 10502 38756
rect 10558 38700 10626 38756
rect 10682 38700 10750 38756
rect 10806 38700 10874 38756
rect 10930 38700 10998 38756
rect 11054 38700 11122 38756
rect 11178 38700 11246 38756
rect 11302 38700 11370 38756
rect 11426 38700 11494 38756
rect 11550 38700 11618 38756
rect 11674 38700 11742 38756
rect 11798 38700 11866 38756
rect 11922 38700 11990 38756
rect 12046 38700 12114 38756
rect 12170 38700 12180 38756
rect 10244 38632 12180 38700
rect 10244 38576 10254 38632
rect 10310 38576 10378 38632
rect 10434 38576 10502 38632
rect 10558 38576 10626 38632
rect 10682 38576 10750 38632
rect 10806 38576 10874 38632
rect 10930 38576 10998 38632
rect 11054 38576 11122 38632
rect 11178 38576 11246 38632
rect 11302 38576 11370 38632
rect 11426 38576 11494 38632
rect 11550 38576 11618 38632
rect 11674 38576 11742 38632
rect 11798 38576 11866 38632
rect 11922 38576 11990 38632
rect 12046 38576 12114 38632
rect 12170 38576 12180 38632
rect 10244 38508 12180 38576
rect 10244 38452 10254 38508
rect 10310 38452 10378 38508
rect 10434 38452 10502 38508
rect 10558 38452 10626 38508
rect 10682 38452 10750 38508
rect 10806 38452 10874 38508
rect 10930 38452 10998 38508
rect 11054 38452 11122 38508
rect 11178 38452 11246 38508
rect 11302 38452 11370 38508
rect 11426 38452 11494 38508
rect 11550 38452 11618 38508
rect 11674 38452 11742 38508
rect 11798 38452 11866 38508
rect 11922 38452 11990 38508
rect 12046 38452 12114 38508
rect 12170 38452 12180 38508
rect 10244 38442 12180 38452
rect 12861 39748 14673 39758
rect 12861 39692 12871 39748
rect 12927 39692 12995 39748
rect 13051 39692 13119 39748
rect 13175 39692 13243 39748
rect 13299 39692 13367 39748
rect 13423 39692 13491 39748
rect 13547 39692 13615 39748
rect 13671 39692 13739 39748
rect 13795 39692 13863 39748
rect 13919 39692 13987 39748
rect 14043 39692 14111 39748
rect 14167 39692 14235 39748
rect 14291 39692 14359 39748
rect 14415 39692 14483 39748
rect 14539 39692 14607 39748
rect 14663 39692 14673 39748
rect 12861 39624 14673 39692
rect 12861 39568 12871 39624
rect 12927 39568 12995 39624
rect 13051 39568 13119 39624
rect 13175 39568 13243 39624
rect 13299 39568 13367 39624
rect 13423 39568 13491 39624
rect 13547 39568 13615 39624
rect 13671 39568 13739 39624
rect 13795 39568 13863 39624
rect 13919 39568 13987 39624
rect 14043 39568 14111 39624
rect 14167 39568 14235 39624
rect 14291 39568 14359 39624
rect 14415 39568 14483 39624
rect 14539 39568 14607 39624
rect 14663 39568 14673 39624
rect 12861 39500 14673 39568
rect 12861 39444 12871 39500
rect 12927 39444 12995 39500
rect 13051 39444 13119 39500
rect 13175 39444 13243 39500
rect 13299 39444 13367 39500
rect 13423 39444 13491 39500
rect 13547 39444 13615 39500
rect 13671 39444 13739 39500
rect 13795 39444 13863 39500
rect 13919 39444 13987 39500
rect 14043 39444 14111 39500
rect 14167 39444 14235 39500
rect 14291 39444 14359 39500
rect 14415 39444 14483 39500
rect 14539 39444 14607 39500
rect 14663 39444 14673 39500
rect 12861 39376 14673 39444
rect 12861 39320 12871 39376
rect 12927 39320 12995 39376
rect 13051 39320 13119 39376
rect 13175 39320 13243 39376
rect 13299 39320 13367 39376
rect 13423 39320 13491 39376
rect 13547 39320 13615 39376
rect 13671 39320 13739 39376
rect 13795 39320 13863 39376
rect 13919 39320 13987 39376
rect 14043 39320 14111 39376
rect 14167 39320 14235 39376
rect 14291 39320 14359 39376
rect 14415 39320 14483 39376
rect 14539 39320 14607 39376
rect 14663 39320 14673 39376
rect 12861 39252 14673 39320
rect 12861 39196 12871 39252
rect 12927 39196 12995 39252
rect 13051 39196 13119 39252
rect 13175 39196 13243 39252
rect 13299 39196 13367 39252
rect 13423 39196 13491 39252
rect 13547 39196 13615 39252
rect 13671 39196 13739 39252
rect 13795 39196 13863 39252
rect 13919 39196 13987 39252
rect 14043 39196 14111 39252
rect 14167 39196 14235 39252
rect 14291 39196 14359 39252
rect 14415 39196 14483 39252
rect 14539 39196 14607 39252
rect 14663 39196 14673 39252
rect 12861 39128 14673 39196
rect 12861 39072 12871 39128
rect 12927 39072 12995 39128
rect 13051 39072 13119 39128
rect 13175 39072 13243 39128
rect 13299 39072 13367 39128
rect 13423 39072 13491 39128
rect 13547 39072 13615 39128
rect 13671 39072 13739 39128
rect 13795 39072 13863 39128
rect 13919 39072 13987 39128
rect 14043 39072 14111 39128
rect 14167 39072 14235 39128
rect 14291 39072 14359 39128
rect 14415 39072 14483 39128
rect 14539 39072 14607 39128
rect 14663 39072 14673 39128
rect 12861 39004 14673 39072
rect 12861 38948 12871 39004
rect 12927 38948 12995 39004
rect 13051 38948 13119 39004
rect 13175 38948 13243 39004
rect 13299 38948 13367 39004
rect 13423 38948 13491 39004
rect 13547 38948 13615 39004
rect 13671 38948 13739 39004
rect 13795 38948 13863 39004
rect 13919 38948 13987 39004
rect 14043 38948 14111 39004
rect 14167 38948 14235 39004
rect 14291 38948 14359 39004
rect 14415 38948 14483 39004
rect 14539 38948 14607 39004
rect 14663 38948 14673 39004
rect 12861 38880 14673 38948
rect 12861 38824 12871 38880
rect 12927 38824 12995 38880
rect 13051 38824 13119 38880
rect 13175 38824 13243 38880
rect 13299 38824 13367 38880
rect 13423 38824 13491 38880
rect 13547 38824 13615 38880
rect 13671 38824 13739 38880
rect 13795 38824 13863 38880
rect 13919 38824 13987 38880
rect 14043 38824 14111 38880
rect 14167 38824 14235 38880
rect 14291 38824 14359 38880
rect 14415 38824 14483 38880
rect 14539 38824 14607 38880
rect 14663 38824 14673 38880
rect 12861 38756 14673 38824
rect 12861 38700 12871 38756
rect 12927 38700 12995 38756
rect 13051 38700 13119 38756
rect 13175 38700 13243 38756
rect 13299 38700 13367 38756
rect 13423 38700 13491 38756
rect 13547 38700 13615 38756
rect 13671 38700 13739 38756
rect 13795 38700 13863 38756
rect 13919 38700 13987 38756
rect 14043 38700 14111 38756
rect 14167 38700 14235 38756
rect 14291 38700 14359 38756
rect 14415 38700 14483 38756
rect 14539 38700 14607 38756
rect 14663 38700 14673 38756
rect 12861 38632 14673 38700
rect 12861 38576 12871 38632
rect 12927 38576 12995 38632
rect 13051 38576 13119 38632
rect 13175 38576 13243 38632
rect 13299 38576 13367 38632
rect 13423 38576 13491 38632
rect 13547 38576 13615 38632
rect 13671 38576 13739 38632
rect 13795 38576 13863 38632
rect 13919 38576 13987 38632
rect 14043 38576 14111 38632
rect 14167 38576 14235 38632
rect 14291 38576 14359 38632
rect 14415 38576 14483 38632
rect 14539 38576 14607 38632
rect 14663 38576 14673 38632
rect 12861 38508 14673 38576
rect 12861 38452 12871 38508
rect 12927 38452 12995 38508
rect 13051 38452 13119 38508
rect 13175 38452 13243 38508
rect 13299 38452 13367 38508
rect 13423 38452 13491 38508
rect 13547 38452 13615 38508
rect 13671 38452 13739 38508
rect 13795 38452 13863 38508
rect 13919 38452 13987 38508
rect 14043 38452 14111 38508
rect 14167 38452 14235 38508
rect 14291 38452 14359 38508
rect 14415 38452 14483 38508
rect 14539 38452 14607 38508
rect 14663 38452 14673 38508
rect 12861 38442 14673 38452
rect 10 38176 86 38186
rect 10 36824 20 38176
rect 76 36824 86 38176
rect 14892 38176 14968 38186
rect 2279 38135 2355 38145
rect 2279 38079 2289 38135
rect 2345 38079 2355 38135
rect 2279 38003 2355 38079
rect 2279 37947 2289 38003
rect 2345 37947 2355 38003
rect 2279 37871 2355 37947
rect 2279 37815 2289 37871
rect 2345 37815 2355 37871
rect 2279 37739 2355 37815
rect 2279 37683 2289 37739
rect 2345 37683 2355 37739
rect 2279 37607 2355 37683
rect 2279 37551 2289 37607
rect 2345 37551 2355 37607
rect 2279 37475 2355 37551
rect 2279 37419 2289 37475
rect 2345 37419 2355 37475
rect 2279 37343 2355 37419
rect 2279 37287 2289 37343
rect 2345 37287 2355 37343
rect 2279 37211 2355 37287
rect 2279 37155 2289 37211
rect 2345 37155 2355 37211
rect 2279 37079 2355 37155
rect 2279 37023 2289 37079
rect 2345 37023 2355 37079
rect 2279 36947 2355 37023
rect 2279 36891 2289 36947
rect 2345 36891 2355 36947
rect 2279 36881 2355 36891
rect 10 36814 86 36824
rect 14892 36824 14902 38176
rect 14958 36824 14968 38176
rect 14892 36814 14968 36824
rect 2481 36554 2681 36564
rect 2481 36498 2491 36554
rect 2547 36498 2615 36554
rect 2671 36498 2681 36554
rect 2481 36430 2681 36498
rect 2481 36374 2491 36430
rect 2547 36374 2615 36430
rect 2671 36374 2681 36430
rect 2481 36306 2681 36374
rect 2481 36250 2491 36306
rect 2547 36250 2615 36306
rect 2671 36250 2681 36306
rect 2481 36182 2681 36250
rect 2481 36126 2491 36182
rect 2547 36126 2615 36182
rect 2671 36126 2681 36182
rect 2481 36058 2681 36126
rect 2481 36002 2491 36058
rect 2547 36002 2615 36058
rect 2671 36002 2681 36058
rect 2481 35934 2681 36002
rect 2481 35878 2491 35934
rect 2547 35878 2615 35934
rect 2671 35878 2681 35934
rect 2481 35810 2681 35878
rect 2481 35754 2491 35810
rect 2547 35754 2615 35810
rect 2671 35754 2681 35810
rect 2481 35686 2681 35754
rect 2481 35630 2491 35686
rect 2547 35630 2615 35686
rect 2671 35630 2681 35686
rect 2481 35562 2681 35630
rect 2481 35506 2491 35562
rect 2547 35506 2615 35562
rect 2671 35506 2681 35562
rect 2481 35438 2681 35506
rect 2481 35382 2491 35438
rect 2547 35382 2615 35438
rect 2671 35382 2681 35438
rect 2481 35314 2681 35382
rect 2481 35258 2491 35314
rect 2547 35258 2615 35314
rect 2671 35258 2681 35314
rect 2481 35190 2681 35258
rect 2481 35134 2491 35190
rect 2547 35134 2615 35190
rect 2671 35134 2681 35190
rect 2481 35066 2681 35134
rect 2481 35010 2491 35066
rect 2547 35010 2615 35066
rect 2671 35010 2681 35066
rect 2481 34942 2681 35010
rect 2481 34886 2491 34942
rect 2547 34886 2615 34942
rect 2671 34886 2681 34942
rect 2481 34818 2681 34886
rect 2481 34762 2491 34818
rect 2547 34762 2615 34818
rect 2671 34762 2681 34818
rect 2481 34694 2681 34762
rect 2481 34638 2491 34694
rect 2547 34638 2615 34694
rect 2671 34638 2681 34694
rect 2481 34570 2681 34638
rect 2481 34514 2491 34570
rect 2547 34514 2615 34570
rect 2671 34514 2681 34570
rect 2481 34446 2681 34514
rect 2481 34390 2491 34446
rect 2547 34390 2615 34446
rect 2671 34390 2681 34446
rect 2481 34322 2681 34390
rect 2481 34266 2491 34322
rect 2547 34266 2615 34322
rect 2671 34266 2681 34322
rect 2481 34198 2681 34266
rect 2481 34142 2491 34198
rect 2547 34142 2615 34198
rect 2671 34142 2681 34198
rect 2481 34074 2681 34142
rect 2481 34018 2491 34074
rect 2547 34018 2615 34074
rect 2671 34018 2681 34074
rect 2481 33950 2681 34018
rect 2481 33894 2491 33950
rect 2547 33894 2615 33950
rect 2671 33894 2681 33950
rect 2481 33826 2681 33894
rect 2481 33770 2491 33826
rect 2547 33770 2615 33826
rect 2671 33770 2681 33826
rect 2481 33702 2681 33770
rect 2481 33646 2491 33702
rect 2547 33646 2615 33702
rect 2671 33646 2681 33702
rect 2481 33636 2681 33646
rect 4851 36554 5051 36564
rect 4851 36498 4861 36554
rect 4917 36498 4985 36554
rect 5041 36498 5051 36554
rect 4851 36430 5051 36498
rect 4851 36374 4861 36430
rect 4917 36374 4985 36430
rect 5041 36374 5051 36430
rect 4851 36306 5051 36374
rect 4851 36250 4861 36306
rect 4917 36250 4985 36306
rect 5041 36250 5051 36306
rect 4851 36182 5051 36250
rect 4851 36126 4861 36182
rect 4917 36126 4985 36182
rect 5041 36126 5051 36182
rect 4851 36058 5051 36126
rect 4851 36002 4861 36058
rect 4917 36002 4985 36058
rect 5041 36002 5051 36058
rect 4851 35934 5051 36002
rect 4851 35878 4861 35934
rect 4917 35878 4985 35934
rect 5041 35878 5051 35934
rect 4851 35810 5051 35878
rect 4851 35754 4861 35810
rect 4917 35754 4985 35810
rect 5041 35754 5051 35810
rect 4851 35686 5051 35754
rect 4851 35630 4861 35686
rect 4917 35630 4985 35686
rect 5041 35630 5051 35686
rect 4851 35562 5051 35630
rect 4851 35506 4861 35562
rect 4917 35506 4985 35562
rect 5041 35506 5051 35562
rect 4851 35438 5051 35506
rect 4851 35382 4861 35438
rect 4917 35382 4985 35438
rect 5041 35382 5051 35438
rect 4851 35314 5051 35382
rect 4851 35258 4861 35314
rect 4917 35258 4985 35314
rect 5041 35258 5051 35314
rect 4851 35190 5051 35258
rect 4851 35134 4861 35190
rect 4917 35134 4985 35190
rect 5041 35134 5051 35190
rect 4851 35066 5051 35134
rect 4851 35010 4861 35066
rect 4917 35010 4985 35066
rect 5041 35010 5051 35066
rect 4851 34942 5051 35010
rect 4851 34886 4861 34942
rect 4917 34886 4985 34942
rect 5041 34886 5051 34942
rect 4851 34818 5051 34886
rect 4851 34762 4861 34818
rect 4917 34762 4985 34818
rect 5041 34762 5051 34818
rect 4851 34694 5051 34762
rect 4851 34638 4861 34694
rect 4917 34638 4985 34694
rect 5041 34638 5051 34694
rect 4851 34570 5051 34638
rect 4851 34514 4861 34570
rect 4917 34514 4985 34570
rect 5041 34514 5051 34570
rect 4851 34446 5051 34514
rect 4851 34390 4861 34446
rect 4917 34390 4985 34446
rect 5041 34390 5051 34446
rect 4851 34322 5051 34390
rect 4851 34266 4861 34322
rect 4917 34266 4985 34322
rect 5041 34266 5051 34322
rect 4851 34198 5051 34266
rect 4851 34142 4861 34198
rect 4917 34142 4985 34198
rect 5041 34142 5051 34198
rect 4851 34074 5051 34142
rect 4851 34018 4861 34074
rect 4917 34018 4985 34074
rect 5041 34018 5051 34074
rect 4851 33950 5051 34018
rect 4851 33894 4861 33950
rect 4917 33894 4985 33950
rect 5041 33894 5051 33950
rect 4851 33826 5051 33894
rect 4851 33770 4861 33826
rect 4917 33770 4985 33826
rect 5041 33770 5051 33826
rect 4851 33702 5051 33770
rect 4851 33646 4861 33702
rect 4917 33646 4985 33702
rect 5041 33646 5051 33702
rect 4851 33636 5051 33646
rect 7265 36554 7713 36564
rect 7265 36498 7275 36554
rect 7331 36498 7399 36554
rect 7455 36498 7523 36554
rect 7579 36498 7647 36554
rect 7703 36498 7713 36554
rect 7265 36430 7713 36498
rect 7265 36374 7275 36430
rect 7331 36374 7399 36430
rect 7455 36374 7523 36430
rect 7579 36374 7647 36430
rect 7703 36374 7713 36430
rect 7265 36306 7713 36374
rect 7265 36250 7275 36306
rect 7331 36250 7399 36306
rect 7455 36250 7523 36306
rect 7579 36250 7647 36306
rect 7703 36250 7713 36306
rect 7265 36182 7713 36250
rect 7265 36126 7275 36182
rect 7331 36126 7399 36182
rect 7455 36126 7523 36182
rect 7579 36126 7647 36182
rect 7703 36126 7713 36182
rect 7265 36058 7713 36126
rect 7265 36002 7275 36058
rect 7331 36002 7399 36058
rect 7455 36002 7523 36058
rect 7579 36002 7647 36058
rect 7703 36002 7713 36058
rect 7265 35934 7713 36002
rect 7265 35878 7275 35934
rect 7331 35878 7399 35934
rect 7455 35878 7523 35934
rect 7579 35878 7647 35934
rect 7703 35878 7713 35934
rect 7265 35810 7713 35878
rect 7265 35754 7275 35810
rect 7331 35754 7399 35810
rect 7455 35754 7523 35810
rect 7579 35754 7647 35810
rect 7703 35754 7713 35810
rect 7265 35686 7713 35754
rect 7265 35630 7275 35686
rect 7331 35630 7399 35686
rect 7455 35630 7523 35686
rect 7579 35630 7647 35686
rect 7703 35630 7713 35686
rect 7265 35562 7713 35630
rect 7265 35506 7275 35562
rect 7331 35506 7399 35562
rect 7455 35506 7523 35562
rect 7579 35506 7647 35562
rect 7703 35506 7713 35562
rect 7265 35438 7713 35506
rect 7265 35382 7275 35438
rect 7331 35382 7399 35438
rect 7455 35382 7523 35438
rect 7579 35382 7647 35438
rect 7703 35382 7713 35438
rect 7265 35314 7713 35382
rect 7265 35258 7275 35314
rect 7331 35258 7399 35314
rect 7455 35258 7523 35314
rect 7579 35258 7647 35314
rect 7703 35258 7713 35314
rect 7265 35190 7713 35258
rect 7265 35134 7275 35190
rect 7331 35134 7399 35190
rect 7455 35134 7523 35190
rect 7579 35134 7647 35190
rect 7703 35134 7713 35190
rect 7265 35066 7713 35134
rect 7265 35010 7275 35066
rect 7331 35010 7399 35066
rect 7455 35010 7523 35066
rect 7579 35010 7647 35066
rect 7703 35010 7713 35066
rect 7265 34942 7713 35010
rect 7265 34886 7275 34942
rect 7331 34886 7399 34942
rect 7455 34886 7523 34942
rect 7579 34886 7647 34942
rect 7703 34886 7713 34942
rect 7265 34818 7713 34886
rect 7265 34762 7275 34818
rect 7331 34762 7399 34818
rect 7455 34762 7523 34818
rect 7579 34762 7647 34818
rect 7703 34762 7713 34818
rect 7265 34694 7713 34762
rect 7265 34638 7275 34694
rect 7331 34638 7399 34694
rect 7455 34638 7523 34694
rect 7579 34638 7647 34694
rect 7703 34638 7713 34694
rect 7265 34570 7713 34638
rect 7265 34514 7275 34570
rect 7331 34514 7399 34570
rect 7455 34514 7523 34570
rect 7579 34514 7647 34570
rect 7703 34514 7713 34570
rect 7265 34446 7713 34514
rect 7265 34390 7275 34446
rect 7331 34390 7399 34446
rect 7455 34390 7523 34446
rect 7579 34390 7647 34446
rect 7703 34390 7713 34446
rect 7265 34322 7713 34390
rect 7265 34266 7275 34322
rect 7331 34266 7399 34322
rect 7455 34266 7523 34322
rect 7579 34266 7647 34322
rect 7703 34266 7713 34322
rect 7265 34198 7713 34266
rect 7265 34142 7275 34198
rect 7331 34142 7399 34198
rect 7455 34142 7523 34198
rect 7579 34142 7647 34198
rect 7703 34142 7713 34198
rect 7265 34074 7713 34142
rect 7265 34018 7275 34074
rect 7331 34018 7399 34074
rect 7455 34018 7523 34074
rect 7579 34018 7647 34074
rect 7703 34018 7713 34074
rect 7265 33950 7713 34018
rect 7265 33894 7275 33950
rect 7331 33894 7399 33950
rect 7455 33894 7523 33950
rect 7579 33894 7647 33950
rect 7703 33894 7713 33950
rect 7265 33826 7713 33894
rect 7265 33770 7275 33826
rect 7331 33770 7399 33826
rect 7455 33770 7523 33826
rect 7579 33770 7647 33826
rect 7703 33770 7713 33826
rect 7265 33702 7713 33770
rect 7265 33646 7275 33702
rect 7331 33646 7399 33702
rect 7455 33646 7523 33702
rect 7579 33646 7647 33702
rect 7703 33646 7713 33702
rect 7265 33636 7713 33646
rect 9927 36554 10127 36564
rect 9927 36498 9937 36554
rect 9993 36498 10061 36554
rect 10117 36498 10127 36554
rect 9927 36430 10127 36498
rect 9927 36374 9937 36430
rect 9993 36374 10061 36430
rect 10117 36374 10127 36430
rect 9927 36306 10127 36374
rect 9927 36250 9937 36306
rect 9993 36250 10061 36306
rect 10117 36250 10127 36306
rect 9927 36182 10127 36250
rect 9927 36126 9937 36182
rect 9993 36126 10061 36182
rect 10117 36126 10127 36182
rect 9927 36058 10127 36126
rect 9927 36002 9937 36058
rect 9993 36002 10061 36058
rect 10117 36002 10127 36058
rect 9927 35934 10127 36002
rect 9927 35878 9937 35934
rect 9993 35878 10061 35934
rect 10117 35878 10127 35934
rect 9927 35810 10127 35878
rect 9927 35754 9937 35810
rect 9993 35754 10061 35810
rect 10117 35754 10127 35810
rect 9927 35686 10127 35754
rect 9927 35630 9937 35686
rect 9993 35630 10061 35686
rect 10117 35630 10127 35686
rect 9927 35562 10127 35630
rect 9927 35506 9937 35562
rect 9993 35506 10061 35562
rect 10117 35506 10127 35562
rect 9927 35438 10127 35506
rect 9927 35382 9937 35438
rect 9993 35382 10061 35438
rect 10117 35382 10127 35438
rect 9927 35314 10127 35382
rect 9927 35258 9937 35314
rect 9993 35258 10061 35314
rect 10117 35258 10127 35314
rect 9927 35190 10127 35258
rect 9927 35134 9937 35190
rect 9993 35134 10061 35190
rect 10117 35134 10127 35190
rect 9927 35066 10127 35134
rect 9927 35010 9937 35066
rect 9993 35010 10061 35066
rect 10117 35010 10127 35066
rect 9927 34942 10127 35010
rect 9927 34886 9937 34942
rect 9993 34886 10061 34942
rect 10117 34886 10127 34942
rect 9927 34818 10127 34886
rect 9927 34762 9937 34818
rect 9993 34762 10061 34818
rect 10117 34762 10127 34818
rect 9927 34694 10127 34762
rect 9927 34638 9937 34694
rect 9993 34638 10061 34694
rect 10117 34638 10127 34694
rect 9927 34570 10127 34638
rect 9927 34514 9937 34570
rect 9993 34514 10061 34570
rect 10117 34514 10127 34570
rect 9927 34446 10127 34514
rect 9927 34390 9937 34446
rect 9993 34390 10061 34446
rect 10117 34390 10127 34446
rect 9927 34322 10127 34390
rect 9927 34266 9937 34322
rect 9993 34266 10061 34322
rect 10117 34266 10127 34322
rect 9927 34198 10127 34266
rect 9927 34142 9937 34198
rect 9993 34142 10061 34198
rect 10117 34142 10127 34198
rect 9927 34074 10127 34142
rect 9927 34018 9937 34074
rect 9993 34018 10061 34074
rect 10117 34018 10127 34074
rect 9927 33950 10127 34018
rect 9927 33894 9937 33950
rect 9993 33894 10061 33950
rect 10117 33894 10127 33950
rect 9927 33826 10127 33894
rect 9927 33770 9937 33826
rect 9993 33770 10061 33826
rect 10117 33770 10127 33826
rect 9927 33702 10127 33770
rect 9927 33646 9937 33702
rect 9993 33646 10061 33702
rect 10117 33646 10127 33702
rect 9927 33636 10127 33646
rect 12297 36554 12497 36564
rect 12297 36498 12307 36554
rect 12363 36498 12431 36554
rect 12487 36498 12497 36554
rect 12297 36430 12497 36498
rect 12297 36374 12307 36430
rect 12363 36374 12431 36430
rect 12487 36374 12497 36430
rect 12297 36306 12497 36374
rect 12297 36250 12307 36306
rect 12363 36250 12431 36306
rect 12487 36250 12497 36306
rect 12297 36182 12497 36250
rect 12297 36126 12307 36182
rect 12363 36126 12431 36182
rect 12487 36126 12497 36182
rect 12297 36058 12497 36126
rect 12297 36002 12307 36058
rect 12363 36002 12431 36058
rect 12487 36002 12497 36058
rect 12297 35934 12497 36002
rect 12297 35878 12307 35934
rect 12363 35878 12431 35934
rect 12487 35878 12497 35934
rect 12297 35810 12497 35878
rect 12297 35754 12307 35810
rect 12363 35754 12431 35810
rect 12487 35754 12497 35810
rect 12297 35686 12497 35754
rect 12297 35630 12307 35686
rect 12363 35630 12431 35686
rect 12487 35630 12497 35686
rect 12297 35562 12497 35630
rect 12297 35506 12307 35562
rect 12363 35506 12431 35562
rect 12487 35506 12497 35562
rect 12297 35438 12497 35506
rect 12297 35382 12307 35438
rect 12363 35382 12431 35438
rect 12487 35382 12497 35438
rect 12297 35314 12497 35382
rect 12297 35258 12307 35314
rect 12363 35258 12431 35314
rect 12487 35258 12497 35314
rect 12297 35190 12497 35258
rect 12297 35134 12307 35190
rect 12363 35134 12431 35190
rect 12487 35134 12497 35190
rect 12297 35066 12497 35134
rect 12297 35010 12307 35066
rect 12363 35010 12431 35066
rect 12487 35010 12497 35066
rect 12297 34942 12497 35010
rect 12297 34886 12307 34942
rect 12363 34886 12431 34942
rect 12487 34886 12497 34942
rect 12297 34818 12497 34886
rect 12297 34762 12307 34818
rect 12363 34762 12431 34818
rect 12487 34762 12497 34818
rect 12297 34694 12497 34762
rect 12297 34638 12307 34694
rect 12363 34638 12431 34694
rect 12487 34638 12497 34694
rect 12297 34570 12497 34638
rect 12297 34514 12307 34570
rect 12363 34514 12431 34570
rect 12487 34514 12497 34570
rect 12297 34446 12497 34514
rect 12297 34390 12307 34446
rect 12363 34390 12431 34446
rect 12487 34390 12497 34446
rect 12297 34322 12497 34390
rect 12297 34266 12307 34322
rect 12363 34266 12431 34322
rect 12487 34266 12497 34322
rect 12297 34198 12497 34266
rect 12297 34142 12307 34198
rect 12363 34142 12431 34198
rect 12487 34142 12497 34198
rect 12297 34074 12497 34142
rect 12297 34018 12307 34074
rect 12363 34018 12431 34074
rect 12487 34018 12497 34074
rect 12297 33950 12497 34018
rect 12297 33894 12307 33950
rect 12363 33894 12431 33950
rect 12487 33894 12497 33950
rect 12297 33826 12497 33894
rect 12297 33770 12307 33826
rect 12363 33770 12431 33826
rect 12487 33770 12497 33826
rect 12297 33702 12497 33770
rect 12297 33646 12307 33702
rect 12363 33646 12431 33702
rect 12487 33646 12497 33702
rect 12297 33636 12497 33646
rect 305 33354 2117 33364
rect 305 33298 315 33354
rect 371 33298 439 33354
rect 495 33298 563 33354
rect 619 33298 687 33354
rect 743 33298 811 33354
rect 867 33298 935 33354
rect 991 33298 1059 33354
rect 1115 33298 1183 33354
rect 1239 33298 1307 33354
rect 1363 33298 1431 33354
rect 1487 33298 1555 33354
rect 1611 33298 1679 33354
rect 1735 33298 1803 33354
rect 1859 33298 1927 33354
rect 1983 33298 2051 33354
rect 2107 33298 2117 33354
rect 305 33230 2117 33298
rect 305 33174 315 33230
rect 371 33174 439 33230
rect 495 33174 563 33230
rect 619 33174 687 33230
rect 743 33174 811 33230
rect 867 33174 935 33230
rect 991 33174 1059 33230
rect 1115 33174 1183 33230
rect 1239 33174 1307 33230
rect 1363 33174 1431 33230
rect 1487 33174 1555 33230
rect 1611 33174 1679 33230
rect 1735 33174 1803 33230
rect 1859 33174 1927 33230
rect 1983 33174 2051 33230
rect 2107 33174 2117 33230
rect 305 33106 2117 33174
rect 305 33050 315 33106
rect 371 33050 439 33106
rect 495 33050 563 33106
rect 619 33050 687 33106
rect 743 33050 811 33106
rect 867 33050 935 33106
rect 991 33050 1059 33106
rect 1115 33050 1183 33106
rect 1239 33050 1307 33106
rect 1363 33050 1431 33106
rect 1487 33050 1555 33106
rect 1611 33050 1679 33106
rect 1735 33050 1803 33106
rect 1859 33050 1927 33106
rect 1983 33050 2051 33106
rect 2107 33050 2117 33106
rect 305 32982 2117 33050
rect 305 32926 315 32982
rect 371 32926 439 32982
rect 495 32926 563 32982
rect 619 32926 687 32982
rect 743 32926 811 32982
rect 867 32926 935 32982
rect 991 32926 1059 32982
rect 1115 32926 1183 32982
rect 1239 32926 1307 32982
rect 1363 32926 1431 32982
rect 1487 32926 1555 32982
rect 1611 32926 1679 32982
rect 1735 32926 1803 32982
rect 1859 32926 1927 32982
rect 1983 32926 2051 32982
rect 2107 32926 2117 32982
rect 305 32858 2117 32926
rect 305 32802 315 32858
rect 371 32802 439 32858
rect 495 32802 563 32858
rect 619 32802 687 32858
rect 743 32802 811 32858
rect 867 32802 935 32858
rect 991 32802 1059 32858
rect 1115 32802 1183 32858
rect 1239 32802 1307 32858
rect 1363 32802 1431 32858
rect 1487 32802 1555 32858
rect 1611 32802 1679 32858
rect 1735 32802 1803 32858
rect 1859 32802 1927 32858
rect 1983 32802 2051 32858
rect 2107 32802 2117 32858
rect 305 32734 2117 32802
rect 305 32678 315 32734
rect 371 32678 439 32734
rect 495 32678 563 32734
rect 619 32678 687 32734
rect 743 32678 811 32734
rect 867 32678 935 32734
rect 991 32678 1059 32734
rect 1115 32678 1183 32734
rect 1239 32678 1307 32734
rect 1363 32678 1431 32734
rect 1487 32678 1555 32734
rect 1611 32678 1679 32734
rect 1735 32678 1803 32734
rect 1859 32678 1927 32734
rect 1983 32678 2051 32734
rect 2107 32678 2117 32734
rect 305 32610 2117 32678
rect 305 32554 315 32610
rect 371 32554 439 32610
rect 495 32554 563 32610
rect 619 32554 687 32610
rect 743 32554 811 32610
rect 867 32554 935 32610
rect 991 32554 1059 32610
rect 1115 32554 1183 32610
rect 1239 32554 1307 32610
rect 1363 32554 1431 32610
rect 1487 32554 1555 32610
rect 1611 32554 1679 32610
rect 1735 32554 1803 32610
rect 1859 32554 1927 32610
rect 1983 32554 2051 32610
rect 2107 32554 2117 32610
rect 305 32486 2117 32554
rect 305 32430 315 32486
rect 371 32430 439 32486
rect 495 32430 563 32486
rect 619 32430 687 32486
rect 743 32430 811 32486
rect 867 32430 935 32486
rect 991 32430 1059 32486
rect 1115 32430 1183 32486
rect 1239 32430 1307 32486
rect 1363 32430 1431 32486
rect 1487 32430 1555 32486
rect 1611 32430 1679 32486
rect 1735 32430 1803 32486
rect 1859 32430 1927 32486
rect 1983 32430 2051 32486
rect 2107 32430 2117 32486
rect 305 32362 2117 32430
rect 305 32306 315 32362
rect 371 32306 439 32362
rect 495 32306 563 32362
rect 619 32306 687 32362
rect 743 32306 811 32362
rect 867 32306 935 32362
rect 991 32306 1059 32362
rect 1115 32306 1183 32362
rect 1239 32306 1307 32362
rect 1363 32306 1431 32362
rect 1487 32306 1555 32362
rect 1611 32306 1679 32362
rect 1735 32306 1803 32362
rect 1859 32306 1927 32362
rect 1983 32306 2051 32362
rect 2107 32306 2117 32362
rect 305 32238 2117 32306
rect 305 32182 315 32238
rect 371 32182 439 32238
rect 495 32182 563 32238
rect 619 32182 687 32238
rect 743 32182 811 32238
rect 867 32182 935 32238
rect 991 32182 1059 32238
rect 1115 32182 1183 32238
rect 1239 32182 1307 32238
rect 1363 32182 1431 32238
rect 1487 32182 1555 32238
rect 1611 32182 1679 32238
rect 1735 32182 1803 32238
rect 1859 32182 1927 32238
rect 1983 32182 2051 32238
rect 2107 32182 2117 32238
rect 305 32114 2117 32182
rect 305 32058 315 32114
rect 371 32058 439 32114
rect 495 32058 563 32114
rect 619 32058 687 32114
rect 743 32058 811 32114
rect 867 32058 935 32114
rect 991 32058 1059 32114
rect 1115 32058 1183 32114
rect 1239 32058 1307 32114
rect 1363 32058 1431 32114
rect 1487 32058 1555 32114
rect 1611 32058 1679 32114
rect 1735 32058 1803 32114
rect 1859 32058 1927 32114
rect 1983 32058 2051 32114
rect 2107 32058 2117 32114
rect 305 31990 2117 32058
rect 305 31934 315 31990
rect 371 31934 439 31990
rect 495 31934 563 31990
rect 619 31934 687 31990
rect 743 31934 811 31990
rect 867 31934 935 31990
rect 991 31934 1059 31990
rect 1115 31934 1183 31990
rect 1239 31934 1307 31990
rect 1363 31934 1431 31990
rect 1487 31934 1555 31990
rect 1611 31934 1679 31990
rect 1735 31934 1803 31990
rect 1859 31934 1927 31990
rect 1983 31934 2051 31990
rect 2107 31934 2117 31990
rect 305 31866 2117 31934
rect 305 31810 315 31866
rect 371 31810 439 31866
rect 495 31810 563 31866
rect 619 31810 687 31866
rect 743 31810 811 31866
rect 867 31810 935 31866
rect 991 31810 1059 31866
rect 1115 31810 1183 31866
rect 1239 31810 1307 31866
rect 1363 31810 1431 31866
rect 1487 31810 1555 31866
rect 1611 31810 1679 31866
rect 1735 31810 1803 31866
rect 1859 31810 1927 31866
rect 1983 31810 2051 31866
rect 2107 31810 2117 31866
rect 305 31742 2117 31810
rect 305 31686 315 31742
rect 371 31686 439 31742
rect 495 31686 563 31742
rect 619 31686 687 31742
rect 743 31686 811 31742
rect 867 31686 935 31742
rect 991 31686 1059 31742
rect 1115 31686 1183 31742
rect 1239 31686 1307 31742
rect 1363 31686 1431 31742
rect 1487 31686 1555 31742
rect 1611 31686 1679 31742
rect 1735 31686 1803 31742
rect 1859 31686 1927 31742
rect 1983 31686 2051 31742
rect 2107 31686 2117 31742
rect 305 31618 2117 31686
rect 305 31562 315 31618
rect 371 31562 439 31618
rect 495 31562 563 31618
rect 619 31562 687 31618
rect 743 31562 811 31618
rect 867 31562 935 31618
rect 991 31562 1059 31618
rect 1115 31562 1183 31618
rect 1239 31562 1307 31618
rect 1363 31562 1431 31618
rect 1487 31562 1555 31618
rect 1611 31562 1679 31618
rect 1735 31562 1803 31618
rect 1859 31562 1927 31618
rect 1983 31562 2051 31618
rect 2107 31562 2117 31618
rect 305 31494 2117 31562
rect 305 31438 315 31494
rect 371 31438 439 31494
rect 495 31438 563 31494
rect 619 31438 687 31494
rect 743 31438 811 31494
rect 867 31438 935 31494
rect 991 31438 1059 31494
rect 1115 31438 1183 31494
rect 1239 31438 1307 31494
rect 1363 31438 1431 31494
rect 1487 31438 1555 31494
rect 1611 31438 1679 31494
rect 1735 31438 1803 31494
rect 1859 31438 1927 31494
rect 1983 31438 2051 31494
rect 2107 31438 2117 31494
rect 305 31370 2117 31438
rect 305 31314 315 31370
rect 371 31314 439 31370
rect 495 31314 563 31370
rect 619 31314 687 31370
rect 743 31314 811 31370
rect 867 31314 935 31370
rect 991 31314 1059 31370
rect 1115 31314 1183 31370
rect 1239 31314 1307 31370
rect 1363 31314 1431 31370
rect 1487 31314 1555 31370
rect 1611 31314 1679 31370
rect 1735 31314 1803 31370
rect 1859 31314 1927 31370
rect 1983 31314 2051 31370
rect 2107 31314 2117 31370
rect 305 31246 2117 31314
rect 305 31190 315 31246
rect 371 31190 439 31246
rect 495 31190 563 31246
rect 619 31190 687 31246
rect 743 31190 811 31246
rect 867 31190 935 31246
rect 991 31190 1059 31246
rect 1115 31190 1183 31246
rect 1239 31190 1307 31246
rect 1363 31190 1431 31246
rect 1487 31190 1555 31246
rect 1611 31190 1679 31246
rect 1735 31190 1803 31246
rect 1859 31190 1927 31246
rect 1983 31190 2051 31246
rect 2107 31190 2117 31246
rect 305 31122 2117 31190
rect 305 31066 315 31122
rect 371 31066 439 31122
rect 495 31066 563 31122
rect 619 31066 687 31122
rect 743 31066 811 31122
rect 867 31066 935 31122
rect 991 31066 1059 31122
rect 1115 31066 1183 31122
rect 1239 31066 1307 31122
rect 1363 31066 1431 31122
rect 1487 31066 1555 31122
rect 1611 31066 1679 31122
rect 1735 31066 1803 31122
rect 1859 31066 1927 31122
rect 1983 31066 2051 31122
rect 2107 31066 2117 31122
rect 305 30998 2117 31066
rect 305 30942 315 30998
rect 371 30942 439 30998
rect 495 30942 563 30998
rect 619 30942 687 30998
rect 743 30942 811 30998
rect 867 30942 935 30998
rect 991 30942 1059 30998
rect 1115 30942 1183 30998
rect 1239 30942 1307 30998
rect 1363 30942 1431 30998
rect 1487 30942 1555 30998
rect 1611 30942 1679 30998
rect 1735 30942 1803 30998
rect 1859 30942 1927 30998
rect 1983 30942 2051 30998
rect 2107 30942 2117 30998
rect 305 30874 2117 30942
rect 305 30818 315 30874
rect 371 30818 439 30874
rect 495 30818 563 30874
rect 619 30818 687 30874
rect 743 30818 811 30874
rect 867 30818 935 30874
rect 991 30818 1059 30874
rect 1115 30818 1183 30874
rect 1239 30818 1307 30874
rect 1363 30818 1431 30874
rect 1487 30818 1555 30874
rect 1611 30818 1679 30874
rect 1735 30818 1803 30874
rect 1859 30818 1927 30874
rect 1983 30818 2051 30874
rect 2107 30818 2117 30874
rect 305 30750 2117 30818
rect 305 30694 315 30750
rect 371 30694 439 30750
rect 495 30694 563 30750
rect 619 30694 687 30750
rect 743 30694 811 30750
rect 867 30694 935 30750
rect 991 30694 1059 30750
rect 1115 30694 1183 30750
rect 1239 30694 1307 30750
rect 1363 30694 1431 30750
rect 1487 30694 1555 30750
rect 1611 30694 1679 30750
rect 1735 30694 1803 30750
rect 1859 30694 1927 30750
rect 1983 30694 2051 30750
rect 2107 30694 2117 30750
rect 305 30626 2117 30694
rect 305 30570 315 30626
rect 371 30570 439 30626
rect 495 30570 563 30626
rect 619 30570 687 30626
rect 743 30570 811 30626
rect 867 30570 935 30626
rect 991 30570 1059 30626
rect 1115 30570 1183 30626
rect 1239 30570 1307 30626
rect 1363 30570 1431 30626
rect 1487 30570 1555 30626
rect 1611 30570 1679 30626
rect 1735 30570 1803 30626
rect 1859 30570 1927 30626
rect 1983 30570 2051 30626
rect 2107 30570 2117 30626
rect 305 30502 2117 30570
rect 305 30446 315 30502
rect 371 30446 439 30502
rect 495 30446 563 30502
rect 619 30446 687 30502
rect 743 30446 811 30502
rect 867 30446 935 30502
rect 991 30446 1059 30502
rect 1115 30446 1183 30502
rect 1239 30446 1307 30502
rect 1363 30446 1431 30502
rect 1487 30446 1555 30502
rect 1611 30446 1679 30502
rect 1735 30446 1803 30502
rect 1859 30446 1927 30502
rect 1983 30446 2051 30502
rect 2107 30446 2117 30502
rect 305 30436 2117 30446
rect 2798 33354 4734 33364
rect 2798 33298 2808 33354
rect 2864 33298 2932 33354
rect 2988 33298 3056 33354
rect 3112 33298 3180 33354
rect 3236 33298 3304 33354
rect 3360 33298 3428 33354
rect 3484 33298 3552 33354
rect 3608 33298 3676 33354
rect 3732 33298 3800 33354
rect 3856 33298 3924 33354
rect 3980 33298 4048 33354
rect 4104 33298 4172 33354
rect 4228 33298 4296 33354
rect 4352 33298 4420 33354
rect 4476 33298 4544 33354
rect 4600 33298 4668 33354
rect 4724 33298 4734 33354
rect 2798 33230 4734 33298
rect 2798 33174 2808 33230
rect 2864 33174 2932 33230
rect 2988 33174 3056 33230
rect 3112 33174 3180 33230
rect 3236 33174 3304 33230
rect 3360 33174 3428 33230
rect 3484 33174 3552 33230
rect 3608 33174 3676 33230
rect 3732 33174 3800 33230
rect 3856 33174 3924 33230
rect 3980 33174 4048 33230
rect 4104 33174 4172 33230
rect 4228 33174 4296 33230
rect 4352 33174 4420 33230
rect 4476 33174 4544 33230
rect 4600 33174 4668 33230
rect 4724 33174 4734 33230
rect 2798 33106 4734 33174
rect 2798 33050 2808 33106
rect 2864 33050 2932 33106
rect 2988 33050 3056 33106
rect 3112 33050 3180 33106
rect 3236 33050 3304 33106
rect 3360 33050 3428 33106
rect 3484 33050 3552 33106
rect 3608 33050 3676 33106
rect 3732 33050 3800 33106
rect 3856 33050 3924 33106
rect 3980 33050 4048 33106
rect 4104 33050 4172 33106
rect 4228 33050 4296 33106
rect 4352 33050 4420 33106
rect 4476 33050 4544 33106
rect 4600 33050 4668 33106
rect 4724 33050 4734 33106
rect 2798 32982 4734 33050
rect 2798 32926 2808 32982
rect 2864 32926 2932 32982
rect 2988 32926 3056 32982
rect 3112 32926 3180 32982
rect 3236 32926 3304 32982
rect 3360 32926 3428 32982
rect 3484 32926 3552 32982
rect 3608 32926 3676 32982
rect 3732 32926 3800 32982
rect 3856 32926 3924 32982
rect 3980 32926 4048 32982
rect 4104 32926 4172 32982
rect 4228 32926 4296 32982
rect 4352 32926 4420 32982
rect 4476 32926 4544 32982
rect 4600 32926 4668 32982
rect 4724 32926 4734 32982
rect 2798 32858 4734 32926
rect 2798 32802 2808 32858
rect 2864 32802 2932 32858
rect 2988 32802 3056 32858
rect 3112 32802 3180 32858
rect 3236 32802 3304 32858
rect 3360 32802 3428 32858
rect 3484 32802 3552 32858
rect 3608 32802 3676 32858
rect 3732 32802 3800 32858
rect 3856 32802 3924 32858
rect 3980 32802 4048 32858
rect 4104 32802 4172 32858
rect 4228 32802 4296 32858
rect 4352 32802 4420 32858
rect 4476 32802 4544 32858
rect 4600 32802 4668 32858
rect 4724 32802 4734 32858
rect 2798 32734 4734 32802
rect 2798 32678 2808 32734
rect 2864 32678 2932 32734
rect 2988 32678 3056 32734
rect 3112 32678 3180 32734
rect 3236 32678 3304 32734
rect 3360 32678 3428 32734
rect 3484 32678 3552 32734
rect 3608 32678 3676 32734
rect 3732 32678 3800 32734
rect 3856 32678 3924 32734
rect 3980 32678 4048 32734
rect 4104 32678 4172 32734
rect 4228 32678 4296 32734
rect 4352 32678 4420 32734
rect 4476 32678 4544 32734
rect 4600 32678 4668 32734
rect 4724 32678 4734 32734
rect 2798 32610 4734 32678
rect 2798 32554 2808 32610
rect 2864 32554 2932 32610
rect 2988 32554 3056 32610
rect 3112 32554 3180 32610
rect 3236 32554 3304 32610
rect 3360 32554 3428 32610
rect 3484 32554 3552 32610
rect 3608 32554 3676 32610
rect 3732 32554 3800 32610
rect 3856 32554 3924 32610
rect 3980 32554 4048 32610
rect 4104 32554 4172 32610
rect 4228 32554 4296 32610
rect 4352 32554 4420 32610
rect 4476 32554 4544 32610
rect 4600 32554 4668 32610
rect 4724 32554 4734 32610
rect 2798 32486 4734 32554
rect 2798 32430 2808 32486
rect 2864 32430 2932 32486
rect 2988 32430 3056 32486
rect 3112 32430 3180 32486
rect 3236 32430 3304 32486
rect 3360 32430 3428 32486
rect 3484 32430 3552 32486
rect 3608 32430 3676 32486
rect 3732 32430 3800 32486
rect 3856 32430 3924 32486
rect 3980 32430 4048 32486
rect 4104 32430 4172 32486
rect 4228 32430 4296 32486
rect 4352 32430 4420 32486
rect 4476 32430 4544 32486
rect 4600 32430 4668 32486
rect 4724 32430 4734 32486
rect 2798 32362 4734 32430
rect 2798 32306 2808 32362
rect 2864 32306 2932 32362
rect 2988 32306 3056 32362
rect 3112 32306 3180 32362
rect 3236 32306 3304 32362
rect 3360 32306 3428 32362
rect 3484 32306 3552 32362
rect 3608 32306 3676 32362
rect 3732 32306 3800 32362
rect 3856 32306 3924 32362
rect 3980 32306 4048 32362
rect 4104 32306 4172 32362
rect 4228 32306 4296 32362
rect 4352 32306 4420 32362
rect 4476 32306 4544 32362
rect 4600 32306 4668 32362
rect 4724 32306 4734 32362
rect 2798 32238 4734 32306
rect 2798 32182 2808 32238
rect 2864 32182 2932 32238
rect 2988 32182 3056 32238
rect 3112 32182 3180 32238
rect 3236 32182 3304 32238
rect 3360 32182 3428 32238
rect 3484 32182 3552 32238
rect 3608 32182 3676 32238
rect 3732 32182 3800 32238
rect 3856 32182 3924 32238
rect 3980 32182 4048 32238
rect 4104 32182 4172 32238
rect 4228 32182 4296 32238
rect 4352 32182 4420 32238
rect 4476 32182 4544 32238
rect 4600 32182 4668 32238
rect 4724 32182 4734 32238
rect 2798 32114 4734 32182
rect 2798 32058 2808 32114
rect 2864 32058 2932 32114
rect 2988 32058 3056 32114
rect 3112 32058 3180 32114
rect 3236 32058 3304 32114
rect 3360 32058 3428 32114
rect 3484 32058 3552 32114
rect 3608 32058 3676 32114
rect 3732 32058 3800 32114
rect 3856 32058 3924 32114
rect 3980 32058 4048 32114
rect 4104 32058 4172 32114
rect 4228 32058 4296 32114
rect 4352 32058 4420 32114
rect 4476 32058 4544 32114
rect 4600 32058 4668 32114
rect 4724 32058 4734 32114
rect 2798 31990 4734 32058
rect 2798 31934 2808 31990
rect 2864 31934 2932 31990
rect 2988 31934 3056 31990
rect 3112 31934 3180 31990
rect 3236 31934 3304 31990
rect 3360 31934 3428 31990
rect 3484 31934 3552 31990
rect 3608 31934 3676 31990
rect 3732 31934 3800 31990
rect 3856 31934 3924 31990
rect 3980 31934 4048 31990
rect 4104 31934 4172 31990
rect 4228 31934 4296 31990
rect 4352 31934 4420 31990
rect 4476 31934 4544 31990
rect 4600 31934 4668 31990
rect 4724 31934 4734 31990
rect 2798 31866 4734 31934
rect 2798 31810 2808 31866
rect 2864 31810 2932 31866
rect 2988 31810 3056 31866
rect 3112 31810 3180 31866
rect 3236 31810 3304 31866
rect 3360 31810 3428 31866
rect 3484 31810 3552 31866
rect 3608 31810 3676 31866
rect 3732 31810 3800 31866
rect 3856 31810 3924 31866
rect 3980 31810 4048 31866
rect 4104 31810 4172 31866
rect 4228 31810 4296 31866
rect 4352 31810 4420 31866
rect 4476 31810 4544 31866
rect 4600 31810 4668 31866
rect 4724 31810 4734 31866
rect 2798 31742 4734 31810
rect 2798 31686 2808 31742
rect 2864 31686 2932 31742
rect 2988 31686 3056 31742
rect 3112 31686 3180 31742
rect 3236 31686 3304 31742
rect 3360 31686 3428 31742
rect 3484 31686 3552 31742
rect 3608 31686 3676 31742
rect 3732 31686 3800 31742
rect 3856 31686 3924 31742
rect 3980 31686 4048 31742
rect 4104 31686 4172 31742
rect 4228 31686 4296 31742
rect 4352 31686 4420 31742
rect 4476 31686 4544 31742
rect 4600 31686 4668 31742
rect 4724 31686 4734 31742
rect 2798 31618 4734 31686
rect 2798 31562 2808 31618
rect 2864 31562 2932 31618
rect 2988 31562 3056 31618
rect 3112 31562 3180 31618
rect 3236 31562 3304 31618
rect 3360 31562 3428 31618
rect 3484 31562 3552 31618
rect 3608 31562 3676 31618
rect 3732 31562 3800 31618
rect 3856 31562 3924 31618
rect 3980 31562 4048 31618
rect 4104 31562 4172 31618
rect 4228 31562 4296 31618
rect 4352 31562 4420 31618
rect 4476 31562 4544 31618
rect 4600 31562 4668 31618
rect 4724 31562 4734 31618
rect 2798 31494 4734 31562
rect 2798 31438 2808 31494
rect 2864 31438 2932 31494
rect 2988 31438 3056 31494
rect 3112 31438 3180 31494
rect 3236 31438 3304 31494
rect 3360 31438 3428 31494
rect 3484 31438 3552 31494
rect 3608 31438 3676 31494
rect 3732 31438 3800 31494
rect 3856 31438 3924 31494
rect 3980 31438 4048 31494
rect 4104 31438 4172 31494
rect 4228 31438 4296 31494
rect 4352 31438 4420 31494
rect 4476 31438 4544 31494
rect 4600 31438 4668 31494
rect 4724 31438 4734 31494
rect 2798 31370 4734 31438
rect 2798 31314 2808 31370
rect 2864 31314 2932 31370
rect 2988 31314 3056 31370
rect 3112 31314 3180 31370
rect 3236 31314 3304 31370
rect 3360 31314 3428 31370
rect 3484 31314 3552 31370
rect 3608 31314 3676 31370
rect 3732 31314 3800 31370
rect 3856 31314 3924 31370
rect 3980 31314 4048 31370
rect 4104 31314 4172 31370
rect 4228 31314 4296 31370
rect 4352 31314 4420 31370
rect 4476 31314 4544 31370
rect 4600 31314 4668 31370
rect 4724 31314 4734 31370
rect 2798 31246 4734 31314
rect 2798 31190 2808 31246
rect 2864 31190 2932 31246
rect 2988 31190 3056 31246
rect 3112 31190 3180 31246
rect 3236 31190 3304 31246
rect 3360 31190 3428 31246
rect 3484 31190 3552 31246
rect 3608 31190 3676 31246
rect 3732 31190 3800 31246
rect 3856 31190 3924 31246
rect 3980 31190 4048 31246
rect 4104 31190 4172 31246
rect 4228 31190 4296 31246
rect 4352 31190 4420 31246
rect 4476 31190 4544 31246
rect 4600 31190 4668 31246
rect 4724 31190 4734 31246
rect 2798 31122 4734 31190
rect 2798 31066 2808 31122
rect 2864 31066 2932 31122
rect 2988 31066 3056 31122
rect 3112 31066 3180 31122
rect 3236 31066 3304 31122
rect 3360 31066 3428 31122
rect 3484 31066 3552 31122
rect 3608 31066 3676 31122
rect 3732 31066 3800 31122
rect 3856 31066 3924 31122
rect 3980 31066 4048 31122
rect 4104 31066 4172 31122
rect 4228 31066 4296 31122
rect 4352 31066 4420 31122
rect 4476 31066 4544 31122
rect 4600 31066 4668 31122
rect 4724 31066 4734 31122
rect 2798 30998 4734 31066
rect 2798 30942 2808 30998
rect 2864 30942 2932 30998
rect 2988 30942 3056 30998
rect 3112 30942 3180 30998
rect 3236 30942 3304 30998
rect 3360 30942 3428 30998
rect 3484 30942 3552 30998
rect 3608 30942 3676 30998
rect 3732 30942 3800 30998
rect 3856 30942 3924 30998
rect 3980 30942 4048 30998
rect 4104 30942 4172 30998
rect 4228 30942 4296 30998
rect 4352 30942 4420 30998
rect 4476 30942 4544 30998
rect 4600 30942 4668 30998
rect 4724 30942 4734 30998
rect 2798 30874 4734 30942
rect 2798 30818 2808 30874
rect 2864 30818 2932 30874
rect 2988 30818 3056 30874
rect 3112 30818 3180 30874
rect 3236 30818 3304 30874
rect 3360 30818 3428 30874
rect 3484 30818 3552 30874
rect 3608 30818 3676 30874
rect 3732 30818 3800 30874
rect 3856 30818 3924 30874
rect 3980 30818 4048 30874
rect 4104 30818 4172 30874
rect 4228 30818 4296 30874
rect 4352 30818 4420 30874
rect 4476 30818 4544 30874
rect 4600 30818 4668 30874
rect 4724 30818 4734 30874
rect 2798 30750 4734 30818
rect 2798 30694 2808 30750
rect 2864 30694 2932 30750
rect 2988 30694 3056 30750
rect 3112 30694 3180 30750
rect 3236 30694 3304 30750
rect 3360 30694 3428 30750
rect 3484 30694 3552 30750
rect 3608 30694 3676 30750
rect 3732 30694 3800 30750
rect 3856 30694 3924 30750
rect 3980 30694 4048 30750
rect 4104 30694 4172 30750
rect 4228 30694 4296 30750
rect 4352 30694 4420 30750
rect 4476 30694 4544 30750
rect 4600 30694 4668 30750
rect 4724 30694 4734 30750
rect 2798 30626 4734 30694
rect 2798 30570 2808 30626
rect 2864 30570 2932 30626
rect 2988 30570 3056 30626
rect 3112 30570 3180 30626
rect 3236 30570 3304 30626
rect 3360 30570 3428 30626
rect 3484 30570 3552 30626
rect 3608 30570 3676 30626
rect 3732 30570 3800 30626
rect 3856 30570 3924 30626
rect 3980 30570 4048 30626
rect 4104 30570 4172 30626
rect 4228 30570 4296 30626
rect 4352 30570 4420 30626
rect 4476 30570 4544 30626
rect 4600 30570 4668 30626
rect 4724 30570 4734 30626
rect 2798 30502 4734 30570
rect 2798 30446 2808 30502
rect 2864 30446 2932 30502
rect 2988 30446 3056 30502
rect 3112 30446 3180 30502
rect 3236 30446 3304 30502
rect 3360 30446 3428 30502
rect 3484 30446 3552 30502
rect 3608 30446 3676 30502
rect 3732 30446 3800 30502
rect 3856 30446 3924 30502
rect 3980 30446 4048 30502
rect 4104 30446 4172 30502
rect 4228 30446 4296 30502
rect 4352 30446 4420 30502
rect 4476 30446 4544 30502
rect 4600 30446 4668 30502
rect 4724 30446 4734 30502
rect 2798 30436 4734 30446
rect 5168 33354 7104 33364
rect 5168 33298 5178 33354
rect 5234 33298 5302 33354
rect 5358 33298 5426 33354
rect 5482 33298 5550 33354
rect 5606 33298 5674 33354
rect 5730 33298 5798 33354
rect 5854 33298 5922 33354
rect 5978 33298 6046 33354
rect 6102 33298 6170 33354
rect 6226 33298 6294 33354
rect 6350 33298 6418 33354
rect 6474 33298 6542 33354
rect 6598 33298 6666 33354
rect 6722 33298 6790 33354
rect 6846 33298 6914 33354
rect 6970 33298 7038 33354
rect 7094 33298 7104 33354
rect 5168 33230 7104 33298
rect 5168 33174 5178 33230
rect 5234 33174 5302 33230
rect 5358 33174 5426 33230
rect 5482 33174 5550 33230
rect 5606 33174 5674 33230
rect 5730 33174 5798 33230
rect 5854 33174 5922 33230
rect 5978 33174 6046 33230
rect 6102 33174 6170 33230
rect 6226 33174 6294 33230
rect 6350 33174 6418 33230
rect 6474 33174 6542 33230
rect 6598 33174 6666 33230
rect 6722 33174 6790 33230
rect 6846 33174 6914 33230
rect 6970 33174 7038 33230
rect 7094 33174 7104 33230
rect 5168 33106 7104 33174
rect 5168 33050 5178 33106
rect 5234 33050 5302 33106
rect 5358 33050 5426 33106
rect 5482 33050 5550 33106
rect 5606 33050 5674 33106
rect 5730 33050 5798 33106
rect 5854 33050 5922 33106
rect 5978 33050 6046 33106
rect 6102 33050 6170 33106
rect 6226 33050 6294 33106
rect 6350 33050 6418 33106
rect 6474 33050 6542 33106
rect 6598 33050 6666 33106
rect 6722 33050 6790 33106
rect 6846 33050 6914 33106
rect 6970 33050 7038 33106
rect 7094 33050 7104 33106
rect 5168 32982 7104 33050
rect 5168 32926 5178 32982
rect 5234 32926 5302 32982
rect 5358 32926 5426 32982
rect 5482 32926 5550 32982
rect 5606 32926 5674 32982
rect 5730 32926 5798 32982
rect 5854 32926 5922 32982
rect 5978 32926 6046 32982
rect 6102 32926 6170 32982
rect 6226 32926 6294 32982
rect 6350 32926 6418 32982
rect 6474 32926 6542 32982
rect 6598 32926 6666 32982
rect 6722 32926 6790 32982
rect 6846 32926 6914 32982
rect 6970 32926 7038 32982
rect 7094 32926 7104 32982
rect 5168 32858 7104 32926
rect 5168 32802 5178 32858
rect 5234 32802 5302 32858
rect 5358 32802 5426 32858
rect 5482 32802 5550 32858
rect 5606 32802 5674 32858
rect 5730 32802 5798 32858
rect 5854 32802 5922 32858
rect 5978 32802 6046 32858
rect 6102 32802 6170 32858
rect 6226 32802 6294 32858
rect 6350 32802 6418 32858
rect 6474 32802 6542 32858
rect 6598 32802 6666 32858
rect 6722 32802 6790 32858
rect 6846 32802 6914 32858
rect 6970 32802 7038 32858
rect 7094 32802 7104 32858
rect 5168 32734 7104 32802
rect 5168 32678 5178 32734
rect 5234 32678 5302 32734
rect 5358 32678 5426 32734
rect 5482 32678 5550 32734
rect 5606 32678 5674 32734
rect 5730 32678 5798 32734
rect 5854 32678 5922 32734
rect 5978 32678 6046 32734
rect 6102 32678 6170 32734
rect 6226 32678 6294 32734
rect 6350 32678 6418 32734
rect 6474 32678 6542 32734
rect 6598 32678 6666 32734
rect 6722 32678 6790 32734
rect 6846 32678 6914 32734
rect 6970 32678 7038 32734
rect 7094 32678 7104 32734
rect 5168 32610 7104 32678
rect 5168 32554 5178 32610
rect 5234 32554 5302 32610
rect 5358 32554 5426 32610
rect 5482 32554 5550 32610
rect 5606 32554 5674 32610
rect 5730 32554 5798 32610
rect 5854 32554 5922 32610
rect 5978 32554 6046 32610
rect 6102 32554 6170 32610
rect 6226 32554 6294 32610
rect 6350 32554 6418 32610
rect 6474 32554 6542 32610
rect 6598 32554 6666 32610
rect 6722 32554 6790 32610
rect 6846 32554 6914 32610
rect 6970 32554 7038 32610
rect 7094 32554 7104 32610
rect 5168 32486 7104 32554
rect 5168 32430 5178 32486
rect 5234 32430 5302 32486
rect 5358 32430 5426 32486
rect 5482 32430 5550 32486
rect 5606 32430 5674 32486
rect 5730 32430 5798 32486
rect 5854 32430 5922 32486
rect 5978 32430 6046 32486
rect 6102 32430 6170 32486
rect 6226 32430 6294 32486
rect 6350 32430 6418 32486
rect 6474 32430 6542 32486
rect 6598 32430 6666 32486
rect 6722 32430 6790 32486
rect 6846 32430 6914 32486
rect 6970 32430 7038 32486
rect 7094 32430 7104 32486
rect 5168 32362 7104 32430
rect 5168 32306 5178 32362
rect 5234 32306 5302 32362
rect 5358 32306 5426 32362
rect 5482 32306 5550 32362
rect 5606 32306 5674 32362
rect 5730 32306 5798 32362
rect 5854 32306 5922 32362
rect 5978 32306 6046 32362
rect 6102 32306 6170 32362
rect 6226 32306 6294 32362
rect 6350 32306 6418 32362
rect 6474 32306 6542 32362
rect 6598 32306 6666 32362
rect 6722 32306 6790 32362
rect 6846 32306 6914 32362
rect 6970 32306 7038 32362
rect 7094 32306 7104 32362
rect 5168 32238 7104 32306
rect 5168 32182 5178 32238
rect 5234 32182 5302 32238
rect 5358 32182 5426 32238
rect 5482 32182 5550 32238
rect 5606 32182 5674 32238
rect 5730 32182 5798 32238
rect 5854 32182 5922 32238
rect 5978 32182 6046 32238
rect 6102 32182 6170 32238
rect 6226 32182 6294 32238
rect 6350 32182 6418 32238
rect 6474 32182 6542 32238
rect 6598 32182 6666 32238
rect 6722 32182 6790 32238
rect 6846 32182 6914 32238
rect 6970 32182 7038 32238
rect 7094 32182 7104 32238
rect 5168 32114 7104 32182
rect 5168 32058 5178 32114
rect 5234 32058 5302 32114
rect 5358 32058 5426 32114
rect 5482 32058 5550 32114
rect 5606 32058 5674 32114
rect 5730 32058 5798 32114
rect 5854 32058 5922 32114
rect 5978 32058 6046 32114
rect 6102 32058 6170 32114
rect 6226 32058 6294 32114
rect 6350 32058 6418 32114
rect 6474 32058 6542 32114
rect 6598 32058 6666 32114
rect 6722 32058 6790 32114
rect 6846 32058 6914 32114
rect 6970 32058 7038 32114
rect 7094 32058 7104 32114
rect 5168 31990 7104 32058
rect 5168 31934 5178 31990
rect 5234 31934 5302 31990
rect 5358 31934 5426 31990
rect 5482 31934 5550 31990
rect 5606 31934 5674 31990
rect 5730 31934 5798 31990
rect 5854 31934 5922 31990
rect 5978 31934 6046 31990
rect 6102 31934 6170 31990
rect 6226 31934 6294 31990
rect 6350 31934 6418 31990
rect 6474 31934 6542 31990
rect 6598 31934 6666 31990
rect 6722 31934 6790 31990
rect 6846 31934 6914 31990
rect 6970 31934 7038 31990
rect 7094 31934 7104 31990
rect 5168 31866 7104 31934
rect 5168 31810 5178 31866
rect 5234 31810 5302 31866
rect 5358 31810 5426 31866
rect 5482 31810 5550 31866
rect 5606 31810 5674 31866
rect 5730 31810 5798 31866
rect 5854 31810 5922 31866
rect 5978 31810 6046 31866
rect 6102 31810 6170 31866
rect 6226 31810 6294 31866
rect 6350 31810 6418 31866
rect 6474 31810 6542 31866
rect 6598 31810 6666 31866
rect 6722 31810 6790 31866
rect 6846 31810 6914 31866
rect 6970 31810 7038 31866
rect 7094 31810 7104 31866
rect 5168 31742 7104 31810
rect 5168 31686 5178 31742
rect 5234 31686 5302 31742
rect 5358 31686 5426 31742
rect 5482 31686 5550 31742
rect 5606 31686 5674 31742
rect 5730 31686 5798 31742
rect 5854 31686 5922 31742
rect 5978 31686 6046 31742
rect 6102 31686 6170 31742
rect 6226 31686 6294 31742
rect 6350 31686 6418 31742
rect 6474 31686 6542 31742
rect 6598 31686 6666 31742
rect 6722 31686 6790 31742
rect 6846 31686 6914 31742
rect 6970 31686 7038 31742
rect 7094 31686 7104 31742
rect 5168 31618 7104 31686
rect 5168 31562 5178 31618
rect 5234 31562 5302 31618
rect 5358 31562 5426 31618
rect 5482 31562 5550 31618
rect 5606 31562 5674 31618
rect 5730 31562 5798 31618
rect 5854 31562 5922 31618
rect 5978 31562 6046 31618
rect 6102 31562 6170 31618
rect 6226 31562 6294 31618
rect 6350 31562 6418 31618
rect 6474 31562 6542 31618
rect 6598 31562 6666 31618
rect 6722 31562 6790 31618
rect 6846 31562 6914 31618
rect 6970 31562 7038 31618
rect 7094 31562 7104 31618
rect 5168 31494 7104 31562
rect 5168 31438 5178 31494
rect 5234 31438 5302 31494
rect 5358 31438 5426 31494
rect 5482 31438 5550 31494
rect 5606 31438 5674 31494
rect 5730 31438 5798 31494
rect 5854 31438 5922 31494
rect 5978 31438 6046 31494
rect 6102 31438 6170 31494
rect 6226 31438 6294 31494
rect 6350 31438 6418 31494
rect 6474 31438 6542 31494
rect 6598 31438 6666 31494
rect 6722 31438 6790 31494
rect 6846 31438 6914 31494
rect 6970 31438 7038 31494
rect 7094 31438 7104 31494
rect 5168 31370 7104 31438
rect 5168 31314 5178 31370
rect 5234 31314 5302 31370
rect 5358 31314 5426 31370
rect 5482 31314 5550 31370
rect 5606 31314 5674 31370
rect 5730 31314 5798 31370
rect 5854 31314 5922 31370
rect 5978 31314 6046 31370
rect 6102 31314 6170 31370
rect 6226 31314 6294 31370
rect 6350 31314 6418 31370
rect 6474 31314 6542 31370
rect 6598 31314 6666 31370
rect 6722 31314 6790 31370
rect 6846 31314 6914 31370
rect 6970 31314 7038 31370
rect 7094 31314 7104 31370
rect 5168 31246 7104 31314
rect 5168 31190 5178 31246
rect 5234 31190 5302 31246
rect 5358 31190 5426 31246
rect 5482 31190 5550 31246
rect 5606 31190 5674 31246
rect 5730 31190 5798 31246
rect 5854 31190 5922 31246
rect 5978 31190 6046 31246
rect 6102 31190 6170 31246
rect 6226 31190 6294 31246
rect 6350 31190 6418 31246
rect 6474 31190 6542 31246
rect 6598 31190 6666 31246
rect 6722 31190 6790 31246
rect 6846 31190 6914 31246
rect 6970 31190 7038 31246
rect 7094 31190 7104 31246
rect 5168 31122 7104 31190
rect 5168 31066 5178 31122
rect 5234 31066 5302 31122
rect 5358 31066 5426 31122
rect 5482 31066 5550 31122
rect 5606 31066 5674 31122
rect 5730 31066 5798 31122
rect 5854 31066 5922 31122
rect 5978 31066 6046 31122
rect 6102 31066 6170 31122
rect 6226 31066 6294 31122
rect 6350 31066 6418 31122
rect 6474 31066 6542 31122
rect 6598 31066 6666 31122
rect 6722 31066 6790 31122
rect 6846 31066 6914 31122
rect 6970 31066 7038 31122
rect 7094 31066 7104 31122
rect 5168 30998 7104 31066
rect 5168 30942 5178 30998
rect 5234 30942 5302 30998
rect 5358 30942 5426 30998
rect 5482 30942 5550 30998
rect 5606 30942 5674 30998
rect 5730 30942 5798 30998
rect 5854 30942 5922 30998
rect 5978 30942 6046 30998
rect 6102 30942 6170 30998
rect 6226 30942 6294 30998
rect 6350 30942 6418 30998
rect 6474 30942 6542 30998
rect 6598 30942 6666 30998
rect 6722 30942 6790 30998
rect 6846 30942 6914 30998
rect 6970 30942 7038 30998
rect 7094 30942 7104 30998
rect 5168 30874 7104 30942
rect 5168 30818 5178 30874
rect 5234 30818 5302 30874
rect 5358 30818 5426 30874
rect 5482 30818 5550 30874
rect 5606 30818 5674 30874
rect 5730 30818 5798 30874
rect 5854 30818 5922 30874
rect 5978 30818 6046 30874
rect 6102 30818 6170 30874
rect 6226 30818 6294 30874
rect 6350 30818 6418 30874
rect 6474 30818 6542 30874
rect 6598 30818 6666 30874
rect 6722 30818 6790 30874
rect 6846 30818 6914 30874
rect 6970 30818 7038 30874
rect 7094 30818 7104 30874
rect 5168 30750 7104 30818
rect 5168 30694 5178 30750
rect 5234 30694 5302 30750
rect 5358 30694 5426 30750
rect 5482 30694 5550 30750
rect 5606 30694 5674 30750
rect 5730 30694 5798 30750
rect 5854 30694 5922 30750
rect 5978 30694 6046 30750
rect 6102 30694 6170 30750
rect 6226 30694 6294 30750
rect 6350 30694 6418 30750
rect 6474 30694 6542 30750
rect 6598 30694 6666 30750
rect 6722 30694 6790 30750
rect 6846 30694 6914 30750
rect 6970 30694 7038 30750
rect 7094 30694 7104 30750
rect 5168 30626 7104 30694
rect 5168 30570 5178 30626
rect 5234 30570 5302 30626
rect 5358 30570 5426 30626
rect 5482 30570 5550 30626
rect 5606 30570 5674 30626
rect 5730 30570 5798 30626
rect 5854 30570 5922 30626
rect 5978 30570 6046 30626
rect 6102 30570 6170 30626
rect 6226 30570 6294 30626
rect 6350 30570 6418 30626
rect 6474 30570 6542 30626
rect 6598 30570 6666 30626
rect 6722 30570 6790 30626
rect 6846 30570 6914 30626
rect 6970 30570 7038 30626
rect 7094 30570 7104 30626
rect 5168 30502 7104 30570
rect 5168 30446 5178 30502
rect 5234 30446 5302 30502
rect 5358 30446 5426 30502
rect 5482 30446 5550 30502
rect 5606 30446 5674 30502
rect 5730 30446 5798 30502
rect 5854 30446 5922 30502
rect 5978 30446 6046 30502
rect 6102 30446 6170 30502
rect 6226 30446 6294 30502
rect 6350 30446 6418 30502
rect 6474 30446 6542 30502
rect 6598 30446 6666 30502
rect 6722 30446 6790 30502
rect 6846 30446 6914 30502
rect 6970 30446 7038 30502
rect 7094 30446 7104 30502
rect 5168 30436 7104 30446
rect 7874 33354 9810 33364
rect 7874 33298 7884 33354
rect 7940 33298 8008 33354
rect 8064 33298 8132 33354
rect 8188 33298 8256 33354
rect 8312 33298 8380 33354
rect 8436 33298 8504 33354
rect 8560 33298 8628 33354
rect 8684 33298 8752 33354
rect 8808 33298 8876 33354
rect 8932 33298 9000 33354
rect 9056 33298 9124 33354
rect 9180 33298 9248 33354
rect 9304 33298 9372 33354
rect 9428 33298 9496 33354
rect 9552 33298 9620 33354
rect 9676 33298 9744 33354
rect 9800 33298 9810 33354
rect 7874 33230 9810 33298
rect 7874 33174 7884 33230
rect 7940 33174 8008 33230
rect 8064 33174 8132 33230
rect 8188 33174 8256 33230
rect 8312 33174 8380 33230
rect 8436 33174 8504 33230
rect 8560 33174 8628 33230
rect 8684 33174 8752 33230
rect 8808 33174 8876 33230
rect 8932 33174 9000 33230
rect 9056 33174 9124 33230
rect 9180 33174 9248 33230
rect 9304 33174 9372 33230
rect 9428 33174 9496 33230
rect 9552 33174 9620 33230
rect 9676 33174 9744 33230
rect 9800 33174 9810 33230
rect 7874 33106 9810 33174
rect 7874 33050 7884 33106
rect 7940 33050 8008 33106
rect 8064 33050 8132 33106
rect 8188 33050 8256 33106
rect 8312 33050 8380 33106
rect 8436 33050 8504 33106
rect 8560 33050 8628 33106
rect 8684 33050 8752 33106
rect 8808 33050 8876 33106
rect 8932 33050 9000 33106
rect 9056 33050 9124 33106
rect 9180 33050 9248 33106
rect 9304 33050 9372 33106
rect 9428 33050 9496 33106
rect 9552 33050 9620 33106
rect 9676 33050 9744 33106
rect 9800 33050 9810 33106
rect 7874 32982 9810 33050
rect 7874 32926 7884 32982
rect 7940 32926 8008 32982
rect 8064 32926 8132 32982
rect 8188 32926 8256 32982
rect 8312 32926 8380 32982
rect 8436 32926 8504 32982
rect 8560 32926 8628 32982
rect 8684 32926 8752 32982
rect 8808 32926 8876 32982
rect 8932 32926 9000 32982
rect 9056 32926 9124 32982
rect 9180 32926 9248 32982
rect 9304 32926 9372 32982
rect 9428 32926 9496 32982
rect 9552 32926 9620 32982
rect 9676 32926 9744 32982
rect 9800 32926 9810 32982
rect 7874 32858 9810 32926
rect 7874 32802 7884 32858
rect 7940 32802 8008 32858
rect 8064 32802 8132 32858
rect 8188 32802 8256 32858
rect 8312 32802 8380 32858
rect 8436 32802 8504 32858
rect 8560 32802 8628 32858
rect 8684 32802 8752 32858
rect 8808 32802 8876 32858
rect 8932 32802 9000 32858
rect 9056 32802 9124 32858
rect 9180 32802 9248 32858
rect 9304 32802 9372 32858
rect 9428 32802 9496 32858
rect 9552 32802 9620 32858
rect 9676 32802 9744 32858
rect 9800 32802 9810 32858
rect 7874 32734 9810 32802
rect 7874 32678 7884 32734
rect 7940 32678 8008 32734
rect 8064 32678 8132 32734
rect 8188 32678 8256 32734
rect 8312 32678 8380 32734
rect 8436 32678 8504 32734
rect 8560 32678 8628 32734
rect 8684 32678 8752 32734
rect 8808 32678 8876 32734
rect 8932 32678 9000 32734
rect 9056 32678 9124 32734
rect 9180 32678 9248 32734
rect 9304 32678 9372 32734
rect 9428 32678 9496 32734
rect 9552 32678 9620 32734
rect 9676 32678 9744 32734
rect 9800 32678 9810 32734
rect 7874 32610 9810 32678
rect 7874 32554 7884 32610
rect 7940 32554 8008 32610
rect 8064 32554 8132 32610
rect 8188 32554 8256 32610
rect 8312 32554 8380 32610
rect 8436 32554 8504 32610
rect 8560 32554 8628 32610
rect 8684 32554 8752 32610
rect 8808 32554 8876 32610
rect 8932 32554 9000 32610
rect 9056 32554 9124 32610
rect 9180 32554 9248 32610
rect 9304 32554 9372 32610
rect 9428 32554 9496 32610
rect 9552 32554 9620 32610
rect 9676 32554 9744 32610
rect 9800 32554 9810 32610
rect 7874 32486 9810 32554
rect 7874 32430 7884 32486
rect 7940 32430 8008 32486
rect 8064 32430 8132 32486
rect 8188 32430 8256 32486
rect 8312 32430 8380 32486
rect 8436 32430 8504 32486
rect 8560 32430 8628 32486
rect 8684 32430 8752 32486
rect 8808 32430 8876 32486
rect 8932 32430 9000 32486
rect 9056 32430 9124 32486
rect 9180 32430 9248 32486
rect 9304 32430 9372 32486
rect 9428 32430 9496 32486
rect 9552 32430 9620 32486
rect 9676 32430 9744 32486
rect 9800 32430 9810 32486
rect 7874 32362 9810 32430
rect 7874 32306 7884 32362
rect 7940 32306 8008 32362
rect 8064 32306 8132 32362
rect 8188 32306 8256 32362
rect 8312 32306 8380 32362
rect 8436 32306 8504 32362
rect 8560 32306 8628 32362
rect 8684 32306 8752 32362
rect 8808 32306 8876 32362
rect 8932 32306 9000 32362
rect 9056 32306 9124 32362
rect 9180 32306 9248 32362
rect 9304 32306 9372 32362
rect 9428 32306 9496 32362
rect 9552 32306 9620 32362
rect 9676 32306 9744 32362
rect 9800 32306 9810 32362
rect 7874 32238 9810 32306
rect 7874 32182 7884 32238
rect 7940 32182 8008 32238
rect 8064 32182 8132 32238
rect 8188 32182 8256 32238
rect 8312 32182 8380 32238
rect 8436 32182 8504 32238
rect 8560 32182 8628 32238
rect 8684 32182 8752 32238
rect 8808 32182 8876 32238
rect 8932 32182 9000 32238
rect 9056 32182 9124 32238
rect 9180 32182 9248 32238
rect 9304 32182 9372 32238
rect 9428 32182 9496 32238
rect 9552 32182 9620 32238
rect 9676 32182 9744 32238
rect 9800 32182 9810 32238
rect 7874 32114 9810 32182
rect 7874 32058 7884 32114
rect 7940 32058 8008 32114
rect 8064 32058 8132 32114
rect 8188 32058 8256 32114
rect 8312 32058 8380 32114
rect 8436 32058 8504 32114
rect 8560 32058 8628 32114
rect 8684 32058 8752 32114
rect 8808 32058 8876 32114
rect 8932 32058 9000 32114
rect 9056 32058 9124 32114
rect 9180 32058 9248 32114
rect 9304 32058 9372 32114
rect 9428 32058 9496 32114
rect 9552 32058 9620 32114
rect 9676 32058 9744 32114
rect 9800 32058 9810 32114
rect 7874 31990 9810 32058
rect 7874 31934 7884 31990
rect 7940 31934 8008 31990
rect 8064 31934 8132 31990
rect 8188 31934 8256 31990
rect 8312 31934 8380 31990
rect 8436 31934 8504 31990
rect 8560 31934 8628 31990
rect 8684 31934 8752 31990
rect 8808 31934 8876 31990
rect 8932 31934 9000 31990
rect 9056 31934 9124 31990
rect 9180 31934 9248 31990
rect 9304 31934 9372 31990
rect 9428 31934 9496 31990
rect 9552 31934 9620 31990
rect 9676 31934 9744 31990
rect 9800 31934 9810 31990
rect 7874 31866 9810 31934
rect 7874 31810 7884 31866
rect 7940 31810 8008 31866
rect 8064 31810 8132 31866
rect 8188 31810 8256 31866
rect 8312 31810 8380 31866
rect 8436 31810 8504 31866
rect 8560 31810 8628 31866
rect 8684 31810 8752 31866
rect 8808 31810 8876 31866
rect 8932 31810 9000 31866
rect 9056 31810 9124 31866
rect 9180 31810 9248 31866
rect 9304 31810 9372 31866
rect 9428 31810 9496 31866
rect 9552 31810 9620 31866
rect 9676 31810 9744 31866
rect 9800 31810 9810 31866
rect 7874 31742 9810 31810
rect 7874 31686 7884 31742
rect 7940 31686 8008 31742
rect 8064 31686 8132 31742
rect 8188 31686 8256 31742
rect 8312 31686 8380 31742
rect 8436 31686 8504 31742
rect 8560 31686 8628 31742
rect 8684 31686 8752 31742
rect 8808 31686 8876 31742
rect 8932 31686 9000 31742
rect 9056 31686 9124 31742
rect 9180 31686 9248 31742
rect 9304 31686 9372 31742
rect 9428 31686 9496 31742
rect 9552 31686 9620 31742
rect 9676 31686 9744 31742
rect 9800 31686 9810 31742
rect 7874 31618 9810 31686
rect 7874 31562 7884 31618
rect 7940 31562 8008 31618
rect 8064 31562 8132 31618
rect 8188 31562 8256 31618
rect 8312 31562 8380 31618
rect 8436 31562 8504 31618
rect 8560 31562 8628 31618
rect 8684 31562 8752 31618
rect 8808 31562 8876 31618
rect 8932 31562 9000 31618
rect 9056 31562 9124 31618
rect 9180 31562 9248 31618
rect 9304 31562 9372 31618
rect 9428 31562 9496 31618
rect 9552 31562 9620 31618
rect 9676 31562 9744 31618
rect 9800 31562 9810 31618
rect 7874 31494 9810 31562
rect 7874 31438 7884 31494
rect 7940 31438 8008 31494
rect 8064 31438 8132 31494
rect 8188 31438 8256 31494
rect 8312 31438 8380 31494
rect 8436 31438 8504 31494
rect 8560 31438 8628 31494
rect 8684 31438 8752 31494
rect 8808 31438 8876 31494
rect 8932 31438 9000 31494
rect 9056 31438 9124 31494
rect 9180 31438 9248 31494
rect 9304 31438 9372 31494
rect 9428 31438 9496 31494
rect 9552 31438 9620 31494
rect 9676 31438 9744 31494
rect 9800 31438 9810 31494
rect 7874 31370 9810 31438
rect 7874 31314 7884 31370
rect 7940 31314 8008 31370
rect 8064 31314 8132 31370
rect 8188 31314 8256 31370
rect 8312 31314 8380 31370
rect 8436 31314 8504 31370
rect 8560 31314 8628 31370
rect 8684 31314 8752 31370
rect 8808 31314 8876 31370
rect 8932 31314 9000 31370
rect 9056 31314 9124 31370
rect 9180 31314 9248 31370
rect 9304 31314 9372 31370
rect 9428 31314 9496 31370
rect 9552 31314 9620 31370
rect 9676 31314 9744 31370
rect 9800 31314 9810 31370
rect 7874 31246 9810 31314
rect 7874 31190 7884 31246
rect 7940 31190 8008 31246
rect 8064 31190 8132 31246
rect 8188 31190 8256 31246
rect 8312 31190 8380 31246
rect 8436 31190 8504 31246
rect 8560 31190 8628 31246
rect 8684 31190 8752 31246
rect 8808 31190 8876 31246
rect 8932 31190 9000 31246
rect 9056 31190 9124 31246
rect 9180 31190 9248 31246
rect 9304 31190 9372 31246
rect 9428 31190 9496 31246
rect 9552 31190 9620 31246
rect 9676 31190 9744 31246
rect 9800 31190 9810 31246
rect 7874 31122 9810 31190
rect 7874 31066 7884 31122
rect 7940 31066 8008 31122
rect 8064 31066 8132 31122
rect 8188 31066 8256 31122
rect 8312 31066 8380 31122
rect 8436 31066 8504 31122
rect 8560 31066 8628 31122
rect 8684 31066 8752 31122
rect 8808 31066 8876 31122
rect 8932 31066 9000 31122
rect 9056 31066 9124 31122
rect 9180 31066 9248 31122
rect 9304 31066 9372 31122
rect 9428 31066 9496 31122
rect 9552 31066 9620 31122
rect 9676 31066 9744 31122
rect 9800 31066 9810 31122
rect 7874 30998 9810 31066
rect 7874 30942 7884 30998
rect 7940 30942 8008 30998
rect 8064 30942 8132 30998
rect 8188 30942 8256 30998
rect 8312 30942 8380 30998
rect 8436 30942 8504 30998
rect 8560 30942 8628 30998
rect 8684 30942 8752 30998
rect 8808 30942 8876 30998
rect 8932 30942 9000 30998
rect 9056 30942 9124 30998
rect 9180 30942 9248 30998
rect 9304 30942 9372 30998
rect 9428 30942 9496 30998
rect 9552 30942 9620 30998
rect 9676 30942 9744 30998
rect 9800 30942 9810 30998
rect 7874 30874 9810 30942
rect 7874 30818 7884 30874
rect 7940 30818 8008 30874
rect 8064 30818 8132 30874
rect 8188 30818 8256 30874
rect 8312 30818 8380 30874
rect 8436 30818 8504 30874
rect 8560 30818 8628 30874
rect 8684 30818 8752 30874
rect 8808 30818 8876 30874
rect 8932 30818 9000 30874
rect 9056 30818 9124 30874
rect 9180 30818 9248 30874
rect 9304 30818 9372 30874
rect 9428 30818 9496 30874
rect 9552 30818 9620 30874
rect 9676 30818 9744 30874
rect 9800 30818 9810 30874
rect 7874 30750 9810 30818
rect 7874 30694 7884 30750
rect 7940 30694 8008 30750
rect 8064 30694 8132 30750
rect 8188 30694 8256 30750
rect 8312 30694 8380 30750
rect 8436 30694 8504 30750
rect 8560 30694 8628 30750
rect 8684 30694 8752 30750
rect 8808 30694 8876 30750
rect 8932 30694 9000 30750
rect 9056 30694 9124 30750
rect 9180 30694 9248 30750
rect 9304 30694 9372 30750
rect 9428 30694 9496 30750
rect 9552 30694 9620 30750
rect 9676 30694 9744 30750
rect 9800 30694 9810 30750
rect 7874 30626 9810 30694
rect 7874 30570 7884 30626
rect 7940 30570 8008 30626
rect 8064 30570 8132 30626
rect 8188 30570 8256 30626
rect 8312 30570 8380 30626
rect 8436 30570 8504 30626
rect 8560 30570 8628 30626
rect 8684 30570 8752 30626
rect 8808 30570 8876 30626
rect 8932 30570 9000 30626
rect 9056 30570 9124 30626
rect 9180 30570 9248 30626
rect 9304 30570 9372 30626
rect 9428 30570 9496 30626
rect 9552 30570 9620 30626
rect 9676 30570 9744 30626
rect 9800 30570 9810 30626
rect 7874 30502 9810 30570
rect 7874 30446 7884 30502
rect 7940 30446 8008 30502
rect 8064 30446 8132 30502
rect 8188 30446 8256 30502
rect 8312 30446 8380 30502
rect 8436 30446 8504 30502
rect 8560 30446 8628 30502
rect 8684 30446 8752 30502
rect 8808 30446 8876 30502
rect 8932 30446 9000 30502
rect 9056 30446 9124 30502
rect 9180 30446 9248 30502
rect 9304 30446 9372 30502
rect 9428 30446 9496 30502
rect 9552 30446 9620 30502
rect 9676 30446 9744 30502
rect 9800 30446 9810 30502
rect 7874 30436 9810 30446
rect 10244 33354 12180 33364
rect 10244 33298 10254 33354
rect 10310 33298 10378 33354
rect 10434 33298 10502 33354
rect 10558 33298 10626 33354
rect 10682 33298 10750 33354
rect 10806 33298 10874 33354
rect 10930 33298 10998 33354
rect 11054 33298 11122 33354
rect 11178 33298 11246 33354
rect 11302 33298 11370 33354
rect 11426 33298 11494 33354
rect 11550 33298 11618 33354
rect 11674 33298 11742 33354
rect 11798 33298 11866 33354
rect 11922 33298 11990 33354
rect 12046 33298 12114 33354
rect 12170 33298 12180 33354
rect 10244 33230 12180 33298
rect 10244 33174 10254 33230
rect 10310 33174 10378 33230
rect 10434 33174 10502 33230
rect 10558 33174 10626 33230
rect 10682 33174 10750 33230
rect 10806 33174 10874 33230
rect 10930 33174 10998 33230
rect 11054 33174 11122 33230
rect 11178 33174 11246 33230
rect 11302 33174 11370 33230
rect 11426 33174 11494 33230
rect 11550 33174 11618 33230
rect 11674 33174 11742 33230
rect 11798 33174 11866 33230
rect 11922 33174 11990 33230
rect 12046 33174 12114 33230
rect 12170 33174 12180 33230
rect 10244 33106 12180 33174
rect 10244 33050 10254 33106
rect 10310 33050 10378 33106
rect 10434 33050 10502 33106
rect 10558 33050 10626 33106
rect 10682 33050 10750 33106
rect 10806 33050 10874 33106
rect 10930 33050 10998 33106
rect 11054 33050 11122 33106
rect 11178 33050 11246 33106
rect 11302 33050 11370 33106
rect 11426 33050 11494 33106
rect 11550 33050 11618 33106
rect 11674 33050 11742 33106
rect 11798 33050 11866 33106
rect 11922 33050 11990 33106
rect 12046 33050 12114 33106
rect 12170 33050 12180 33106
rect 10244 32982 12180 33050
rect 10244 32926 10254 32982
rect 10310 32926 10378 32982
rect 10434 32926 10502 32982
rect 10558 32926 10626 32982
rect 10682 32926 10750 32982
rect 10806 32926 10874 32982
rect 10930 32926 10998 32982
rect 11054 32926 11122 32982
rect 11178 32926 11246 32982
rect 11302 32926 11370 32982
rect 11426 32926 11494 32982
rect 11550 32926 11618 32982
rect 11674 32926 11742 32982
rect 11798 32926 11866 32982
rect 11922 32926 11990 32982
rect 12046 32926 12114 32982
rect 12170 32926 12180 32982
rect 10244 32858 12180 32926
rect 10244 32802 10254 32858
rect 10310 32802 10378 32858
rect 10434 32802 10502 32858
rect 10558 32802 10626 32858
rect 10682 32802 10750 32858
rect 10806 32802 10874 32858
rect 10930 32802 10998 32858
rect 11054 32802 11122 32858
rect 11178 32802 11246 32858
rect 11302 32802 11370 32858
rect 11426 32802 11494 32858
rect 11550 32802 11618 32858
rect 11674 32802 11742 32858
rect 11798 32802 11866 32858
rect 11922 32802 11990 32858
rect 12046 32802 12114 32858
rect 12170 32802 12180 32858
rect 10244 32734 12180 32802
rect 10244 32678 10254 32734
rect 10310 32678 10378 32734
rect 10434 32678 10502 32734
rect 10558 32678 10626 32734
rect 10682 32678 10750 32734
rect 10806 32678 10874 32734
rect 10930 32678 10998 32734
rect 11054 32678 11122 32734
rect 11178 32678 11246 32734
rect 11302 32678 11370 32734
rect 11426 32678 11494 32734
rect 11550 32678 11618 32734
rect 11674 32678 11742 32734
rect 11798 32678 11866 32734
rect 11922 32678 11990 32734
rect 12046 32678 12114 32734
rect 12170 32678 12180 32734
rect 10244 32610 12180 32678
rect 10244 32554 10254 32610
rect 10310 32554 10378 32610
rect 10434 32554 10502 32610
rect 10558 32554 10626 32610
rect 10682 32554 10750 32610
rect 10806 32554 10874 32610
rect 10930 32554 10998 32610
rect 11054 32554 11122 32610
rect 11178 32554 11246 32610
rect 11302 32554 11370 32610
rect 11426 32554 11494 32610
rect 11550 32554 11618 32610
rect 11674 32554 11742 32610
rect 11798 32554 11866 32610
rect 11922 32554 11990 32610
rect 12046 32554 12114 32610
rect 12170 32554 12180 32610
rect 10244 32486 12180 32554
rect 10244 32430 10254 32486
rect 10310 32430 10378 32486
rect 10434 32430 10502 32486
rect 10558 32430 10626 32486
rect 10682 32430 10750 32486
rect 10806 32430 10874 32486
rect 10930 32430 10998 32486
rect 11054 32430 11122 32486
rect 11178 32430 11246 32486
rect 11302 32430 11370 32486
rect 11426 32430 11494 32486
rect 11550 32430 11618 32486
rect 11674 32430 11742 32486
rect 11798 32430 11866 32486
rect 11922 32430 11990 32486
rect 12046 32430 12114 32486
rect 12170 32430 12180 32486
rect 10244 32362 12180 32430
rect 10244 32306 10254 32362
rect 10310 32306 10378 32362
rect 10434 32306 10502 32362
rect 10558 32306 10626 32362
rect 10682 32306 10750 32362
rect 10806 32306 10874 32362
rect 10930 32306 10998 32362
rect 11054 32306 11122 32362
rect 11178 32306 11246 32362
rect 11302 32306 11370 32362
rect 11426 32306 11494 32362
rect 11550 32306 11618 32362
rect 11674 32306 11742 32362
rect 11798 32306 11866 32362
rect 11922 32306 11990 32362
rect 12046 32306 12114 32362
rect 12170 32306 12180 32362
rect 10244 32238 12180 32306
rect 10244 32182 10254 32238
rect 10310 32182 10378 32238
rect 10434 32182 10502 32238
rect 10558 32182 10626 32238
rect 10682 32182 10750 32238
rect 10806 32182 10874 32238
rect 10930 32182 10998 32238
rect 11054 32182 11122 32238
rect 11178 32182 11246 32238
rect 11302 32182 11370 32238
rect 11426 32182 11494 32238
rect 11550 32182 11618 32238
rect 11674 32182 11742 32238
rect 11798 32182 11866 32238
rect 11922 32182 11990 32238
rect 12046 32182 12114 32238
rect 12170 32182 12180 32238
rect 10244 32114 12180 32182
rect 10244 32058 10254 32114
rect 10310 32058 10378 32114
rect 10434 32058 10502 32114
rect 10558 32058 10626 32114
rect 10682 32058 10750 32114
rect 10806 32058 10874 32114
rect 10930 32058 10998 32114
rect 11054 32058 11122 32114
rect 11178 32058 11246 32114
rect 11302 32058 11370 32114
rect 11426 32058 11494 32114
rect 11550 32058 11618 32114
rect 11674 32058 11742 32114
rect 11798 32058 11866 32114
rect 11922 32058 11990 32114
rect 12046 32058 12114 32114
rect 12170 32058 12180 32114
rect 10244 31990 12180 32058
rect 10244 31934 10254 31990
rect 10310 31934 10378 31990
rect 10434 31934 10502 31990
rect 10558 31934 10626 31990
rect 10682 31934 10750 31990
rect 10806 31934 10874 31990
rect 10930 31934 10998 31990
rect 11054 31934 11122 31990
rect 11178 31934 11246 31990
rect 11302 31934 11370 31990
rect 11426 31934 11494 31990
rect 11550 31934 11618 31990
rect 11674 31934 11742 31990
rect 11798 31934 11866 31990
rect 11922 31934 11990 31990
rect 12046 31934 12114 31990
rect 12170 31934 12180 31990
rect 10244 31866 12180 31934
rect 10244 31810 10254 31866
rect 10310 31810 10378 31866
rect 10434 31810 10502 31866
rect 10558 31810 10626 31866
rect 10682 31810 10750 31866
rect 10806 31810 10874 31866
rect 10930 31810 10998 31866
rect 11054 31810 11122 31866
rect 11178 31810 11246 31866
rect 11302 31810 11370 31866
rect 11426 31810 11494 31866
rect 11550 31810 11618 31866
rect 11674 31810 11742 31866
rect 11798 31810 11866 31866
rect 11922 31810 11990 31866
rect 12046 31810 12114 31866
rect 12170 31810 12180 31866
rect 10244 31742 12180 31810
rect 10244 31686 10254 31742
rect 10310 31686 10378 31742
rect 10434 31686 10502 31742
rect 10558 31686 10626 31742
rect 10682 31686 10750 31742
rect 10806 31686 10874 31742
rect 10930 31686 10998 31742
rect 11054 31686 11122 31742
rect 11178 31686 11246 31742
rect 11302 31686 11370 31742
rect 11426 31686 11494 31742
rect 11550 31686 11618 31742
rect 11674 31686 11742 31742
rect 11798 31686 11866 31742
rect 11922 31686 11990 31742
rect 12046 31686 12114 31742
rect 12170 31686 12180 31742
rect 10244 31618 12180 31686
rect 10244 31562 10254 31618
rect 10310 31562 10378 31618
rect 10434 31562 10502 31618
rect 10558 31562 10626 31618
rect 10682 31562 10750 31618
rect 10806 31562 10874 31618
rect 10930 31562 10998 31618
rect 11054 31562 11122 31618
rect 11178 31562 11246 31618
rect 11302 31562 11370 31618
rect 11426 31562 11494 31618
rect 11550 31562 11618 31618
rect 11674 31562 11742 31618
rect 11798 31562 11866 31618
rect 11922 31562 11990 31618
rect 12046 31562 12114 31618
rect 12170 31562 12180 31618
rect 10244 31494 12180 31562
rect 10244 31438 10254 31494
rect 10310 31438 10378 31494
rect 10434 31438 10502 31494
rect 10558 31438 10626 31494
rect 10682 31438 10750 31494
rect 10806 31438 10874 31494
rect 10930 31438 10998 31494
rect 11054 31438 11122 31494
rect 11178 31438 11246 31494
rect 11302 31438 11370 31494
rect 11426 31438 11494 31494
rect 11550 31438 11618 31494
rect 11674 31438 11742 31494
rect 11798 31438 11866 31494
rect 11922 31438 11990 31494
rect 12046 31438 12114 31494
rect 12170 31438 12180 31494
rect 10244 31370 12180 31438
rect 10244 31314 10254 31370
rect 10310 31314 10378 31370
rect 10434 31314 10502 31370
rect 10558 31314 10626 31370
rect 10682 31314 10750 31370
rect 10806 31314 10874 31370
rect 10930 31314 10998 31370
rect 11054 31314 11122 31370
rect 11178 31314 11246 31370
rect 11302 31314 11370 31370
rect 11426 31314 11494 31370
rect 11550 31314 11618 31370
rect 11674 31314 11742 31370
rect 11798 31314 11866 31370
rect 11922 31314 11990 31370
rect 12046 31314 12114 31370
rect 12170 31314 12180 31370
rect 10244 31246 12180 31314
rect 10244 31190 10254 31246
rect 10310 31190 10378 31246
rect 10434 31190 10502 31246
rect 10558 31190 10626 31246
rect 10682 31190 10750 31246
rect 10806 31190 10874 31246
rect 10930 31190 10998 31246
rect 11054 31190 11122 31246
rect 11178 31190 11246 31246
rect 11302 31190 11370 31246
rect 11426 31190 11494 31246
rect 11550 31190 11618 31246
rect 11674 31190 11742 31246
rect 11798 31190 11866 31246
rect 11922 31190 11990 31246
rect 12046 31190 12114 31246
rect 12170 31190 12180 31246
rect 10244 31122 12180 31190
rect 10244 31066 10254 31122
rect 10310 31066 10378 31122
rect 10434 31066 10502 31122
rect 10558 31066 10626 31122
rect 10682 31066 10750 31122
rect 10806 31066 10874 31122
rect 10930 31066 10998 31122
rect 11054 31066 11122 31122
rect 11178 31066 11246 31122
rect 11302 31066 11370 31122
rect 11426 31066 11494 31122
rect 11550 31066 11618 31122
rect 11674 31066 11742 31122
rect 11798 31066 11866 31122
rect 11922 31066 11990 31122
rect 12046 31066 12114 31122
rect 12170 31066 12180 31122
rect 10244 30998 12180 31066
rect 10244 30942 10254 30998
rect 10310 30942 10378 30998
rect 10434 30942 10502 30998
rect 10558 30942 10626 30998
rect 10682 30942 10750 30998
rect 10806 30942 10874 30998
rect 10930 30942 10998 30998
rect 11054 30942 11122 30998
rect 11178 30942 11246 30998
rect 11302 30942 11370 30998
rect 11426 30942 11494 30998
rect 11550 30942 11618 30998
rect 11674 30942 11742 30998
rect 11798 30942 11866 30998
rect 11922 30942 11990 30998
rect 12046 30942 12114 30998
rect 12170 30942 12180 30998
rect 10244 30874 12180 30942
rect 10244 30818 10254 30874
rect 10310 30818 10378 30874
rect 10434 30818 10502 30874
rect 10558 30818 10626 30874
rect 10682 30818 10750 30874
rect 10806 30818 10874 30874
rect 10930 30818 10998 30874
rect 11054 30818 11122 30874
rect 11178 30818 11246 30874
rect 11302 30818 11370 30874
rect 11426 30818 11494 30874
rect 11550 30818 11618 30874
rect 11674 30818 11742 30874
rect 11798 30818 11866 30874
rect 11922 30818 11990 30874
rect 12046 30818 12114 30874
rect 12170 30818 12180 30874
rect 10244 30750 12180 30818
rect 10244 30694 10254 30750
rect 10310 30694 10378 30750
rect 10434 30694 10502 30750
rect 10558 30694 10626 30750
rect 10682 30694 10750 30750
rect 10806 30694 10874 30750
rect 10930 30694 10998 30750
rect 11054 30694 11122 30750
rect 11178 30694 11246 30750
rect 11302 30694 11370 30750
rect 11426 30694 11494 30750
rect 11550 30694 11618 30750
rect 11674 30694 11742 30750
rect 11798 30694 11866 30750
rect 11922 30694 11990 30750
rect 12046 30694 12114 30750
rect 12170 30694 12180 30750
rect 10244 30626 12180 30694
rect 10244 30570 10254 30626
rect 10310 30570 10378 30626
rect 10434 30570 10502 30626
rect 10558 30570 10626 30626
rect 10682 30570 10750 30626
rect 10806 30570 10874 30626
rect 10930 30570 10998 30626
rect 11054 30570 11122 30626
rect 11178 30570 11246 30626
rect 11302 30570 11370 30626
rect 11426 30570 11494 30626
rect 11550 30570 11618 30626
rect 11674 30570 11742 30626
rect 11798 30570 11866 30626
rect 11922 30570 11990 30626
rect 12046 30570 12114 30626
rect 12170 30570 12180 30626
rect 10244 30502 12180 30570
rect 10244 30446 10254 30502
rect 10310 30446 10378 30502
rect 10434 30446 10502 30502
rect 10558 30446 10626 30502
rect 10682 30446 10750 30502
rect 10806 30446 10874 30502
rect 10930 30446 10998 30502
rect 11054 30446 11122 30502
rect 11178 30446 11246 30502
rect 11302 30446 11370 30502
rect 11426 30446 11494 30502
rect 11550 30446 11618 30502
rect 11674 30446 11742 30502
rect 11798 30446 11866 30502
rect 11922 30446 11990 30502
rect 12046 30446 12114 30502
rect 12170 30446 12180 30502
rect 10244 30436 12180 30446
rect 12861 33354 14673 33364
rect 12861 33298 12871 33354
rect 12927 33298 12995 33354
rect 13051 33298 13119 33354
rect 13175 33298 13243 33354
rect 13299 33298 13367 33354
rect 13423 33298 13491 33354
rect 13547 33298 13615 33354
rect 13671 33298 13739 33354
rect 13795 33298 13863 33354
rect 13919 33298 13987 33354
rect 14043 33298 14111 33354
rect 14167 33298 14235 33354
rect 14291 33298 14359 33354
rect 14415 33298 14483 33354
rect 14539 33298 14607 33354
rect 14663 33298 14673 33354
rect 12861 33230 14673 33298
rect 12861 33174 12871 33230
rect 12927 33174 12995 33230
rect 13051 33174 13119 33230
rect 13175 33174 13243 33230
rect 13299 33174 13367 33230
rect 13423 33174 13491 33230
rect 13547 33174 13615 33230
rect 13671 33174 13739 33230
rect 13795 33174 13863 33230
rect 13919 33174 13987 33230
rect 14043 33174 14111 33230
rect 14167 33174 14235 33230
rect 14291 33174 14359 33230
rect 14415 33174 14483 33230
rect 14539 33174 14607 33230
rect 14663 33174 14673 33230
rect 12861 33106 14673 33174
rect 12861 33050 12871 33106
rect 12927 33050 12995 33106
rect 13051 33050 13119 33106
rect 13175 33050 13243 33106
rect 13299 33050 13367 33106
rect 13423 33050 13491 33106
rect 13547 33050 13615 33106
rect 13671 33050 13739 33106
rect 13795 33050 13863 33106
rect 13919 33050 13987 33106
rect 14043 33050 14111 33106
rect 14167 33050 14235 33106
rect 14291 33050 14359 33106
rect 14415 33050 14483 33106
rect 14539 33050 14607 33106
rect 14663 33050 14673 33106
rect 12861 32982 14673 33050
rect 12861 32926 12871 32982
rect 12927 32926 12995 32982
rect 13051 32926 13119 32982
rect 13175 32926 13243 32982
rect 13299 32926 13367 32982
rect 13423 32926 13491 32982
rect 13547 32926 13615 32982
rect 13671 32926 13739 32982
rect 13795 32926 13863 32982
rect 13919 32926 13987 32982
rect 14043 32926 14111 32982
rect 14167 32926 14235 32982
rect 14291 32926 14359 32982
rect 14415 32926 14483 32982
rect 14539 32926 14607 32982
rect 14663 32926 14673 32982
rect 12861 32858 14673 32926
rect 12861 32802 12871 32858
rect 12927 32802 12995 32858
rect 13051 32802 13119 32858
rect 13175 32802 13243 32858
rect 13299 32802 13367 32858
rect 13423 32802 13491 32858
rect 13547 32802 13615 32858
rect 13671 32802 13739 32858
rect 13795 32802 13863 32858
rect 13919 32802 13987 32858
rect 14043 32802 14111 32858
rect 14167 32802 14235 32858
rect 14291 32802 14359 32858
rect 14415 32802 14483 32858
rect 14539 32802 14607 32858
rect 14663 32802 14673 32858
rect 12861 32734 14673 32802
rect 12861 32678 12871 32734
rect 12927 32678 12995 32734
rect 13051 32678 13119 32734
rect 13175 32678 13243 32734
rect 13299 32678 13367 32734
rect 13423 32678 13491 32734
rect 13547 32678 13615 32734
rect 13671 32678 13739 32734
rect 13795 32678 13863 32734
rect 13919 32678 13987 32734
rect 14043 32678 14111 32734
rect 14167 32678 14235 32734
rect 14291 32678 14359 32734
rect 14415 32678 14483 32734
rect 14539 32678 14607 32734
rect 14663 32678 14673 32734
rect 12861 32610 14673 32678
rect 12861 32554 12871 32610
rect 12927 32554 12995 32610
rect 13051 32554 13119 32610
rect 13175 32554 13243 32610
rect 13299 32554 13367 32610
rect 13423 32554 13491 32610
rect 13547 32554 13615 32610
rect 13671 32554 13739 32610
rect 13795 32554 13863 32610
rect 13919 32554 13987 32610
rect 14043 32554 14111 32610
rect 14167 32554 14235 32610
rect 14291 32554 14359 32610
rect 14415 32554 14483 32610
rect 14539 32554 14607 32610
rect 14663 32554 14673 32610
rect 12861 32486 14673 32554
rect 12861 32430 12871 32486
rect 12927 32430 12995 32486
rect 13051 32430 13119 32486
rect 13175 32430 13243 32486
rect 13299 32430 13367 32486
rect 13423 32430 13491 32486
rect 13547 32430 13615 32486
rect 13671 32430 13739 32486
rect 13795 32430 13863 32486
rect 13919 32430 13987 32486
rect 14043 32430 14111 32486
rect 14167 32430 14235 32486
rect 14291 32430 14359 32486
rect 14415 32430 14483 32486
rect 14539 32430 14607 32486
rect 14663 32430 14673 32486
rect 12861 32362 14673 32430
rect 12861 32306 12871 32362
rect 12927 32306 12995 32362
rect 13051 32306 13119 32362
rect 13175 32306 13243 32362
rect 13299 32306 13367 32362
rect 13423 32306 13491 32362
rect 13547 32306 13615 32362
rect 13671 32306 13739 32362
rect 13795 32306 13863 32362
rect 13919 32306 13987 32362
rect 14043 32306 14111 32362
rect 14167 32306 14235 32362
rect 14291 32306 14359 32362
rect 14415 32306 14483 32362
rect 14539 32306 14607 32362
rect 14663 32306 14673 32362
rect 12861 32238 14673 32306
rect 12861 32182 12871 32238
rect 12927 32182 12995 32238
rect 13051 32182 13119 32238
rect 13175 32182 13243 32238
rect 13299 32182 13367 32238
rect 13423 32182 13491 32238
rect 13547 32182 13615 32238
rect 13671 32182 13739 32238
rect 13795 32182 13863 32238
rect 13919 32182 13987 32238
rect 14043 32182 14111 32238
rect 14167 32182 14235 32238
rect 14291 32182 14359 32238
rect 14415 32182 14483 32238
rect 14539 32182 14607 32238
rect 14663 32182 14673 32238
rect 12861 32114 14673 32182
rect 12861 32058 12871 32114
rect 12927 32058 12995 32114
rect 13051 32058 13119 32114
rect 13175 32058 13243 32114
rect 13299 32058 13367 32114
rect 13423 32058 13491 32114
rect 13547 32058 13615 32114
rect 13671 32058 13739 32114
rect 13795 32058 13863 32114
rect 13919 32058 13987 32114
rect 14043 32058 14111 32114
rect 14167 32058 14235 32114
rect 14291 32058 14359 32114
rect 14415 32058 14483 32114
rect 14539 32058 14607 32114
rect 14663 32058 14673 32114
rect 12861 31990 14673 32058
rect 12861 31934 12871 31990
rect 12927 31934 12995 31990
rect 13051 31934 13119 31990
rect 13175 31934 13243 31990
rect 13299 31934 13367 31990
rect 13423 31934 13491 31990
rect 13547 31934 13615 31990
rect 13671 31934 13739 31990
rect 13795 31934 13863 31990
rect 13919 31934 13987 31990
rect 14043 31934 14111 31990
rect 14167 31934 14235 31990
rect 14291 31934 14359 31990
rect 14415 31934 14483 31990
rect 14539 31934 14607 31990
rect 14663 31934 14673 31990
rect 12861 31866 14673 31934
rect 12861 31810 12871 31866
rect 12927 31810 12995 31866
rect 13051 31810 13119 31866
rect 13175 31810 13243 31866
rect 13299 31810 13367 31866
rect 13423 31810 13491 31866
rect 13547 31810 13615 31866
rect 13671 31810 13739 31866
rect 13795 31810 13863 31866
rect 13919 31810 13987 31866
rect 14043 31810 14111 31866
rect 14167 31810 14235 31866
rect 14291 31810 14359 31866
rect 14415 31810 14483 31866
rect 14539 31810 14607 31866
rect 14663 31810 14673 31866
rect 12861 31742 14673 31810
rect 12861 31686 12871 31742
rect 12927 31686 12995 31742
rect 13051 31686 13119 31742
rect 13175 31686 13243 31742
rect 13299 31686 13367 31742
rect 13423 31686 13491 31742
rect 13547 31686 13615 31742
rect 13671 31686 13739 31742
rect 13795 31686 13863 31742
rect 13919 31686 13987 31742
rect 14043 31686 14111 31742
rect 14167 31686 14235 31742
rect 14291 31686 14359 31742
rect 14415 31686 14483 31742
rect 14539 31686 14607 31742
rect 14663 31686 14673 31742
rect 12861 31618 14673 31686
rect 12861 31562 12871 31618
rect 12927 31562 12995 31618
rect 13051 31562 13119 31618
rect 13175 31562 13243 31618
rect 13299 31562 13367 31618
rect 13423 31562 13491 31618
rect 13547 31562 13615 31618
rect 13671 31562 13739 31618
rect 13795 31562 13863 31618
rect 13919 31562 13987 31618
rect 14043 31562 14111 31618
rect 14167 31562 14235 31618
rect 14291 31562 14359 31618
rect 14415 31562 14483 31618
rect 14539 31562 14607 31618
rect 14663 31562 14673 31618
rect 12861 31494 14673 31562
rect 12861 31438 12871 31494
rect 12927 31438 12995 31494
rect 13051 31438 13119 31494
rect 13175 31438 13243 31494
rect 13299 31438 13367 31494
rect 13423 31438 13491 31494
rect 13547 31438 13615 31494
rect 13671 31438 13739 31494
rect 13795 31438 13863 31494
rect 13919 31438 13987 31494
rect 14043 31438 14111 31494
rect 14167 31438 14235 31494
rect 14291 31438 14359 31494
rect 14415 31438 14483 31494
rect 14539 31438 14607 31494
rect 14663 31438 14673 31494
rect 12861 31370 14673 31438
rect 12861 31314 12871 31370
rect 12927 31314 12995 31370
rect 13051 31314 13119 31370
rect 13175 31314 13243 31370
rect 13299 31314 13367 31370
rect 13423 31314 13491 31370
rect 13547 31314 13615 31370
rect 13671 31314 13739 31370
rect 13795 31314 13863 31370
rect 13919 31314 13987 31370
rect 14043 31314 14111 31370
rect 14167 31314 14235 31370
rect 14291 31314 14359 31370
rect 14415 31314 14483 31370
rect 14539 31314 14607 31370
rect 14663 31314 14673 31370
rect 12861 31246 14673 31314
rect 12861 31190 12871 31246
rect 12927 31190 12995 31246
rect 13051 31190 13119 31246
rect 13175 31190 13243 31246
rect 13299 31190 13367 31246
rect 13423 31190 13491 31246
rect 13547 31190 13615 31246
rect 13671 31190 13739 31246
rect 13795 31190 13863 31246
rect 13919 31190 13987 31246
rect 14043 31190 14111 31246
rect 14167 31190 14235 31246
rect 14291 31190 14359 31246
rect 14415 31190 14483 31246
rect 14539 31190 14607 31246
rect 14663 31190 14673 31246
rect 12861 31122 14673 31190
rect 12861 31066 12871 31122
rect 12927 31066 12995 31122
rect 13051 31066 13119 31122
rect 13175 31066 13243 31122
rect 13299 31066 13367 31122
rect 13423 31066 13491 31122
rect 13547 31066 13615 31122
rect 13671 31066 13739 31122
rect 13795 31066 13863 31122
rect 13919 31066 13987 31122
rect 14043 31066 14111 31122
rect 14167 31066 14235 31122
rect 14291 31066 14359 31122
rect 14415 31066 14483 31122
rect 14539 31066 14607 31122
rect 14663 31066 14673 31122
rect 12861 30998 14673 31066
rect 12861 30942 12871 30998
rect 12927 30942 12995 30998
rect 13051 30942 13119 30998
rect 13175 30942 13243 30998
rect 13299 30942 13367 30998
rect 13423 30942 13491 30998
rect 13547 30942 13615 30998
rect 13671 30942 13739 30998
rect 13795 30942 13863 30998
rect 13919 30942 13987 30998
rect 14043 30942 14111 30998
rect 14167 30942 14235 30998
rect 14291 30942 14359 30998
rect 14415 30942 14483 30998
rect 14539 30942 14607 30998
rect 14663 30942 14673 30998
rect 12861 30874 14673 30942
rect 12861 30818 12871 30874
rect 12927 30818 12995 30874
rect 13051 30818 13119 30874
rect 13175 30818 13243 30874
rect 13299 30818 13367 30874
rect 13423 30818 13491 30874
rect 13547 30818 13615 30874
rect 13671 30818 13739 30874
rect 13795 30818 13863 30874
rect 13919 30818 13987 30874
rect 14043 30818 14111 30874
rect 14167 30818 14235 30874
rect 14291 30818 14359 30874
rect 14415 30818 14483 30874
rect 14539 30818 14607 30874
rect 14663 30818 14673 30874
rect 12861 30750 14673 30818
rect 12861 30694 12871 30750
rect 12927 30694 12995 30750
rect 13051 30694 13119 30750
rect 13175 30694 13243 30750
rect 13299 30694 13367 30750
rect 13423 30694 13491 30750
rect 13547 30694 13615 30750
rect 13671 30694 13739 30750
rect 13795 30694 13863 30750
rect 13919 30694 13987 30750
rect 14043 30694 14111 30750
rect 14167 30694 14235 30750
rect 14291 30694 14359 30750
rect 14415 30694 14483 30750
rect 14539 30694 14607 30750
rect 14663 30694 14673 30750
rect 12861 30626 14673 30694
rect 12861 30570 12871 30626
rect 12927 30570 12995 30626
rect 13051 30570 13119 30626
rect 13175 30570 13243 30626
rect 13299 30570 13367 30626
rect 13423 30570 13491 30626
rect 13547 30570 13615 30626
rect 13671 30570 13739 30626
rect 13795 30570 13863 30626
rect 13919 30570 13987 30626
rect 14043 30570 14111 30626
rect 14167 30570 14235 30626
rect 14291 30570 14359 30626
rect 14415 30570 14483 30626
rect 14539 30570 14607 30626
rect 14663 30570 14673 30626
rect 12861 30502 14673 30570
rect 12861 30446 12871 30502
rect 12927 30446 12995 30502
rect 13051 30446 13119 30502
rect 13175 30446 13243 30502
rect 13299 30446 13367 30502
rect 13423 30446 13491 30502
rect 13547 30446 13615 30502
rect 13671 30446 13739 30502
rect 13795 30446 13863 30502
rect 13919 30446 13987 30502
rect 14043 30446 14111 30502
rect 14167 30446 14235 30502
rect 14291 30446 14359 30502
rect 14415 30446 14483 30502
rect 14539 30446 14607 30502
rect 14663 30446 14673 30502
rect 12861 30436 14673 30446
rect 305 30148 2117 30158
rect 305 30092 315 30148
rect 371 30092 439 30148
rect 495 30092 563 30148
rect 619 30092 687 30148
rect 743 30092 811 30148
rect 867 30092 935 30148
rect 991 30092 1059 30148
rect 1115 30092 1183 30148
rect 1239 30092 1307 30148
rect 1363 30092 1431 30148
rect 1487 30092 1555 30148
rect 1611 30092 1679 30148
rect 1735 30092 1803 30148
rect 1859 30092 1927 30148
rect 1983 30092 2051 30148
rect 2107 30092 2117 30148
rect 305 30024 2117 30092
rect 305 29968 315 30024
rect 371 29968 439 30024
rect 495 29968 563 30024
rect 619 29968 687 30024
rect 743 29968 811 30024
rect 867 29968 935 30024
rect 991 29968 1059 30024
rect 1115 29968 1183 30024
rect 1239 29968 1307 30024
rect 1363 29968 1431 30024
rect 1487 29968 1555 30024
rect 1611 29968 1679 30024
rect 1735 29968 1803 30024
rect 1859 29968 1927 30024
rect 1983 29968 2051 30024
rect 2107 29968 2117 30024
rect 305 29900 2117 29968
rect 305 29844 315 29900
rect 371 29844 439 29900
rect 495 29844 563 29900
rect 619 29844 687 29900
rect 743 29844 811 29900
rect 867 29844 935 29900
rect 991 29844 1059 29900
rect 1115 29844 1183 29900
rect 1239 29844 1307 29900
rect 1363 29844 1431 29900
rect 1487 29844 1555 29900
rect 1611 29844 1679 29900
rect 1735 29844 1803 29900
rect 1859 29844 1927 29900
rect 1983 29844 2051 29900
rect 2107 29844 2117 29900
rect 305 29776 2117 29844
rect 305 29720 315 29776
rect 371 29720 439 29776
rect 495 29720 563 29776
rect 619 29720 687 29776
rect 743 29720 811 29776
rect 867 29720 935 29776
rect 991 29720 1059 29776
rect 1115 29720 1183 29776
rect 1239 29720 1307 29776
rect 1363 29720 1431 29776
rect 1487 29720 1555 29776
rect 1611 29720 1679 29776
rect 1735 29720 1803 29776
rect 1859 29720 1927 29776
rect 1983 29720 2051 29776
rect 2107 29720 2117 29776
rect 305 29652 2117 29720
rect 305 29596 315 29652
rect 371 29596 439 29652
rect 495 29596 563 29652
rect 619 29596 687 29652
rect 743 29596 811 29652
rect 867 29596 935 29652
rect 991 29596 1059 29652
rect 1115 29596 1183 29652
rect 1239 29596 1307 29652
rect 1363 29596 1431 29652
rect 1487 29596 1555 29652
rect 1611 29596 1679 29652
rect 1735 29596 1803 29652
rect 1859 29596 1927 29652
rect 1983 29596 2051 29652
rect 2107 29596 2117 29652
rect 305 29528 2117 29596
rect 305 29472 315 29528
rect 371 29472 439 29528
rect 495 29472 563 29528
rect 619 29472 687 29528
rect 743 29472 811 29528
rect 867 29472 935 29528
rect 991 29472 1059 29528
rect 1115 29472 1183 29528
rect 1239 29472 1307 29528
rect 1363 29472 1431 29528
rect 1487 29472 1555 29528
rect 1611 29472 1679 29528
rect 1735 29472 1803 29528
rect 1859 29472 1927 29528
rect 1983 29472 2051 29528
rect 2107 29472 2117 29528
rect 305 29404 2117 29472
rect 305 29348 315 29404
rect 371 29348 439 29404
rect 495 29348 563 29404
rect 619 29348 687 29404
rect 743 29348 811 29404
rect 867 29348 935 29404
rect 991 29348 1059 29404
rect 1115 29348 1183 29404
rect 1239 29348 1307 29404
rect 1363 29348 1431 29404
rect 1487 29348 1555 29404
rect 1611 29348 1679 29404
rect 1735 29348 1803 29404
rect 1859 29348 1927 29404
rect 1983 29348 2051 29404
rect 2107 29348 2117 29404
rect 305 29280 2117 29348
rect 305 29224 315 29280
rect 371 29224 439 29280
rect 495 29224 563 29280
rect 619 29224 687 29280
rect 743 29224 811 29280
rect 867 29224 935 29280
rect 991 29224 1059 29280
rect 1115 29224 1183 29280
rect 1239 29224 1307 29280
rect 1363 29224 1431 29280
rect 1487 29224 1555 29280
rect 1611 29224 1679 29280
rect 1735 29224 1803 29280
rect 1859 29224 1927 29280
rect 1983 29224 2051 29280
rect 2107 29224 2117 29280
rect 305 29156 2117 29224
rect 305 29100 315 29156
rect 371 29100 439 29156
rect 495 29100 563 29156
rect 619 29100 687 29156
rect 743 29100 811 29156
rect 867 29100 935 29156
rect 991 29100 1059 29156
rect 1115 29100 1183 29156
rect 1239 29100 1307 29156
rect 1363 29100 1431 29156
rect 1487 29100 1555 29156
rect 1611 29100 1679 29156
rect 1735 29100 1803 29156
rect 1859 29100 1927 29156
rect 1983 29100 2051 29156
rect 2107 29100 2117 29156
rect 305 29032 2117 29100
rect 305 28976 315 29032
rect 371 28976 439 29032
rect 495 28976 563 29032
rect 619 28976 687 29032
rect 743 28976 811 29032
rect 867 28976 935 29032
rect 991 28976 1059 29032
rect 1115 28976 1183 29032
rect 1239 28976 1307 29032
rect 1363 28976 1431 29032
rect 1487 28976 1555 29032
rect 1611 28976 1679 29032
rect 1735 28976 1803 29032
rect 1859 28976 1927 29032
rect 1983 28976 2051 29032
rect 2107 28976 2117 29032
rect 305 28908 2117 28976
rect 305 28852 315 28908
rect 371 28852 439 28908
rect 495 28852 563 28908
rect 619 28852 687 28908
rect 743 28852 811 28908
rect 867 28852 935 28908
rect 991 28852 1059 28908
rect 1115 28852 1183 28908
rect 1239 28852 1307 28908
rect 1363 28852 1431 28908
rect 1487 28852 1555 28908
rect 1611 28852 1679 28908
rect 1735 28852 1803 28908
rect 1859 28852 1927 28908
rect 1983 28852 2051 28908
rect 2107 28852 2117 28908
rect 305 28842 2117 28852
rect 2798 30148 4734 30158
rect 2798 30092 2808 30148
rect 2864 30092 2932 30148
rect 2988 30092 3056 30148
rect 3112 30092 3180 30148
rect 3236 30092 3304 30148
rect 3360 30092 3428 30148
rect 3484 30092 3552 30148
rect 3608 30092 3676 30148
rect 3732 30092 3800 30148
rect 3856 30092 3924 30148
rect 3980 30092 4048 30148
rect 4104 30092 4172 30148
rect 4228 30092 4296 30148
rect 4352 30092 4420 30148
rect 4476 30092 4544 30148
rect 4600 30092 4668 30148
rect 4724 30092 4734 30148
rect 2798 30024 4734 30092
rect 2798 29968 2808 30024
rect 2864 29968 2932 30024
rect 2988 29968 3056 30024
rect 3112 29968 3180 30024
rect 3236 29968 3304 30024
rect 3360 29968 3428 30024
rect 3484 29968 3552 30024
rect 3608 29968 3676 30024
rect 3732 29968 3800 30024
rect 3856 29968 3924 30024
rect 3980 29968 4048 30024
rect 4104 29968 4172 30024
rect 4228 29968 4296 30024
rect 4352 29968 4420 30024
rect 4476 29968 4544 30024
rect 4600 29968 4668 30024
rect 4724 29968 4734 30024
rect 2798 29900 4734 29968
rect 2798 29844 2808 29900
rect 2864 29844 2932 29900
rect 2988 29844 3056 29900
rect 3112 29844 3180 29900
rect 3236 29844 3304 29900
rect 3360 29844 3428 29900
rect 3484 29844 3552 29900
rect 3608 29844 3676 29900
rect 3732 29844 3800 29900
rect 3856 29844 3924 29900
rect 3980 29844 4048 29900
rect 4104 29844 4172 29900
rect 4228 29844 4296 29900
rect 4352 29844 4420 29900
rect 4476 29844 4544 29900
rect 4600 29844 4668 29900
rect 4724 29844 4734 29900
rect 2798 29776 4734 29844
rect 2798 29720 2808 29776
rect 2864 29720 2932 29776
rect 2988 29720 3056 29776
rect 3112 29720 3180 29776
rect 3236 29720 3304 29776
rect 3360 29720 3428 29776
rect 3484 29720 3552 29776
rect 3608 29720 3676 29776
rect 3732 29720 3800 29776
rect 3856 29720 3924 29776
rect 3980 29720 4048 29776
rect 4104 29720 4172 29776
rect 4228 29720 4296 29776
rect 4352 29720 4420 29776
rect 4476 29720 4544 29776
rect 4600 29720 4668 29776
rect 4724 29720 4734 29776
rect 2798 29652 4734 29720
rect 2798 29596 2808 29652
rect 2864 29596 2932 29652
rect 2988 29596 3056 29652
rect 3112 29596 3180 29652
rect 3236 29596 3304 29652
rect 3360 29596 3428 29652
rect 3484 29596 3552 29652
rect 3608 29596 3676 29652
rect 3732 29596 3800 29652
rect 3856 29596 3924 29652
rect 3980 29596 4048 29652
rect 4104 29596 4172 29652
rect 4228 29596 4296 29652
rect 4352 29596 4420 29652
rect 4476 29596 4544 29652
rect 4600 29596 4668 29652
rect 4724 29596 4734 29652
rect 2798 29528 4734 29596
rect 2798 29472 2808 29528
rect 2864 29472 2932 29528
rect 2988 29472 3056 29528
rect 3112 29472 3180 29528
rect 3236 29472 3304 29528
rect 3360 29472 3428 29528
rect 3484 29472 3552 29528
rect 3608 29472 3676 29528
rect 3732 29472 3800 29528
rect 3856 29472 3924 29528
rect 3980 29472 4048 29528
rect 4104 29472 4172 29528
rect 4228 29472 4296 29528
rect 4352 29472 4420 29528
rect 4476 29472 4544 29528
rect 4600 29472 4668 29528
rect 4724 29472 4734 29528
rect 2798 29404 4734 29472
rect 2798 29348 2808 29404
rect 2864 29348 2932 29404
rect 2988 29348 3056 29404
rect 3112 29348 3180 29404
rect 3236 29348 3304 29404
rect 3360 29348 3428 29404
rect 3484 29348 3552 29404
rect 3608 29348 3676 29404
rect 3732 29348 3800 29404
rect 3856 29348 3924 29404
rect 3980 29348 4048 29404
rect 4104 29348 4172 29404
rect 4228 29348 4296 29404
rect 4352 29348 4420 29404
rect 4476 29348 4544 29404
rect 4600 29348 4668 29404
rect 4724 29348 4734 29404
rect 2798 29280 4734 29348
rect 2798 29224 2808 29280
rect 2864 29224 2932 29280
rect 2988 29224 3056 29280
rect 3112 29224 3180 29280
rect 3236 29224 3304 29280
rect 3360 29224 3428 29280
rect 3484 29224 3552 29280
rect 3608 29224 3676 29280
rect 3732 29224 3800 29280
rect 3856 29224 3924 29280
rect 3980 29224 4048 29280
rect 4104 29224 4172 29280
rect 4228 29224 4296 29280
rect 4352 29224 4420 29280
rect 4476 29224 4544 29280
rect 4600 29224 4668 29280
rect 4724 29224 4734 29280
rect 2798 29156 4734 29224
rect 2798 29100 2808 29156
rect 2864 29100 2932 29156
rect 2988 29100 3056 29156
rect 3112 29100 3180 29156
rect 3236 29100 3304 29156
rect 3360 29100 3428 29156
rect 3484 29100 3552 29156
rect 3608 29100 3676 29156
rect 3732 29100 3800 29156
rect 3856 29100 3924 29156
rect 3980 29100 4048 29156
rect 4104 29100 4172 29156
rect 4228 29100 4296 29156
rect 4352 29100 4420 29156
rect 4476 29100 4544 29156
rect 4600 29100 4668 29156
rect 4724 29100 4734 29156
rect 2798 29032 4734 29100
rect 2798 28976 2808 29032
rect 2864 28976 2932 29032
rect 2988 28976 3056 29032
rect 3112 28976 3180 29032
rect 3236 28976 3304 29032
rect 3360 28976 3428 29032
rect 3484 28976 3552 29032
rect 3608 28976 3676 29032
rect 3732 28976 3800 29032
rect 3856 28976 3924 29032
rect 3980 28976 4048 29032
rect 4104 28976 4172 29032
rect 4228 28976 4296 29032
rect 4352 28976 4420 29032
rect 4476 28976 4544 29032
rect 4600 28976 4668 29032
rect 4724 28976 4734 29032
rect 2798 28908 4734 28976
rect 2798 28852 2808 28908
rect 2864 28852 2932 28908
rect 2988 28852 3056 28908
rect 3112 28852 3180 28908
rect 3236 28852 3304 28908
rect 3360 28852 3428 28908
rect 3484 28852 3552 28908
rect 3608 28852 3676 28908
rect 3732 28852 3800 28908
rect 3856 28852 3924 28908
rect 3980 28852 4048 28908
rect 4104 28852 4172 28908
rect 4228 28852 4296 28908
rect 4352 28852 4420 28908
rect 4476 28852 4544 28908
rect 4600 28852 4668 28908
rect 4724 28852 4734 28908
rect 2798 28842 4734 28852
rect 5168 30148 7104 30158
rect 5168 30092 5178 30148
rect 5234 30092 5302 30148
rect 5358 30092 5426 30148
rect 5482 30092 5550 30148
rect 5606 30092 5674 30148
rect 5730 30092 5798 30148
rect 5854 30092 5922 30148
rect 5978 30092 6046 30148
rect 6102 30092 6170 30148
rect 6226 30092 6294 30148
rect 6350 30092 6418 30148
rect 6474 30092 6542 30148
rect 6598 30092 6666 30148
rect 6722 30092 6790 30148
rect 6846 30092 6914 30148
rect 6970 30092 7038 30148
rect 7094 30092 7104 30148
rect 5168 30024 7104 30092
rect 5168 29968 5178 30024
rect 5234 29968 5302 30024
rect 5358 29968 5426 30024
rect 5482 29968 5550 30024
rect 5606 29968 5674 30024
rect 5730 29968 5798 30024
rect 5854 29968 5922 30024
rect 5978 29968 6046 30024
rect 6102 29968 6170 30024
rect 6226 29968 6294 30024
rect 6350 29968 6418 30024
rect 6474 29968 6542 30024
rect 6598 29968 6666 30024
rect 6722 29968 6790 30024
rect 6846 29968 6914 30024
rect 6970 29968 7038 30024
rect 7094 29968 7104 30024
rect 5168 29900 7104 29968
rect 5168 29844 5178 29900
rect 5234 29844 5302 29900
rect 5358 29844 5426 29900
rect 5482 29844 5550 29900
rect 5606 29844 5674 29900
rect 5730 29844 5798 29900
rect 5854 29844 5922 29900
rect 5978 29844 6046 29900
rect 6102 29844 6170 29900
rect 6226 29844 6294 29900
rect 6350 29844 6418 29900
rect 6474 29844 6542 29900
rect 6598 29844 6666 29900
rect 6722 29844 6790 29900
rect 6846 29844 6914 29900
rect 6970 29844 7038 29900
rect 7094 29844 7104 29900
rect 5168 29776 7104 29844
rect 5168 29720 5178 29776
rect 5234 29720 5302 29776
rect 5358 29720 5426 29776
rect 5482 29720 5550 29776
rect 5606 29720 5674 29776
rect 5730 29720 5798 29776
rect 5854 29720 5922 29776
rect 5978 29720 6046 29776
rect 6102 29720 6170 29776
rect 6226 29720 6294 29776
rect 6350 29720 6418 29776
rect 6474 29720 6542 29776
rect 6598 29720 6666 29776
rect 6722 29720 6790 29776
rect 6846 29720 6914 29776
rect 6970 29720 7038 29776
rect 7094 29720 7104 29776
rect 5168 29652 7104 29720
rect 5168 29596 5178 29652
rect 5234 29596 5302 29652
rect 5358 29596 5426 29652
rect 5482 29596 5550 29652
rect 5606 29596 5674 29652
rect 5730 29596 5798 29652
rect 5854 29596 5922 29652
rect 5978 29596 6046 29652
rect 6102 29596 6170 29652
rect 6226 29596 6294 29652
rect 6350 29596 6418 29652
rect 6474 29596 6542 29652
rect 6598 29596 6666 29652
rect 6722 29596 6790 29652
rect 6846 29596 6914 29652
rect 6970 29596 7038 29652
rect 7094 29596 7104 29652
rect 5168 29528 7104 29596
rect 5168 29472 5178 29528
rect 5234 29472 5302 29528
rect 5358 29472 5426 29528
rect 5482 29472 5550 29528
rect 5606 29472 5674 29528
rect 5730 29472 5798 29528
rect 5854 29472 5922 29528
rect 5978 29472 6046 29528
rect 6102 29472 6170 29528
rect 6226 29472 6294 29528
rect 6350 29472 6418 29528
rect 6474 29472 6542 29528
rect 6598 29472 6666 29528
rect 6722 29472 6790 29528
rect 6846 29472 6914 29528
rect 6970 29472 7038 29528
rect 7094 29472 7104 29528
rect 5168 29404 7104 29472
rect 5168 29348 5178 29404
rect 5234 29348 5302 29404
rect 5358 29348 5426 29404
rect 5482 29348 5550 29404
rect 5606 29348 5674 29404
rect 5730 29348 5798 29404
rect 5854 29348 5922 29404
rect 5978 29348 6046 29404
rect 6102 29348 6170 29404
rect 6226 29348 6294 29404
rect 6350 29348 6418 29404
rect 6474 29348 6542 29404
rect 6598 29348 6666 29404
rect 6722 29348 6790 29404
rect 6846 29348 6914 29404
rect 6970 29348 7038 29404
rect 7094 29348 7104 29404
rect 5168 29280 7104 29348
rect 5168 29224 5178 29280
rect 5234 29224 5302 29280
rect 5358 29224 5426 29280
rect 5482 29224 5550 29280
rect 5606 29224 5674 29280
rect 5730 29224 5798 29280
rect 5854 29224 5922 29280
rect 5978 29224 6046 29280
rect 6102 29224 6170 29280
rect 6226 29224 6294 29280
rect 6350 29224 6418 29280
rect 6474 29224 6542 29280
rect 6598 29224 6666 29280
rect 6722 29224 6790 29280
rect 6846 29224 6914 29280
rect 6970 29224 7038 29280
rect 7094 29224 7104 29280
rect 5168 29156 7104 29224
rect 5168 29100 5178 29156
rect 5234 29100 5302 29156
rect 5358 29100 5426 29156
rect 5482 29100 5550 29156
rect 5606 29100 5674 29156
rect 5730 29100 5798 29156
rect 5854 29100 5922 29156
rect 5978 29100 6046 29156
rect 6102 29100 6170 29156
rect 6226 29100 6294 29156
rect 6350 29100 6418 29156
rect 6474 29100 6542 29156
rect 6598 29100 6666 29156
rect 6722 29100 6790 29156
rect 6846 29100 6914 29156
rect 6970 29100 7038 29156
rect 7094 29100 7104 29156
rect 5168 29032 7104 29100
rect 5168 28976 5178 29032
rect 5234 28976 5302 29032
rect 5358 28976 5426 29032
rect 5482 28976 5550 29032
rect 5606 28976 5674 29032
rect 5730 28976 5798 29032
rect 5854 28976 5922 29032
rect 5978 28976 6046 29032
rect 6102 28976 6170 29032
rect 6226 28976 6294 29032
rect 6350 28976 6418 29032
rect 6474 28976 6542 29032
rect 6598 28976 6666 29032
rect 6722 28976 6790 29032
rect 6846 28976 6914 29032
rect 6970 28976 7038 29032
rect 7094 28976 7104 29032
rect 5168 28908 7104 28976
rect 5168 28852 5178 28908
rect 5234 28852 5302 28908
rect 5358 28852 5426 28908
rect 5482 28852 5550 28908
rect 5606 28852 5674 28908
rect 5730 28852 5798 28908
rect 5854 28852 5922 28908
rect 5978 28852 6046 28908
rect 6102 28852 6170 28908
rect 6226 28852 6294 28908
rect 6350 28852 6418 28908
rect 6474 28852 6542 28908
rect 6598 28852 6666 28908
rect 6722 28852 6790 28908
rect 6846 28852 6914 28908
rect 6970 28852 7038 28908
rect 7094 28852 7104 28908
rect 5168 28842 7104 28852
rect 7874 30148 9810 30158
rect 7874 30092 7884 30148
rect 7940 30092 8008 30148
rect 8064 30092 8132 30148
rect 8188 30092 8256 30148
rect 8312 30092 8380 30148
rect 8436 30092 8504 30148
rect 8560 30092 8628 30148
rect 8684 30092 8752 30148
rect 8808 30092 8876 30148
rect 8932 30092 9000 30148
rect 9056 30092 9124 30148
rect 9180 30092 9248 30148
rect 9304 30092 9372 30148
rect 9428 30092 9496 30148
rect 9552 30092 9620 30148
rect 9676 30092 9744 30148
rect 9800 30092 9810 30148
rect 7874 30024 9810 30092
rect 7874 29968 7884 30024
rect 7940 29968 8008 30024
rect 8064 29968 8132 30024
rect 8188 29968 8256 30024
rect 8312 29968 8380 30024
rect 8436 29968 8504 30024
rect 8560 29968 8628 30024
rect 8684 29968 8752 30024
rect 8808 29968 8876 30024
rect 8932 29968 9000 30024
rect 9056 29968 9124 30024
rect 9180 29968 9248 30024
rect 9304 29968 9372 30024
rect 9428 29968 9496 30024
rect 9552 29968 9620 30024
rect 9676 29968 9744 30024
rect 9800 29968 9810 30024
rect 7874 29900 9810 29968
rect 7874 29844 7884 29900
rect 7940 29844 8008 29900
rect 8064 29844 8132 29900
rect 8188 29844 8256 29900
rect 8312 29844 8380 29900
rect 8436 29844 8504 29900
rect 8560 29844 8628 29900
rect 8684 29844 8752 29900
rect 8808 29844 8876 29900
rect 8932 29844 9000 29900
rect 9056 29844 9124 29900
rect 9180 29844 9248 29900
rect 9304 29844 9372 29900
rect 9428 29844 9496 29900
rect 9552 29844 9620 29900
rect 9676 29844 9744 29900
rect 9800 29844 9810 29900
rect 7874 29776 9810 29844
rect 7874 29720 7884 29776
rect 7940 29720 8008 29776
rect 8064 29720 8132 29776
rect 8188 29720 8256 29776
rect 8312 29720 8380 29776
rect 8436 29720 8504 29776
rect 8560 29720 8628 29776
rect 8684 29720 8752 29776
rect 8808 29720 8876 29776
rect 8932 29720 9000 29776
rect 9056 29720 9124 29776
rect 9180 29720 9248 29776
rect 9304 29720 9372 29776
rect 9428 29720 9496 29776
rect 9552 29720 9620 29776
rect 9676 29720 9744 29776
rect 9800 29720 9810 29776
rect 7874 29652 9810 29720
rect 7874 29596 7884 29652
rect 7940 29596 8008 29652
rect 8064 29596 8132 29652
rect 8188 29596 8256 29652
rect 8312 29596 8380 29652
rect 8436 29596 8504 29652
rect 8560 29596 8628 29652
rect 8684 29596 8752 29652
rect 8808 29596 8876 29652
rect 8932 29596 9000 29652
rect 9056 29596 9124 29652
rect 9180 29596 9248 29652
rect 9304 29596 9372 29652
rect 9428 29596 9496 29652
rect 9552 29596 9620 29652
rect 9676 29596 9744 29652
rect 9800 29596 9810 29652
rect 7874 29528 9810 29596
rect 7874 29472 7884 29528
rect 7940 29472 8008 29528
rect 8064 29472 8132 29528
rect 8188 29472 8256 29528
rect 8312 29472 8380 29528
rect 8436 29472 8504 29528
rect 8560 29472 8628 29528
rect 8684 29472 8752 29528
rect 8808 29472 8876 29528
rect 8932 29472 9000 29528
rect 9056 29472 9124 29528
rect 9180 29472 9248 29528
rect 9304 29472 9372 29528
rect 9428 29472 9496 29528
rect 9552 29472 9620 29528
rect 9676 29472 9744 29528
rect 9800 29472 9810 29528
rect 7874 29404 9810 29472
rect 7874 29348 7884 29404
rect 7940 29348 8008 29404
rect 8064 29348 8132 29404
rect 8188 29348 8256 29404
rect 8312 29348 8380 29404
rect 8436 29348 8504 29404
rect 8560 29348 8628 29404
rect 8684 29348 8752 29404
rect 8808 29348 8876 29404
rect 8932 29348 9000 29404
rect 9056 29348 9124 29404
rect 9180 29348 9248 29404
rect 9304 29348 9372 29404
rect 9428 29348 9496 29404
rect 9552 29348 9620 29404
rect 9676 29348 9744 29404
rect 9800 29348 9810 29404
rect 7874 29280 9810 29348
rect 7874 29224 7884 29280
rect 7940 29224 8008 29280
rect 8064 29224 8132 29280
rect 8188 29224 8256 29280
rect 8312 29224 8380 29280
rect 8436 29224 8504 29280
rect 8560 29224 8628 29280
rect 8684 29224 8752 29280
rect 8808 29224 8876 29280
rect 8932 29224 9000 29280
rect 9056 29224 9124 29280
rect 9180 29224 9248 29280
rect 9304 29224 9372 29280
rect 9428 29224 9496 29280
rect 9552 29224 9620 29280
rect 9676 29224 9744 29280
rect 9800 29224 9810 29280
rect 7874 29156 9810 29224
rect 7874 29100 7884 29156
rect 7940 29100 8008 29156
rect 8064 29100 8132 29156
rect 8188 29100 8256 29156
rect 8312 29100 8380 29156
rect 8436 29100 8504 29156
rect 8560 29100 8628 29156
rect 8684 29100 8752 29156
rect 8808 29100 8876 29156
rect 8932 29100 9000 29156
rect 9056 29100 9124 29156
rect 9180 29100 9248 29156
rect 9304 29100 9372 29156
rect 9428 29100 9496 29156
rect 9552 29100 9620 29156
rect 9676 29100 9744 29156
rect 9800 29100 9810 29156
rect 7874 29032 9810 29100
rect 7874 28976 7884 29032
rect 7940 28976 8008 29032
rect 8064 28976 8132 29032
rect 8188 28976 8256 29032
rect 8312 28976 8380 29032
rect 8436 28976 8504 29032
rect 8560 28976 8628 29032
rect 8684 28976 8752 29032
rect 8808 28976 8876 29032
rect 8932 28976 9000 29032
rect 9056 28976 9124 29032
rect 9180 28976 9248 29032
rect 9304 28976 9372 29032
rect 9428 28976 9496 29032
rect 9552 28976 9620 29032
rect 9676 28976 9744 29032
rect 9800 28976 9810 29032
rect 7874 28908 9810 28976
rect 7874 28852 7884 28908
rect 7940 28852 8008 28908
rect 8064 28852 8132 28908
rect 8188 28852 8256 28908
rect 8312 28852 8380 28908
rect 8436 28852 8504 28908
rect 8560 28852 8628 28908
rect 8684 28852 8752 28908
rect 8808 28852 8876 28908
rect 8932 28852 9000 28908
rect 9056 28852 9124 28908
rect 9180 28852 9248 28908
rect 9304 28852 9372 28908
rect 9428 28852 9496 28908
rect 9552 28852 9620 28908
rect 9676 28852 9744 28908
rect 9800 28852 9810 28908
rect 7874 28842 9810 28852
rect 10244 30148 12180 30158
rect 10244 30092 10254 30148
rect 10310 30092 10378 30148
rect 10434 30092 10502 30148
rect 10558 30092 10626 30148
rect 10682 30092 10750 30148
rect 10806 30092 10874 30148
rect 10930 30092 10998 30148
rect 11054 30092 11122 30148
rect 11178 30092 11246 30148
rect 11302 30092 11370 30148
rect 11426 30092 11494 30148
rect 11550 30092 11618 30148
rect 11674 30092 11742 30148
rect 11798 30092 11866 30148
rect 11922 30092 11990 30148
rect 12046 30092 12114 30148
rect 12170 30092 12180 30148
rect 10244 30024 12180 30092
rect 10244 29968 10254 30024
rect 10310 29968 10378 30024
rect 10434 29968 10502 30024
rect 10558 29968 10626 30024
rect 10682 29968 10750 30024
rect 10806 29968 10874 30024
rect 10930 29968 10998 30024
rect 11054 29968 11122 30024
rect 11178 29968 11246 30024
rect 11302 29968 11370 30024
rect 11426 29968 11494 30024
rect 11550 29968 11618 30024
rect 11674 29968 11742 30024
rect 11798 29968 11866 30024
rect 11922 29968 11990 30024
rect 12046 29968 12114 30024
rect 12170 29968 12180 30024
rect 10244 29900 12180 29968
rect 10244 29844 10254 29900
rect 10310 29844 10378 29900
rect 10434 29844 10502 29900
rect 10558 29844 10626 29900
rect 10682 29844 10750 29900
rect 10806 29844 10874 29900
rect 10930 29844 10998 29900
rect 11054 29844 11122 29900
rect 11178 29844 11246 29900
rect 11302 29844 11370 29900
rect 11426 29844 11494 29900
rect 11550 29844 11618 29900
rect 11674 29844 11742 29900
rect 11798 29844 11866 29900
rect 11922 29844 11990 29900
rect 12046 29844 12114 29900
rect 12170 29844 12180 29900
rect 10244 29776 12180 29844
rect 10244 29720 10254 29776
rect 10310 29720 10378 29776
rect 10434 29720 10502 29776
rect 10558 29720 10626 29776
rect 10682 29720 10750 29776
rect 10806 29720 10874 29776
rect 10930 29720 10998 29776
rect 11054 29720 11122 29776
rect 11178 29720 11246 29776
rect 11302 29720 11370 29776
rect 11426 29720 11494 29776
rect 11550 29720 11618 29776
rect 11674 29720 11742 29776
rect 11798 29720 11866 29776
rect 11922 29720 11990 29776
rect 12046 29720 12114 29776
rect 12170 29720 12180 29776
rect 10244 29652 12180 29720
rect 10244 29596 10254 29652
rect 10310 29596 10378 29652
rect 10434 29596 10502 29652
rect 10558 29596 10626 29652
rect 10682 29596 10750 29652
rect 10806 29596 10874 29652
rect 10930 29596 10998 29652
rect 11054 29596 11122 29652
rect 11178 29596 11246 29652
rect 11302 29596 11370 29652
rect 11426 29596 11494 29652
rect 11550 29596 11618 29652
rect 11674 29596 11742 29652
rect 11798 29596 11866 29652
rect 11922 29596 11990 29652
rect 12046 29596 12114 29652
rect 12170 29596 12180 29652
rect 10244 29528 12180 29596
rect 10244 29472 10254 29528
rect 10310 29472 10378 29528
rect 10434 29472 10502 29528
rect 10558 29472 10626 29528
rect 10682 29472 10750 29528
rect 10806 29472 10874 29528
rect 10930 29472 10998 29528
rect 11054 29472 11122 29528
rect 11178 29472 11246 29528
rect 11302 29472 11370 29528
rect 11426 29472 11494 29528
rect 11550 29472 11618 29528
rect 11674 29472 11742 29528
rect 11798 29472 11866 29528
rect 11922 29472 11990 29528
rect 12046 29472 12114 29528
rect 12170 29472 12180 29528
rect 10244 29404 12180 29472
rect 10244 29348 10254 29404
rect 10310 29348 10378 29404
rect 10434 29348 10502 29404
rect 10558 29348 10626 29404
rect 10682 29348 10750 29404
rect 10806 29348 10874 29404
rect 10930 29348 10998 29404
rect 11054 29348 11122 29404
rect 11178 29348 11246 29404
rect 11302 29348 11370 29404
rect 11426 29348 11494 29404
rect 11550 29348 11618 29404
rect 11674 29348 11742 29404
rect 11798 29348 11866 29404
rect 11922 29348 11990 29404
rect 12046 29348 12114 29404
rect 12170 29348 12180 29404
rect 10244 29280 12180 29348
rect 10244 29224 10254 29280
rect 10310 29224 10378 29280
rect 10434 29224 10502 29280
rect 10558 29224 10626 29280
rect 10682 29224 10750 29280
rect 10806 29224 10874 29280
rect 10930 29224 10998 29280
rect 11054 29224 11122 29280
rect 11178 29224 11246 29280
rect 11302 29224 11370 29280
rect 11426 29224 11494 29280
rect 11550 29224 11618 29280
rect 11674 29224 11742 29280
rect 11798 29224 11866 29280
rect 11922 29224 11990 29280
rect 12046 29224 12114 29280
rect 12170 29224 12180 29280
rect 10244 29156 12180 29224
rect 10244 29100 10254 29156
rect 10310 29100 10378 29156
rect 10434 29100 10502 29156
rect 10558 29100 10626 29156
rect 10682 29100 10750 29156
rect 10806 29100 10874 29156
rect 10930 29100 10998 29156
rect 11054 29100 11122 29156
rect 11178 29100 11246 29156
rect 11302 29100 11370 29156
rect 11426 29100 11494 29156
rect 11550 29100 11618 29156
rect 11674 29100 11742 29156
rect 11798 29100 11866 29156
rect 11922 29100 11990 29156
rect 12046 29100 12114 29156
rect 12170 29100 12180 29156
rect 10244 29032 12180 29100
rect 10244 28976 10254 29032
rect 10310 28976 10378 29032
rect 10434 28976 10502 29032
rect 10558 28976 10626 29032
rect 10682 28976 10750 29032
rect 10806 28976 10874 29032
rect 10930 28976 10998 29032
rect 11054 28976 11122 29032
rect 11178 28976 11246 29032
rect 11302 28976 11370 29032
rect 11426 28976 11494 29032
rect 11550 28976 11618 29032
rect 11674 28976 11742 29032
rect 11798 28976 11866 29032
rect 11922 28976 11990 29032
rect 12046 28976 12114 29032
rect 12170 28976 12180 29032
rect 10244 28908 12180 28976
rect 10244 28852 10254 28908
rect 10310 28852 10378 28908
rect 10434 28852 10502 28908
rect 10558 28852 10626 28908
rect 10682 28852 10750 28908
rect 10806 28852 10874 28908
rect 10930 28852 10998 28908
rect 11054 28852 11122 28908
rect 11178 28852 11246 28908
rect 11302 28852 11370 28908
rect 11426 28852 11494 28908
rect 11550 28852 11618 28908
rect 11674 28852 11742 28908
rect 11798 28852 11866 28908
rect 11922 28852 11990 28908
rect 12046 28852 12114 28908
rect 12170 28852 12180 28908
rect 10244 28842 12180 28852
rect 12861 30148 14673 30158
rect 12861 30092 12871 30148
rect 12927 30092 12995 30148
rect 13051 30092 13119 30148
rect 13175 30092 13243 30148
rect 13299 30092 13367 30148
rect 13423 30092 13491 30148
rect 13547 30092 13615 30148
rect 13671 30092 13739 30148
rect 13795 30092 13863 30148
rect 13919 30092 13987 30148
rect 14043 30092 14111 30148
rect 14167 30092 14235 30148
rect 14291 30092 14359 30148
rect 14415 30092 14483 30148
rect 14539 30092 14607 30148
rect 14663 30092 14673 30148
rect 12861 30024 14673 30092
rect 12861 29968 12871 30024
rect 12927 29968 12995 30024
rect 13051 29968 13119 30024
rect 13175 29968 13243 30024
rect 13299 29968 13367 30024
rect 13423 29968 13491 30024
rect 13547 29968 13615 30024
rect 13671 29968 13739 30024
rect 13795 29968 13863 30024
rect 13919 29968 13987 30024
rect 14043 29968 14111 30024
rect 14167 29968 14235 30024
rect 14291 29968 14359 30024
rect 14415 29968 14483 30024
rect 14539 29968 14607 30024
rect 14663 29968 14673 30024
rect 12861 29900 14673 29968
rect 12861 29844 12871 29900
rect 12927 29844 12995 29900
rect 13051 29844 13119 29900
rect 13175 29844 13243 29900
rect 13299 29844 13367 29900
rect 13423 29844 13491 29900
rect 13547 29844 13615 29900
rect 13671 29844 13739 29900
rect 13795 29844 13863 29900
rect 13919 29844 13987 29900
rect 14043 29844 14111 29900
rect 14167 29844 14235 29900
rect 14291 29844 14359 29900
rect 14415 29844 14483 29900
rect 14539 29844 14607 29900
rect 14663 29844 14673 29900
rect 12861 29776 14673 29844
rect 12861 29720 12871 29776
rect 12927 29720 12995 29776
rect 13051 29720 13119 29776
rect 13175 29720 13243 29776
rect 13299 29720 13367 29776
rect 13423 29720 13491 29776
rect 13547 29720 13615 29776
rect 13671 29720 13739 29776
rect 13795 29720 13863 29776
rect 13919 29720 13987 29776
rect 14043 29720 14111 29776
rect 14167 29720 14235 29776
rect 14291 29720 14359 29776
rect 14415 29720 14483 29776
rect 14539 29720 14607 29776
rect 14663 29720 14673 29776
rect 12861 29652 14673 29720
rect 12861 29596 12871 29652
rect 12927 29596 12995 29652
rect 13051 29596 13119 29652
rect 13175 29596 13243 29652
rect 13299 29596 13367 29652
rect 13423 29596 13491 29652
rect 13547 29596 13615 29652
rect 13671 29596 13739 29652
rect 13795 29596 13863 29652
rect 13919 29596 13987 29652
rect 14043 29596 14111 29652
rect 14167 29596 14235 29652
rect 14291 29596 14359 29652
rect 14415 29596 14483 29652
rect 14539 29596 14607 29652
rect 14663 29596 14673 29652
rect 12861 29528 14673 29596
rect 12861 29472 12871 29528
rect 12927 29472 12995 29528
rect 13051 29472 13119 29528
rect 13175 29472 13243 29528
rect 13299 29472 13367 29528
rect 13423 29472 13491 29528
rect 13547 29472 13615 29528
rect 13671 29472 13739 29528
rect 13795 29472 13863 29528
rect 13919 29472 13987 29528
rect 14043 29472 14111 29528
rect 14167 29472 14235 29528
rect 14291 29472 14359 29528
rect 14415 29472 14483 29528
rect 14539 29472 14607 29528
rect 14663 29472 14673 29528
rect 12861 29404 14673 29472
rect 12861 29348 12871 29404
rect 12927 29348 12995 29404
rect 13051 29348 13119 29404
rect 13175 29348 13243 29404
rect 13299 29348 13367 29404
rect 13423 29348 13491 29404
rect 13547 29348 13615 29404
rect 13671 29348 13739 29404
rect 13795 29348 13863 29404
rect 13919 29348 13987 29404
rect 14043 29348 14111 29404
rect 14167 29348 14235 29404
rect 14291 29348 14359 29404
rect 14415 29348 14483 29404
rect 14539 29348 14607 29404
rect 14663 29348 14673 29404
rect 12861 29280 14673 29348
rect 12861 29224 12871 29280
rect 12927 29224 12995 29280
rect 13051 29224 13119 29280
rect 13175 29224 13243 29280
rect 13299 29224 13367 29280
rect 13423 29224 13491 29280
rect 13547 29224 13615 29280
rect 13671 29224 13739 29280
rect 13795 29224 13863 29280
rect 13919 29224 13987 29280
rect 14043 29224 14111 29280
rect 14167 29224 14235 29280
rect 14291 29224 14359 29280
rect 14415 29224 14483 29280
rect 14539 29224 14607 29280
rect 14663 29224 14673 29280
rect 12861 29156 14673 29224
rect 12861 29100 12871 29156
rect 12927 29100 12995 29156
rect 13051 29100 13119 29156
rect 13175 29100 13243 29156
rect 13299 29100 13367 29156
rect 13423 29100 13491 29156
rect 13547 29100 13615 29156
rect 13671 29100 13739 29156
rect 13795 29100 13863 29156
rect 13919 29100 13987 29156
rect 14043 29100 14111 29156
rect 14167 29100 14235 29156
rect 14291 29100 14359 29156
rect 14415 29100 14483 29156
rect 14539 29100 14607 29156
rect 14663 29100 14673 29156
rect 12861 29032 14673 29100
rect 12861 28976 12871 29032
rect 12927 28976 12995 29032
rect 13051 28976 13119 29032
rect 13175 28976 13243 29032
rect 13299 28976 13367 29032
rect 13423 28976 13491 29032
rect 13547 28976 13615 29032
rect 13671 28976 13739 29032
rect 13795 28976 13863 29032
rect 13919 28976 13987 29032
rect 14043 28976 14111 29032
rect 14167 28976 14235 29032
rect 14291 28976 14359 29032
rect 14415 28976 14483 29032
rect 14539 28976 14607 29032
rect 14663 28976 14673 29032
rect 12861 28908 14673 28976
rect 12861 28852 12871 28908
rect 12927 28852 12995 28908
rect 13051 28852 13119 28908
rect 13175 28852 13243 28908
rect 13299 28852 13367 28908
rect 13423 28852 13491 28908
rect 13547 28852 13615 28908
rect 13671 28852 13739 28908
rect 13795 28852 13863 28908
rect 13919 28852 13987 28908
rect 14043 28852 14111 28908
rect 14167 28852 14235 28908
rect 14291 28852 14359 28908
rect 14415 28852 14483 28908
rect 14539 28852 14607 28908
rect 14663 28852 14673 28908
rect 12861 28842 14673 28852
rect 2481 28548 2681 28558
rect 2481 28492 2491 28548
rect 2547 28492 2615 28548
rect 2671 28492 2681 28548
rect 2481 28424 2681 28492
rect 2481 28368 2491 28424
rect 2547 28368 2615 28424
rect 2671 28368 2681 28424
rect 2481 28300 2681 28368
rect 2481 28244 2491 28300
rect 2547 28244 2615 28300
rect 2671 28244 2681 28300
rect 2481 28176 2681 28244
rect 2481 28120 2491 28176
rect 2547 28120 2615 28176
rect 2671 28120 2681 28176
rect 2481 28052 2681 28120
rect 2481 27996 2491 28052
rect 2547 27996 2615 28052
rect 2671 27996 2681 28052
rect 2481 27928 2681 27996
rect 2481 27872 2491 27928
rect 2547 27872 2615 27928
rect 2671 27872 2681 27928
rect 2481 27804 2681 27872
rect 2481 27748 2491 27804
rect 2547 27748 2615 27804
rect 2671 27748 2681 27804
rect 2481 27680 2681 27748
rect 2481 27624 2491 27680
rect 2547 27624 2615 27680
rect 2671 27624 2681 27680
rect 2481 27556 2681 27624
rect 2481 27500 2491 27556
rect 2547 27500 2615 27556
rect 2671 27500 2681 27556
rect 2481 27432 2681 27500
rect 2481 27376 2491 27432
rect 2547 27376 2615 27432
rect 2671 27376 2681 27432
rect 2481 27308 2681 27376
rect 2481 27252 2491 27308
rect 2547 27252 2615 27308
rect 2671 27252 2681 27308
rect 2481 27242 2681 27252
rect 4851 28548 5051 28558
rect 4851 28492 4861 28548
rect 4917 28492 4985 28548
rect 5041 28492 5051 28548
rect 4851 28424 5051 28492
rect 4851 28368 4861 28424
rect 4917 28368 4985 28424
rect 5041 28368 5051 28424
rect 4851 28300 5051 28368
rect 4851 28244 4861 28300
rect 4917 28244 4985 28300
rect 5041 28244 5051 28300
rect 4851 28176 5051 28244
rect 4851 28120 4861 28176
rect 4917 28120 4985 28176
rect 5041 28120 5051 28176
rect 4851 28052 5051 28120
rect 4851 27996 4861 28052
rect 4917 27996 4985 28052
rect 5041 27996 5051 28052
rect 4851 27928 5051 27996
rect 4851 27872 4861 27928
rect 4917 27872 4985 27928
rect 5041 27872 5051 27928
rect 4851 27804 5051 27872
rect 4851 27748 4861 27804
rect 4917 27748 4985 27804
rect 5041 27748 5051 27804
rect 4851 27680 5051 27748
rect 4851 27624 4861 27680
rect 4917 27624 4985 27680
rect 5041 27624 5051 27680
rect 4851 27556 5051 27624
rect 4851 27500 4861 27556
rect 4917 27500 4985 27556
rect 5041 27500 5051 27556
rect 4851 27432 5051 27500
rect 4851 27376 4861 27432
rect 4917 27376 4985 27432
rect 5041 27376 5051 27432
rect 4851 27308 5051 27376
rect 4851 27252 4861 27308
rect 4917 27252 4985 27308
rect 5041 27252 5051 27308
rect 4851 27242 5051 27252
rect 7265 28548 7713 28558
rect 7265 28492 7275 28548
rect 7331 28492 7399 28548
rect 7455 28492 7523 28548
rect 7579 28492 7647 28548
rect 7703 28492 7713 28548
rect 7265 28424 7713 28492
rect 7265 28368 7275 28424
rect 7331 28368 7399 28424
rect 7455 28368 7523 28424
rect 7579 28368 7647 28424
rect 7703 28368 7713 28424
rect 7265 28300 7713 28368
rect 7265 28244 7275 28300
rect 7331 28244 7399 28300
rect 7455 28244 7523 28300
rect 7579 28244 7647 28300
rect 7703 28244 7713 28300
rect 7265 28176 7713 28244
rect 7265 28120 7275 28176
rect 7331 28120 7399 28176
rect 7455 28120 7523 28176
rect 7579 28120 7647 28176
rect 7703 28120 7713 28176
rect 7265 28052 7713 28120
rect 7265 27996 7275 28052
rect 7331 27996 7399 28052
rect 7455 27996 7523 28052
rect 7579 27996 7647 28052
rect 7703 27996 7713 28052
rect 7265 27928 7713 27996
rect 7265 27872 7275 27928
rect 7331 27872 7399 27928
rect 7455 27872 7523 27928
rect 7579 27872 7647 27928
rect 7703 27872 7713 27928
rect 7265 27804 7713 27872
rect 7265 27748 7275 27804
rect 7331 27748 7399 27804
rect 7455 27748 7523 27804
rect 7579 27748 7647 27804
rect 7703 27748 7713 27804
rect 7265 27680 7713 27748
rect 7265 27624 7275 27680
rect 7331 27624 7399 27680
rect 7455 27624 7523 27680
rect 7579 27624 7647 27680
rect 7703 27624 7713 27680
rect 7265 27556 7713 27624
rect 7265 27500 7275 27556
rect 7331 27500 7399 27556
rect 7455 27500 7523 27556
rect 7579 27500 7647 27556
rect 7703 27500 7713 27556
rect 7265 27432 7713 27500
rect 7265 27376 7275 27432
rect 7331 27376 7399 27432
rect 7455 27376 7523 27432
rect 7579 27376 7647 27432
rect 7703 27376 7713 27432
rect 7265 27308 7713 27376
rect 7265 27252 7275 27308
rect 7331 27252 7399 27308
rect 7455 27252 7523 27308
rect 7579 27252 7647 27308
rect 7703 27252 7713 27308
rect 7265 27242 7713 27252
rect 9927 28548 10127 28558
rect 9927 28492 9937 28548
rect 9993 28492 10061 28548
rect 10117 28492 10127 28548
rect 9927 28424 10127 28492
rect 9927 28368 9937 28424
rect 9993 28368 10061 28424
rect 10117 28368 10127 28424
rect 9927 28300 10127 28368
rect 9927 28244 9937 28300
rect 9993 28244 10061 28300
rect 10117 28244 10127 28300
rect 9927 28176 10127 28244
rect 9927 28120 9937 28176
rect 9993 28120 10061 28176
rect 10117 28120 10127 28176
rect 9927 28052 10127 28120
rect 9927 27996 9937 28052
rect 9993 27996 10061 28052
rect 10117 27996 10127 28052
rect 9927 27928 10127 27996
rect 9927 27872 9937 27928
rect 9993 27872 10061 27928
rect 10117 27872 10127 27928
rect 9927 27804 10127 27872
rect 9927 27748 9937 27804
rect 9993 27748 10061 27804
rect 10117 27748 10127 27804
rect 9927 27680 10127 27748
rect 9927 27624 9937 27680
rect 9993 27624 10061 27680
rect 10117 27624 10127 27680
rect 9927 27556 10127 27624
rect 9927 27500 9937 27556
rect 9993 27500 10061 27556
rect 10117 27500 10127 27556
rect 9927 27432 10127 27500
rect 9927 27376 9937 27432
rect 9993 27376 10061 27432
rect 10117 27376 10127 27432
rect 9927 27308 10127 27376
rect 9927 27252 9937 27308
rect 9993 27252 10061 27308
rect 10117 27252 10127 27308
rect 9927 27242 10127 27252
rect 12297 28548 12497 28558
rect 12297 28492 12307 28548
rect 12363 28492 12431 28548
rect 12487 28492 12497 28548
rect 12297 28424 12497 28492
rect 12297 28368 12307 28424
rect 12363 28368 12431 28424
rect 12487 28368 12497 28424
rect 12297 28300 12497 28368
rect 12297 28244 12307 28300
rect 12363 28244 12431 28300
rect 12487 28244 12497 28300
rect 12297 28176 12497 28244
rect 12297 28120 12307 28176
rect 12363 28120 12431 28176
rect 12487 28120 12497 28176
rect 12297 28052 12497 28120
rect 12297 27996 12307 28052
rect 12363 27996 12431 28052
rect 12487 27996 12497 28052
rect 12297 27928 12497 27996
rect 12297 27872 12307 27928
rect 12363 27872 12431 27928
rect 12487 27872 12497 27928
rect 12297 27804 12497 27872
rect 12297 27748 12307 27804
rect 12363 27748 12431 27804
rect 12487 27748 12497 27804
rect 12297 27680 12497 27748
rect 12297 27624 12307 27680
rect 12363 27624 12431 27680
rect 12487 27624 12497 27680
rect 12297 27556 12497 27624
rect 12297 27500 12307 27556
rect 12363 27500 12431 27556
rect 12487 27500 12497 27556
rect 12297 27432 12497 27500
rect 12297 27376 12307 27432
rect 12363 27376 12431 27432
rect 12487 27376 12497 27432
rect 12297 27308 12497 27376
rect 12297 27252 12307 27308
rect 12363 27252 12431 27308
rect 12487 27252 12497 27308
rect 12297 27242 12497 27252
rect 305 26954 2117 26964
rect 305 26898 315 26954
rect 371 26898 439 26954
rect 495 26898 563 26954
rect 619 26898 687 26954
rect 743 26898 811 26954
rect 867 26898 935 26954
rect 991 26898 1059 26954
rect 1115 26898 1183 26954
rect 1239 26898 1307 26954
rect 1363 26898 1431 26954
rect 1487 26898 1555 26954
rect 1611 26898 1679 26954
rect 1735 26898 1803 26954
rect 1859 26898 1927 26954
rect 1983 26898 2051 26954
rect 2107 26898 2117 26954
rect 305 26830 2117 26898
rect 305 26774 315 26830
rect 371 26774 439 26830
rect 495 26774 563 26830
rect 619 26774 687 26830
rect 743 26774 811 26830
rect 867 26774 935 26830
rect 991 26774 1059 26830
rect 1115 26774 1183 26830
rect 1239 26774 1307 26830
rect 1363 26774 1431 26830
rect 1487 26774 1555 26830
rect 1611 26774 1679 26830
rect 1735 26774 1803 26830
rect 1859 26774 1927 26830
rect 1983 26774 2051 26830
rect 2107 26774 2117 26830
rect 305 26706 2117 26774
rect 305 26650 315 26706
rect 371 26650 439 26706
rect 495 26650 563 26706
rect 619 26650 687 26706
rect 743 26650 811 26706
rect 867 26650 935 26706
rect 991 26650 1059 26706
rect 1115 26650 1183 26706
rect 1239 26650 1307 26706
rect 1363 26650 1431 26706
rect 1487 26650 1555 26706
rect 1611 26650 1679 26706
rect 1735 26650 1803 26706
rect 1859 26650 1927 26706
rect 1983 26650 2051 26706
rect 2107 26650 2117 26706
rect 305 26582 2117 26650
rect 305 26526 315 26582
rect 371 26526 439 26582
rect 495 26526 563 26582
rect 619 26526 687 26582
rect 743 26526 811 26582
rect 867 26526 935 26582
rect 991 26526 1059 26582
rect 1115 26526 1183 26582
rect 1239 26526 1307 26582
rect 1363 26526 1431 26582
rect 1487 26526 1555 26582
rect 1611 26526 1679 26582
rect 1735 26526 1803 26582
rect 1859 26526 1927 26582
rect 1983 26526 2051 26582
rect 2107 26526 2117 26582
rect 305 26458 2117 26526
rect 305 26402 315 26458
rect 371 26402 439 26458
rect 495 26402 563 26458
rect 619 26402 687 26458
rect 743 26402 811 26458
rect 867 26402 935 26458
rect 991 26402 1059 26458
rect 1115 26402 1183 26458
rect 1239 26402 1307 26458
rect 1363 26402 1431 26458
rect 1487 26402 1555 26458
rect 1611 26402 1679 26458
rect 1735 26402 1803 26458
rect 1859 26402 1927 26458
rect 1983 26402 2051 26458
rect 2107 26402 2117 26458
rect 305 26334 2117 26402
rect 305 26278 315 26334
rect 371 26278 439 26334
rect 495 26278 563 26334
rect 619 26278 687 26334
rect 743 26278 811 26334
rect 867 26278 935 26334
rect 991 26278 1059 26334
rect 1115 26278 1183 26334
rect 1239 26278 1307 26334
rect 1363 26278 1431 26334
rect 1487 26278 1555 26334
rect 1611 26278 1679 26334
rect 1735 26278 1803 26334
rect 1859 26278 1927 26334
rect 1983 26278 2051 26334
rect 2107 26278 2117 26334
rect 305 26210 2117 26278
rect 305 26154 315 26210
rect 371 26154 439 26210
rect 495 26154 563 26210
rect 619 26154 687 26210
rect 743 26154 811 26210
rect 867 26154 935 26210
rect 991 26154 1059 26210
rect 1115 26154 1183 26210
rect 1239 26154 1307 26210
rect 1363 26154 1431 26210
rect 1487 26154 1555 26210
rect 1611 26154 1679 26210
rect 1735 26154 1803 26210
rect 1859 26154 1927 26210
rect 1983 26154 2051 26210
rect 2107 26154 2117 26210
rect 305 26086 2117 26154
rect 305 26030 315 26086
rect 371 26030 439 26086
rect 495 26030 563 26086
rect 619 26030 687 26086
rect 743 26030 811 26086
rect 867 26030 935 26086
rect 991 26030 1059 26086
rect 1115 26030 1183 26086
rect 1239 26030 1307 26086
rect 1363 26030 1431 26086
rect 1487 26030 1555 26086
rect 1611 26030 1679 26086
rect 1735 26030 1803 26086
rect 1859 26030 1927 26086
rect 1983 26030 2051 26086
rect 2107 26030 2117 26086
rect 305 25962 2117 26030
rect 305 25906 315 25962
rect 371 25906 439 25962
rect 495 25906 563 25962
rect 619 25906 687 25962
rect 743 25906 811 25962
rect 867 25906 935 25962
rect 991 25906 1059 25962
rect 1115 25906 1183 25962
rect 1239 25906 1307 25962
rect 1363 25906 1431 25962
rect 1487 25906 1555 25962
rect 1611 25906 1679 25962
rect 1735 25906 1803 25962
rect 1859 25906 1927 25962
rect 1983 25906 2051 25962
rect 2107 25906 2117 25962
rect 305 25838 2117 25906
rect 305 25782 315 25838
rect 371 25782 439 25838
rect 495 25782 563 25838
rect 619 25782 687 25838
rect 743 25782 811 25838
rect 867 25782 935 25838
rect 991 25782 1059 25838
rect 1115 25782 1183 25838
rect 1239 25782 1307 25838
rect 1363 25782 1431 25838
rect 1487 25782 1555 25838
rect 1611 25782 1679 25838
rect 1735 25782 1803 25838
rect 1859 25782 1927 25838
rect 1983 25782 2051 25838
rect 2107 25782 2117 25838
rect 305 25714 2117 25782
rect 305 25658 315 25714
rect 371 25658 439 25714
rect 495 25658 563 25714
rect 619 25658 687 25714
rect 743 25658 811 25714
rect 867 25658 935 25714
rect 991 25658 1059 25714
rect 1115 25658 1183 25714
rect 1239 25658 1307 25714
rect 1363 25658 1431 25714
rect 1487 25658 1555 25714
rect 1611 25658 1679 25714
rect 1735 25658 1803 25714
rect 1859 25658 1927 25714
rect 1983 25658 2051 25714
rect 2107 25658 2117 25714
rect 305 25590 2117 25658
rect 305 25534 315 25590
rect 371 25534 439 25590
rect 495 25534 563 25590
rect 619 25534 687 25590
rect 743 25534 811 25590
rect 867 25534 935 25590
rect 991 25534 1059 25590
rect 1115 25534 1183 25590
rect 1239 25534 1307 25590
rect 1363 25534 1431 25590
rect 1487 25534 1555 25590
rect 1611 25534 1679 25590
rect 1735 25534 1803 25590
rect 1859 25534 1927 25590
rect 1983 25534 2051 25590
rect 2107 25534 2117 25590
rect 305 25466 2117 25534
rect 305 25410 315 25466
rect 371 25410 439 25466
rect 495 25410 563 25466
rect 619 25410 687 25466
rect 743 25410 811 25466
rect 867 25410 935 25466
rect 991 25410 1059 25466
rect 1115 25410 1183 25466
rect 1239 25410 1307 25466
rect 1363 25410 1431 25466
rect 1487 25410 1555 25466
rect 1611 25410 1679 25466
rect 1735 25410 1803 25466
rect 1859 25410 1927 25466
rect 1983 25410 2051 25466
rect 2107 25410 2117 25466
rect 305 25342 2117 25410
rect 305 25286 315 25342
rect 371 25286 439 25342
rect 495 25286 563 25342
rect 619 25286 687 25342
rect 743 25286 811 25342
rect 867 25286 935 25342
rect 991 25286 1059 25342
rect 1115 25286 1183 25342
rect 1239 25286 1307 25342
rect 1363 25286 1431 25342
rect 1487 25286 1555 25342
rect 1611 25286 1679 25342
rect 1735 25286 1803 25342
rect 1859 25286 1927 25342
rect 1983 25286 2051 25342
rect 2107 25286 2117 25342
rect 305 25218 2117 25286
rect 305 25162 315 25218
rect 371 25162 439 25218
rect 495 25162 563 25218
rect 619 25162 687 25218
rect 743 25162 811 25218
rect 867 25162 935 25218
rect 991 25162 1059 25218
rect 1115 25162 1183 25218
rect 1239 25162 1307 25218
rect 1363 25162 1431 25218
rect 1487 25162 1555 25218
rect 1611 25162 1679 25218
rect 1735 25162 1803 25218
rect 1859 25162 1927 25218
rect 1983 25162 2051 25218
rect 2107 25162 2117 25218
rect 305 25094 2117 25162
rect 305 25038 315 25094
rect 371 25038 439 25094
rect 495 25038 563 25094
rect 619 25038 687 25094
rect 743 25038 811 25094
rect 867 25038 935 25094
rect 991 25038 1059 25094
rect 1115 25038 1183 25094
rect 1239 25038 1307 25094
rect 1363 25038 1431 25094
rect 1487 25038 1555 25094
rect 1611 25038 1679 25094
rect 1735 25038 1803 25094
rect 1859 25038 1927 25094
rect 1983 25038 2051 25094
rect 2107 25038 2117 25094
rect 305 24970 2117 25038
rect 305 24914 315 24970
rect 371 24914 439 24970
rect 495 24914 563 24970
rect 619 24914 687 24970
rect 743 24914 811 24970
rect 867 24914 935 24970
rect 991 24914 1059 24970
rect 1115 24914 1183 24970
rect 1239 24914 1307 24970
rect 1363 24914 1431 24970
rect 1487 24914 1555 24970
rect 1611 24914 1679 24970
rect 1735 24914 1803 24970
rect 1859 24914 1927 24970
rect 1983 24914 2051 24970
rect 2107 24914 2117 24970
rect 305 24846 2117 24914
rect 305 24790 315 24846
rect 371 24790 439 24846
rect 495 24790 563 24846
rect 619 24790 687 24846
rect 743 24790 811 24846
rect 867 24790 935 24846
rect 991 24790 1059 24846
rect 1115 24790 1183 24846
rect 1239 24790 1307 24846
rect 1363 24790 1431 24846
rect 1487 24790 1555 24846
rect 1611 24790 1679 24846
rect 1735 24790 1803 24846
rect 1859 24790 1927 24846
rect 1983 24790 2051 24846
rect 2107 24790 2117 24846
rect 305 24722 2117 24790
rect 305 24666 315 24722
rect 371 24666 439 24722
rect 495 24666 563 24722
rect 619 24666 687 24722
rect 743 24666 811 24722
rect 867 24666 935 24722
rect 991 24666 1059 24722
rect 1115 24666 1183 24722
rect 1239 24666 1307 24722
rect 1363 24666 1431 24722
rect 1487 24666 1555 24722
rect 1611 24666 1679 24722
rect 1735 24666 1803 24722
rect 1859 24666 1927 24722
rect 1983 24666 2051 24722
rect 2107 24666 2117 24722
rect 305 24598 2117 24666
rect 305 24542 315 24598
rect 371 24542 439 24598
rect 495 24542 563 24598
rect 619 24542 687 24598
rect 743 24542 811 24598
rect 867 24542 935 24598
rect 991 24542 1059 24598
rect 1115 24542 1183 24598
rect 1239 24542 1307 24598
rect 1363 24542 1431 24598
rect 1487 24542 1555 24598
rect 1611 24542 1679 24598
rect 1735 24542 1803 24598
rect 1859 24542 1927 24598
rect 1983 24542 2051 24598
rect 2107 24542 2117 24598
rect 305 24474 2117 24542
rect 305 24418 315 24474
rect 371 24418 439 24474
rect 495 24418 563 24474
rect 619 24418 687 24474
rect 743 24418 811 24474
rect 867 24418 935 24474
rect 991 24418 1059 24474
rect 1115 24418 1183 24474
rect 1239 24418 1307 24474
rect 1363 24418 1431 24474
rect 1487 24418 1555 24474
rect 1611 24418 1679 24474
rect 1735 24418 1803 24474
rect 1859 24418 1927 24474
rect 1983 24418 2051 24474
rect 2107 24418 2117 24474
rect 305 24350 2117 24418
rect 305 24294 315 24350
rect 371 24294 439 24350
rect 495 24294 563 24350
rect 619 24294 687 24350
rect 743 24294 811 24350
rect 867 24294 935 24350
rect 991 24294 1059 24350
rect 1115 24294 1183 24350
rect 1239 24294 1307 24350
rect 1363 24294 1431 24350
rect 1487 24294 1555 24350
rect 1611 24294 1679 24350
rect 1735 24294 1803 24350
rect 1859 24294 1927 24350
rect 1983 24294 2051 24350
rect 2107 24294 2117 24350
rect 305 24226 2117 24294
rect 305 24170 315 24226
rect 371 24170 439 24226
rect 495 24170 563 24226
rect 619 24170 687 24226
rect 743 24170 811 24226
rect 867 24170 935 24226
rect 991 24170 1059 24226
rect 1115 24170 1183 24226
rect 1239 24170 1307 24226
rect 1363 24170 1431 24226
rect 1487 24170 1555 24226
rect 1611 24170 1679 24226
rect 1735 24170 1803 24226
rect 1859 24170 1927 24226
rect 1983 24170 2051 24226
rect 2107 24170 2117 24226
rect 305 24102 2117 24170
rect 305 24046 315 24102
rect 371 24046 439 24102
rect 495 24046 563 24102
rect 619 24046 687 24102
rect 743 24046 811 24102
rect 867 24046 935 24102
rect 991 24046 1059 24102
rect 1115 24046 1183 24102
rect 1239 24046 1307 24102
rect 1363 24046 1431 24102
rect 1487 24046 1555 24102
rect 1611 24046 1679 24102
rect 1735 24046 1803 24102
rect 1859 24046 1927 24102
rect 1983 24046 2051 24102
rect 2107 24046 2117 24102
rect 305 24036 2117 24046
rect 2798 26954 4734 26964
rect 2798 26898 2808 26954
rect 2864 26898 2932 26954
rect 2988 26898 3056 26954
rect 3112 26898 3180 26954
rect 3236 26898 3304 26954
rect 3360 26898 3428 26954
rect 3484 26898 3552 26954
rect 3608 26898 3676 26954
rect 3732 26898 3800 26954
rect 3856 26898 3924 26954
rect 3980 26898 4048 26954
rect 4104 26898 4172 26954
rect 4228 26898 4296 26954
rect 4352 26898 4420 26954
rect 4476 26898 4544 26954
rect 4600 26898 4668 26954
rect 4724 26898 4734 26954
rect 2798 26830 4734 26898
rect 2798 26774 2808 26830
rect 2864 26774 2932 26830
rect 2988 26774 3056 26830
rect 3112 26774 3180 26830
rect 3236 26774 3304 26830
rect 3360 26774 3428 26830
rect 3484 26774 3552 26830
rect 3608 26774 3676 26830
rect 3732 26774 3800 26830
rect 3856 26774 3924 26830
rect 3980 26774 4048 26830
rect 4104 26774 4172 26830
rect 4228 26774 4296 26830
rect 4352 26774 4420 26830
rect 4476 26774 4544 26830
rect 4600 26774 4668 26830
rect 4724 26774 4734 26830
rect 2798 26706 4734 26774
rect 2798 26650 2808 26706
rect 2864 26650 2932 26706
rect 2988 26650 3056 26706
rect 3112 26650 3180 26706
rect 3236 26650 3304 26706
rect 3360 26650 3428 26706
rect 3484 26650 3552 26706
rect 3608 26650 3676 26706
rect 3732 26650 3800 26706
rect 3856 26650 3924 26706
rect 3980 26650 4048 26706
rect 4104 26650 4172 26706
rect 4228 26650 4296 26706
rect 4352 26650 4420 26706
rect 4476 26650 4544 26706
rect 4600 26650 4668 26706
rect 4724 26650 4734 26706
rect 2798 26582 4734 26650
rect 2798 26526 2808 26582
rect 2864 26526 2932 26582
rect 2988 26526 3056 26582
rect 3112 26526 3180 26582
rect 3236 26526 3304 26582
rect 3360 26526 3428 26582
rect 3484 26526 3552 26582
rect 3608 26526 3676 26582
rect 3732 26526 3800 26582
rect 3856 26526 3924 26582
rect 3980 26526 4048 26582
rect 4104 26526 4172 26582
rect 4228 26526 4296 26582
rect 4352 26526 4420 26582
rect 4476 26526 4544 26582
rect 4600 26526 4668 26582
rect 4724 26526 4734 26582
rect 2798 26458 4734 26526
rect 2798 26402 2808 26458
rect 2864 26402 2932 26458
rect 2988 26402 3056 26458
rect 3112 26402 3180 26458
rect 3236 26402 3304 26458
rect 3360 26402 3428 26458
rect 3484 26402 3552 26458
rect 3608 26402 3676 26458
rect 3732 26402 3800 26458
rect 3856 26402 3924 26458
rect 3980 26402 4048 26458
rect 4104 26402 4172 26458
rect 4228 26402 4296 26458
rect 4352 26402 4420 26458
rect 4476 26402 4544 26458
rect 4600 26402 4668 26458
rect 4724 26402 4734 26458
rect 2798 26334 4734 26402
rect 2798 26278 2808 26334
rect 2864 26278 2932 26334
rect 2988 26278 3056 26334
rect 3112 26278 3180 26334
rect 3236 26278 3304 26334
rect 3360 26278 3428 26334
rect 3484 26278 3552 26334
rect 3608 26278 3676 26334
rect 3732 26278 3800 26334
rect 3856 26278 3924 26334
rect 3980 26278 4048 26334
rect 4104 26278 4172 26334
rect 4228 26278 4296 26334
rect 4352 26278 4420 26334
rect 4476 26278 4544 26334
rect 4600 26278 4668 26334
rect 4724 26278 4734 26334
rect 2798 26210 4734 26278
rect 2798 26154 2808 26210
rect 2864 26154 2932 26210
rect 2988 26154 3056 26210
rect 3112 26154 3180 26210
rect 3236 26154 3304 26210
rect 3360 26154 3428 26210
rect 3484 26154 3552 26210
rect 3608 26154 3676 26210
rect 3732 26154 3800 26210
rect 3856 26154 3924 26210
rect 3980 26154 4048 26210
rect 4104 26154 4172 26210
rect 4228 26154 4296 26210
rect 4352 26154 4420 26210
rect 4476 26154 4544 26210
rect 4600 26154 4668 26210
rect 4724 26154 4734 26210
rect 2798 26086 4734 26154
rect 2798 26030 2808 26086
rect 2864 26030 2932 26086
rect 2988 26030 3056 26086
rect 3112 26030 3180 26086
rect 3236 26030 3304 26086
rect 3360 26030 3428 26086
rect 3484 26030 3552 26086
rect 3608 26030 3676 26086
rect 3732 26030 3800 26086
rect 3856 26030 3924 26086
rect 3980 26030 4048 26086
rect 4104 26030 4172 26086
rect 4228 26030 4296 26086
rect 4352 26030 4420 26086
rect 4476 26030 4544 26086
rect 4600 26030 4668 26086
rect 4724 26030 4734 26086
rect 2798 25962 4734 26030
rect 2798 25906 2808 25962
rect 2864 25906 2932 25962
rect 2988 25906 3056 25962
rect 3112 25906 3180 25962
rect 3236 25906 3304 25962
rect 3360 25906 3428 25962
rect 3484 25906 3552 25962
rect 3608 25906 3676 25962
rect 3732 25906 3800 25962
rect 3856 25906 3924 25962
rect 3980 25906 4048 25962
rect 4104 25906 4172 25962
rect 4228 25906 4296 25962
rect 4352 25906 4420 25962
rect 4476 25906 4544 25962
rect 4600 25906 4668 25962
rect 4724 25906 4734 25962
rect 2798 25838 4734 25906
rect 2798 25782 2808 25838
rect 2864 25782 2932 25838
rect 2988 25782 3056 25838
rect 3112 25782 3180 25838
rect 3236 25782 3304 25838
rect 3360 25782 3428 25838
rect 3484 25782 3552 25838
rect 3608 25782 3676 25838
rect 3732 25782 3800 25838
rect 3856 25782 3924 25838
rect 3980 25782 4048 25838
rect 4104 25782 4172 25838
rect 4228 25782 4296 25838
rect 4352 25782 4420 25838
rect 4476 25782 4544 25838
rect 4600 25782 4668 25838
rect 4724 25782 4734 25838
rect 2798 25714 4734 25782
rect 2798 25658 2808 25714
rect 2864 25658 2932 25714
rect 2988 25658 3056 25714
rect 3112 25658 3180 25714
rect 3236 25658 3304 25714
rect 3360 25658 3428 25714
rect 3484 25658 3552 25714
rect 3608 25658 3676 25714
rect 3732 25658 3800 25714
rect 3856 25658 3924 25714
rect 3980 25658 4048 25714
rect 4104 25658 4172 25714
rect 4228 25658 4296 25714
rect 4352 25658 4420 25714
rect 4476 25658 4544 25714
rect 4600 25658 4668 25714
rect 4724 25658 4734 25714
rect 2798 25590 4734 25658
rect 2798 25534 2808 25590
rect 2864 25534 2932 25590
rect 2988 25534 3056 25590
rect 3112 25534 3180 25590
rect 3236 25534 3304 25590
rect 3360 25534 3428 25590
rect 3484 25534 3552 25590
rect 3608 25534 3676 25590
rect 3732 25534 3800 25590
rect 3856 25534 3924 25590
rect 3980 25534 4048 25590
rect 4104 25534 4172 25590
rect 4228 25534 4296 25590
rect 4352 25534 4420 25590
rect 4476 25534 4544 25590
rect 4600 25534 4668 25590
rect 4724 25534 4734 25590
rect 2798 25466 4734 25534
rect 2798 25410 2808 25466
rect 2864 25410 2932 25466
rect 2988 25410 3056 25466
rect 3112 25410 3180 25466
rect 3236 25410 3304 25466
rect 3360 25410 3428 25466
rect 3484 25410 3552 25466
rect 3608 25410 3676 25466
rect 3732 25410 3800 25466
rect 3856 25410 3924 25466
rect 3980 25410 4048 25466
rect 4104 25410 4172 25466
rect 4228 25410 4296 25466
rect 4352 25410 4420 25466
rect 4476 25410 4544 25466
rect 4600 25410 4668 25466
rect 4724 25410 4734 25466
rect 2798 25342 4734 25410
rect 2798 25286 2808 25342
rect 2864 25286 2932 25342
rect 2988 25286 3056 25342
rect 3112 25286 3180 25342
rect 3236 25286 3304 25342
rect 3360 25286 3428 25342
rect 3484 25286 3552 25342
rect 3608 25286 3676 25342
rect 3732 25286 3800 25342
rect 3856 25286 3924 25342
rect 3980 25286 4048 25342
rect 4104 25286 4172 25342
rect 4228 25286 4296 25342
rect 4352 25286 4420 25342
rect 4476 25286 4544 25342
rect 4600 25286 4668 25342
rect 4724 25286 4734 25342
rect 2798 25218 4734 25286
rect 2798 25162 2808 25218
rect 2864 25162 2932 25218
rect 2988 25162 3056 25218
rect 3112 25162 3180 25218
rect 3236 25162 3304 25218
rect 3360 25162 3428 25218
rect 3484 25162 3552 25218
rect 3608 25162 3676 25218
rect 3732 25162 3800 25218
rect 3856 25162 3924 25218
rect 3980 25162 4048 25218
rect 4104 25162 4172 25218
rect 4228 25162 4296 25218
rect 4352 25162 4420 25218
rect 4476 25162 4544 25218
rect 4600 25162 4668 25218
rect 4724 25162 4734 25218
rect 2798 25094 4734 25162
rect 2798 25038 2808 25094
rect 2864 25038 2932 25094
rect 2988 25038 3056 25094
rect 3112 25038 3180 25094
rect 3236 25038 3304 25094
rect 3360 25038 3428 25094
rect 3484 25038 3552 25094
rect 3608 25038 3676 25094
rect 3732 25038 3800 25094
rect 3856 25038 3924 25094
rect 3980 25038 4048 25094
rect 4104 25038 4172 25094
rect 4228 25038 4296 25094
rect 4352 25038 4420 25094
rect 4476 25038 4544 25094
rect 4600 25038 4668 25094
rect 4724 25038 4734 25094
rect 2798 24970 4734 25038
rect 2798 24914 2808 24970
rect 2864 24914 2932 24970
rect 2988 24914 3056 24970
rect 3112 24914 3180 24970
rect 3236 24914 3304 24970
rect 3360 24914 3428 24970
rect 3484 24914 3552 24970
rect 3608 24914 3676 24970
rect 3732 24914 3800 24970
rect 3856 24914 3924 24970
rect 3980 24914 4048 24970
rect 4104 24914 4172 24970
rect 4228 24914 4296 24970
rect 4352 24914 4420 24970
rect 4476 24914 4544 24970
rect 4600 24914 4668 24970
rect 4724 24914 4734 24970
rect 2798 24846 4734 24914
rect 2798 24790 2808 24846
rect 2864 24790 2932 24846
rect 2988 24790 3056 24846
rect 3112 24790 3180 24846
rect 3236 24790 3304 24846
rect 3360 24790 3428 24846
rect 3484 24790 3552 24846
rect 3608 24790 3676 24846
rect 3732 24790 3800 24846
rect 3856 24790 3924 24846
rect 3980 24790 4048 24846
rect 4104 24790 4172 24846
rect 4228 24790 4296 24846
rect 4352 24790 4420 24846
rect 4476 24790 4544 24846
rect 4600 24790 4668 24846
rect 4724 24790 4734 24846
rect 2798 24722 4734 24790
rect 2798 24666 2808 24722
rect 2864 24666 2932 24722
rect 2988 24666 3056 24722
rect 3112 24666 3180 24722
rect 3236 24666 3304 24722
rect 3360 24666 3428 24722
rect 3484 24666 3552 24722
rect 3608 24666 3676 24722
rect 3732 24666 3800 24722
rect 3856 24666 3924 24722
rect 3980 24666 4048 24722
rect 4104 24666 4172 24722
rect 4228 24666 4296 24722
rect 4352 24666 4420 24722
rect 4476 24666 4544 24722
rect 4600 24666 4668 24722
rect 4724 24666 4734 24722
rect 2798 24598 4734 24666
rect 2798 24542 2808 24598
rect 2864 24542 2932 24598
rect 2988 24542 3056 24598
rect 3112 24542 3180 24598
rect 3236 24542 3304 24598
rect 3360 24542 3428 24598
rect 3484 24542 3552 24598
rect 3608 24542 3676 24598
rect 3732 24542 3800 24598
rect 3856 24542 3924 24598
rect 3980 24542 4048 24598
rect 4104 24542 4172 24598
rect 4228 24542 4296 24598
rect 4352 24542 4420 24598
rect 4476 24542 4544 24598
rect 4600 24542 4668 24598
rect 4724 24542 4734 24598
rect 2798 24474 4734 24542
rect 2798 24418 2808 24474
rect 2864 24418 2932 24474
rect 2988 24418 3056 24474
rect 3112 24418 3180 24474
rect 3236 24418 3304 24474
rect 3360 24418 3428 24474
rect 3484 24418 3552 24474
rect 3608 24418 3676 24474
rect 3732 24418 3800 24474
rect 3856 24418 3924 24474
rect 3980 24418 4048 24474
rect 4104 24418 4172 24474
rect 4228 24418 4296 24474
rect 4352 24418 4420 24474
rect 4476 24418 4544 24474
rect 4600 24418 4668 24474
rect 4724 24418 4734 24474
rect 2798 24350 4734 24418
rect 2798 24294 2808 24350
rect 2864 24294 2932 24350
rect 2988 24294 3056 24350
rect 3112 24294 3180 24350
rect 3236 24294 3304 24350
rect 3360 24294 3428 24350
rect 3484 24294 3552 24350
rect 3608 24294 3676 24350
rect 3732 24294 3800 24350
rect 3856 24294 3924 24350
rect 3980 24294 4048 24350
rect 4104 24294 4172 24350
rect 4228 24294 4296 24350
rect 4352 24294 4420 24350
rect 4476 24294 4544 24350
rect 4600 24294 4668 24350
rect 4724 24294 4734 24350
rect 2798 24226 4734 24294
rect 2798 24170 2808 24226
rect 2864 24170 2932 24226
rect 2988 24170 3056 24226
rect 3112 24170 3180 24226
rect 3236 24170 3304 24226
rect 3360 24170 3428 24226
rect 3484 24170 3552 24226
rect 3608 24170 3676 24226
rect 3732 24170 3800 24226
rect 3856 24170 3924 24226
rect 3980 24170 4048 24226
rect 4104 24170 4172 24226
rect 4228 24170 4296 24226
rect 4352 24170 4420 24226
rect 4476 24170 4544 24226
rect 4600 24170 4668 24226
rect 4724 24170 4734 24226
rect 2798 24102 4734 24170
rect 2798 24046 2808 24102
rect 2864 24046 2932 24102
rect 2988 24046 3056 24102
rect 3112 24046 3180 24102
rect 3236 24046 3304 24102
rect 3360 24046 3428 24102
rect 3484 24046 3552 24102
rect 3608 24046 3676 24102
rect 3732 24046 3800 24102
rect 3856 24046 3924 24102
rect 3980 24046 4048 24102
rect 4104 24046 4172 24102
rect 4228 24046 4296 24102
rect 4352 24046 4420 24102
rect 4476 24046 4544 24102
rect 4600 24046 4668 24102
rect 4724 24046 4734 24102
rect 2798 24036 4734 24046
rect 5168 26954 7104 26964
rect 5168 26898 5178 26954
rect 5234 26898 5302 26954
rect 5358 26898 5426 26954
rect 5482 26898 5550 26954
rect 5606 26898 5674 26954
rect 5730 26898 5798 26954
rect 5854 26898 5922 26954
rect 5978 26898 6046 26954
rect 6102 26898 6170 26954
rect 6226 26898 6294 26954
rect 6350 26898 6418 26954
rect 6474 26898 6542 26954
rect 6598 26898 6666 26954
rect 6722 26898 6790 26954
rect 6846 26898 6914 26954
rect 6970 26898 7038 26954
rect 7094 26898 7104 26954
rect 5168 26830 7104 26898
rect 5168 26774 5178 26830
rect 5234 26774 5302 26830
rect 5358 26774 5426 26830
rect 5482 26774 5550 26830
rect 5606 26774 5674 26830
rect 5730 26774 5798 26830
rect 5854 26774 5922 26830
rect 5978 26774 6046 26830
rect 6102 26774 6170 26830
rect 6226 26774 6294 26830
rect 6350 26774 6418 26830
rect 6474 26774 6542 26830
rect 6598 26774 6666 26830
rect 6722 26774 6790 26830
rect 6846 26774 6914 26830
rect 6970 26774 7038 26830
rect 7094 26774 7104 26830
rect 5168 26706 7104 26774
rect 5168 26650 5178 26706
rect 5234 26650 5302 26706
rect 5358 26650 5426 26706
rect 5482 26650 5550 26706
rect 5606 26650 5674 26706
rect 5730 26650 5798 26706
rect 5854 26650 5922 26706
rect 5978 26650 6046 26706
rect 6102 26650 6170 26706
rect 6226 26650 6294 26706
rect 6350 26650 6418 26706
rect 6474 26650 6542 26706
rect 6598 26650 6666 26706
rect 6722 26650 6790 26706
rect 6846 26650 6914 26706
rect 6970 26650 7038 26706
rect 7094 26650 7104 26706
rect 5168 26582 7104 26650
rect 5168 26526 5178 26582
rect 5234 26526 5302 26582
rect 5358 26526 5426 26582
rect 5482 26526 5550 26582
rect 5606 26526 5674 26582
rect 5730 26526 5798 26582
rect 5854 26526 5922 26582
rect 5978 26526 6046 26582
rect 6102 26526 6170 26582
rect 6226 26526 6294 26582
rect 6350 26526 6418 26582
rect 6474 26526 6542 26582
rect 6598 26526 6666 26582
rect 6722 26526 6790 26582
rect 6846 26526 6914 26582
rect 6970 26526 7038 26582
rect 7094 26526 7104 26582
rect 5168 26458 7104 26526
rect 5168 26402 5178 26458
rect 5234 26402 5302 26458
rect 5358 26402 5426 26458
rect 5482 26402 5550 26458
rect 5606 26402 5674 26458
rect 5730 26402 5798 26458
rect 5854 26402 5922 26458
rect 5978 26402 6046 26458
rect 6102 26402 6170 26458
rect 6226 26402 6294 26458
rect 6350 26402 6418 26458
rect 6474 26402 6542 26458
rect 6598 26402 6666 26458
rect 6722 26402 6790 26458
rect 6846 26402 6914 26458
rect 6970 26402 7038 26458
rect 7094 26402 7104 26458
rect 5168 26334 7104 26402
rect 5168 26278 5178 26334
rect 5234 26278 5302 26334
rect 5358 26278 5426 26334
rect 5482 26278 5550 26334
rect 5606 26278 5674 26334
rect 5730 26278 5798 26334
rect 5854 26278 5922 26334
rect 5978 26278 6046 26334
rect 6102 26278 6170 26334
rect 6226 26278 6294 26334
rect 6350 26278 6418 26334
rect 6474 26278 6542 26334
rect 6598 26278 6666 26334
rect 6722 26278 6790 26334
rect 6846 26278 6914 26334
rect 6970 26278 7038 26334
rect 7094 26278 7104 26334
rect 5168 26210 7104 26278
rect 5168 26154 5178 26210
rect 5234 26154 5302 26210
rect 5358 26154 5426 26210
rect 5482 26154 5550 26210
rect 5606 26154 5674 26210
rect 5730 26154 5798 26210
rect 5854 26154 5922 26210
rect 5978 26154 6046 26210
rect 6102 26154 6170 26210
rect 6226 26154 6294 26210
rect 6350 26154 6418 26210
rect 6474 26154 6542 26210
rect 6598 26154 6666 26210
rect 6722 26154 6790 26210
rect 6846 26154 6914 26210
rect 6970 26154 7038 26210
rect 7094 26154 7104 26210
rect 5168 26086 7104 26154
rect 5168 26030 5178 26086
rect 5234 26030 5302 26086
rect 5358 26030 5426 26086
rect 5482 26030 5550 26086
rect 5606 26030 5674 26086
rect 5730 26030 5798 26086
rect 5854 26030 5922 26086
rect 5978 26030 6046 26086
rect 6102 26030 6170 26086
rect 6226 26030 6294 26086
rect 6350 26030 6418 26086
rect 6474 26030 6542 26086
rect 6598 26030 6666 26086
rect 6722 26030 6790 26086
rect 6846 26030 6914 26086
rect 6970 26030 7038 26086
rect 7094 26030 7104 26086
rect 5168 25962 7104 26030
rect 5168 25906 5178 25962
rect 5234 25906 5302 25962
rect 5358 25906 5426 25962
rect 5482 25906 5550 25962
rect 5606 25906 5674 25962
rect 5730 25906 5798 25962
rect 5854 25906 5922 25962
rect 5978 25906 6046 25962
rect 6102 25906 6170 25962
rect 6226 25906 6294 25962
rect 6350 25906 6418 25962
rect 6474 25906 6542 25962
rect 6598 25906 6666 25962
rect 6722 25906 6790 25962
rect 6846 25906 6914 25962
rect 6970 25906 7038 25962
rect 7094 25906 7104 25962
rect 5168 25838 7104 25906
rect 5168 25782 5178 25838
rect 5234 25782 5302 25838
rect 5358 25782 5426 25838
rect 5482 25782 5550 25838
rect 5606 25782 5674 25838
rect 5730 25782 5798 25838
rect 5854 25782 5922 25838
rect 5978 25782 6046 25838
rect 6102 25782 6170 25838
rect 6226 25782 6294 25838
rect 6350 25782 6418 25838
rect 6474 25782 6542 25838
rect 6598 25782 6666 25838
rect 6722 25782 6790 25838
rect 6846 25782 6914 25838
rect 6970 25782 7038 25838
rect 7094 25782 7104 25838
rect 5168 25714 7104 25782
rect 5168 25658 5178 25714
rect 5234 25658 5302 25714
rect 5358 25658 5426 25714
rect 5482 25658 5550 25714
rect 5606 25658 5674 25714
rect 5730 25658 5798 25714
rect 5854 25658 5922 25714
rect 5978 25658 6046 25714
rect 6102 25658 6170 25714
rect 6226 25658 6294 25714
rect 6350 25658 6418 25714
rect 6474 25658 6542 25714
rect 6598 25658 6666 25714
rect 6722 25658 6790 25714
rect 6846 25658 6914 25714
rect 6970 25658 7038 25714
rect 7094 25658 7104 25714
rect 5168 25590 7104 25658
rect 5168 25534 5178 25590
rect 5234 25534 5302 25590
rect 5358 25534 5426 25590
rect 5482 25534 5550 25590
rect 5606 25534 5674 25590
rect 5730 25534 5798 25590
rect 5854 25534 5922 25590
rect 5978 25534 6046 25590
rect 6102 25534 6170 25590
rect 6226 25534 6294 25590
rect 6350 25534 6418 25590
rect 6474 25534 6542 25590
rect 6598 25534 6666 25590
rect 6722 25534 6790 25590
rect 6846 25534 6914 25590
rect 6970 25534 7038 25590
rect 7094 25534 7104 25590
rect 5168 25466 7104 25534
rect 5168 25410 5178 25466
rect 5234 25410 5302 25466
rect 5358 25410 5426 25466
rect 5482 25410 5550 25466
rect 5606 25410 5674 25466
rect 5730 25410 5798 25466
rect 5854 25410 5922 25466
rect 5978 25410 6046 25466
rect 6102 25410 6170 25466
rect 6226 25410 6294 25466
rect 6350 25410 6418 25466
rect 6474 25410 6542 25466
rect 6598 25410 6666 25466
rect 6722 25410 6790 25466
rect 6846 25410 6914 25466
rect 6970 25410 7038 25466
rect 7094 25410 7104 25466
rect 5168 25342 7104 25410
rect 5168 25286 5178 25342
rect 5234 25286 5302 25342
rect 5358 25286 5426 25342
rect 5482 25286 5550 25342
rect 5606 25286 5674 25342
rect 5730 25286 5798 25342
rect 5854 25286 5922 25342
rect 5978 25286 6046 25342
rect 6102 25286 6170 25342
rect 6226 25286 6294 25342
rect 6350 25286 6418 25342
rect 6474 25286 6542 25342
rect 6598 25286 6666 25342
rect 6722 25286 6790 25342
rect 6846 25286 6914 25342
rect 6970 25286 7038 25342
rect 7094 25286 7104 25342
rect 5168 25218 7104 25286
rect 5168 25162 5178 25218
rect 5234 25162 5302 25218
rect 5358 25162 5426 25218
rect 5482 25162 5550 25218
rect 5606 25162 5674 25218
rect 5730 25162 5798 25218
rect 5854 25162 5922 25218
rect 5978 25162 6046 25218
rect 6102 25162 6170 25218
rect 6226 25162 6294 25218
rect 6350 25162 6418 25218
rect 6474 25162 6542 25218
rect 6598 25162 6666 25218
rect 6722 25162 6790 25218
rect 6846 25162 6914 25218
rect 6970 25162 7038 25218
rect 7094 25162 7104 25218
rect 5168 25094 7104 25162
rect 5168 25038 5178 25094
rect 5234 25038 5302 25094
rect 5358 25038 5426 25094
rect 5482 25038 5550 25094
rect 5606 25038 5674 25094
rect 5730 25038 5798 25094
rect 5854 25038 5922 25094
rect 5978 25038 6046 25094
rect 6102 25038 6170 25094
rect 6226 25038 6294 25094
rect 6350 25038 6418 25094
rect 6474 25038 6542 25094
rect 6598 25038 6666 25094
rect 6722 25038 6790 25094
rect 6846 25038 6914 25094
rect 6970 25038 7038 25094
rect 7094 25038 7104 25094
rect 5168 24970 7104 25038
rect 5168 24914 5178 24970
rect 5234 24914 5302 24970
rect 5358 24914 5426 24970
rect 5482 24914 5550 24970
rect 5606 24914 5674 24970
rect 5730 24914 5798 24970
rect 5854 24914 5922 24970
rect 5978 24914 6046 24970
rect 6102 24914 6170 24970
rect 6226 24914 6294 24970
rect 6350 24914 6418 24970
rect 6474 24914 6542 24970
rect 6598 24914 6666 24970
rect 6722 24914 6790 24970
rect 6846 24914 6914 24970
rect 6970 24914 7038 24970
rect 7094 24914 7104 24970
rect 5168 24846 7104 24914
rect 5168 24790 5178 24846
rect 5234 24790 5302 24846
rect 5358 24790 5426 24846
rect 5482 24790 5550 24846
rect 5606 24790 5674 24846
rect 5730 24790 5798 24846
rect 5854 24790 5922 24846
rect 5978 24790 6046 24846
rect 6102 24790 6170 24846
rect 6226 24790 6294 24846
rect 6350 24790 6418 24846
rect 6474 24790 6542 24846
rect 6598 24790 6666 24846
rect 6722 24790 6790 24846
rect 6846 24790 6914 24846
rect 6970 24790 7038 24846
rect 7094 24790 7104 24846
rect 5168 24722 7104 24790
rect 5168 24666 5178 24722
rect 5234 24666 5302 24722
rect 5358 24666 5426 24722
rect 5482 24666 5550 24722
rect 5606 24666 5674 24722
rect 5730 24666 5798 24722
rect 5854 24666 5922 24722
rect 5978 24666 6046 24722
rect 6102 24666 6170 24722
rect 6226 24666 6294 24722
rect 6350 24666 6418 24722
rect 6474 24666 6542 24722
rect 6598 24666 6666 24722
rect 6722 24666 6790 24722
rect 6846 24666 6914 24722
rect 6970 24666 7038 24722
rect 7094 24666 7104 24722
rect 5168 24598 7104 24666
rect 5168 24542 5178 24598
rect 5234 24542 5302 24598
rect 5358 24542 5426 24598
rect 5482 24542 5550 24598
rect 5606 24542 5674 24598
rect 5730 24542 5798 24598
rect 5854 24542 5922 24598
rect 5978 24542 6046 24598
rect 6102 24542 6170 24598
rect 6226 24542 6294 24598
rect 6350 24542 6418 24598
rect 6474 24542 6542 24598
rect 6598 24542 6666 24598
rect 6722 24542 6790 24598
rect 6846 24542 6914 24598
rect 6970 24542 7038 24598
rect 7094 24542 7104 24598
rect 5168 24474 7104 24542
rect 5168 24418 5178 24474
rect 5234 24418 5302 24474
rect 5358 24418 5426 24474
rect 5482 24418 5550 24474
rect 5606 24418 5674 24474
rect 5730 24418 5798 24474
rect 5854 24418 5922 24474
rect 5978 24418 6046 24474
rect 6102 24418 6170 24474
rect 6226 24418 6294 24474
rect 6350 24418 6418 24474
rect 6474 24418 6542 24474
rect 6598 24418 6666 24474
rect 6722 24418 6790 24474
rect 6846 24418 6914 24474
rect 6970 24418 7038 24474
rect 7094 24418 7104 24474
rect 5168 24350 7104 24418
rect 5168 24294 5178 24350
rect 5234 24294 5302 24350
rect 5358 24294 5426 24350
rect 5482 24294 5550 24350
rect 5606 24294 5674 24350
rect 5730 24294 5798 24350
rect 5854 24294 5922 24350
rect 5978 24294 6046 24350
rect 6102 24294 6170 24350
rect 6226 24294 6294 24350
rect 6350 24294 6418 24350
rect 6474 24294 6542 24350
rect 6598 24294 6666 24350
rect 6722 24294 6790 24350
rect 6846 24294 6914 24350
rect 6970 24294 7038 24350
rect 7094 24294 7104 24350
rect 5168 24226 7104 24294
rect 5168 24170 5178 24226
rect 5234 24170 5302 24226
rect 5358 24170 5426 24226
rect 5482 24170 5550 24226
rect 5606 24170 5674 24226
rect 5730 24170 5798 24226
rect 5854 24170 5922 24226
rect 5978 24170 6046 24226
rect 6102 24170 6170 24226
rect 6226 24170 6294 24226
rect 6350 24170 6418 24226
rect 6474 24170 6542 24226
rect 6598 24170 6666 24226
rect 6722 24170 6790 24226
rect 6846 24170 6914 24226
rect 6970 24170 7038 24226
rect 7094 24170 7104 24226
rect 5168 24102 7104 24170
rect 5168 24046 5178 24102
rect 5234 24046 5302 24102
rect 5358 24046 5426 24102
rect 5482 24046 5550 24102
rect 5606 24046 5674 24102
rect 5730 24046 5798 24102
rect 5854 24046 5922 24102
rect 5978 24046 6046 24102
rect 6102 24046 6170 24102
rect 6226 24046 6294 24102
rect 6350 24046 6418 24102
rect 6474 24046 6542 24102
rect 6598 24046 6666 24102
rect 6722 24046 6790 24102
rect 6846 24046 6914 24102
rect 6970 24046 7038 24102
rect 7094 24046 7104 24102
rect 5168 24036 7104 24046
rect 7874 26954 9810 26964
rect 7874 26898 7884 26954
rect 7940 26898 8008 26954
rect 8064 26898 8132 26954
rect 8188 26898 8256 26954
rect 8312 26898 8380 26954
rect 8436 26898 8504 26954
rect 8560 26898 8628 26954
rect 8684 26898 8752 26954
rect 8808 26898 8876 26954
rect 8932 26898 9000 26954
rect 9056 26898 9124 26954
rect 9180 26898 9248 26954
rect 9304 26898 9372 26954
rect 9428 26898 9496 26954
rect 9552 26898 9620 26954
rect 9676 26898 9744 26954
rect 9800 26898 9810 26954
rect 7874 26830 9810 26898
rect 7874 26774 7884 26830
rect 7940 26774 8008 26830
rect 8064 26774 8132 26830
rect 8188 26774 8256 26830
rect 8312 26774 8380 26830
rect 8436 26774 8504 26830
rect 8560 26774 8628 26830
rect 8684 26774 8752 26830
rect 8808 26774 8876 26830
rect 8932 26774 9000 26830
rect 9056 26774 9124 26830
rect 9180 26774 9248 26830
rect 9304 26774 9372 26830
rect 9428 26774 9496 26830
rect 9552 26774 9620 26830
rect 9676 26774 9744 26830
rect 9800 26774 9810 26830
rect 7874 26706 9810 26774
rect 7874 26650 7884 26706
rect 7940 26650 8008 26706
rect 8064 26650 8132 26706
rect 8188 26650 8256 26706
rect 8312 26650 8380 26706
rect 8436 26650 8504 26706
rect 8560 26650 8628 26706
rect 8684 26650 8752 26706
rect 8808 26650 8876 26706
rect 8932 26650 9000 26706
rect 9056 26650 9124 26706
rect 9180 26650 9248 26706
rect 9304 26650 9372 26706
rect 9428 26650 9496 26706
rect 9552 26650 9620 26706
rect 9676 26650 9744 26706
rect 9800 26650 9810 26706
rect 7874 26582 9810 26650
rect 7874 26526 7884 26582
rect 7940 26526 8008 26582
rect 8064 26526 8132 26582
rect 8188 26526 8256 26582
rect 8312 26526 8380 26582
rect 8436 26526 8504 26582
rect 8560 26526 8628 26582
rect 8684 26526 8752 26582
rect 8808 26526 8876 26582
rect 8932 26526 9000 26582
rect 9056 26526 9124 26582
rect 9180 26526 9248 26582
rect 9304 26526 9372 26582
rect 9428 26526 9496 26582
rect 9552 26526 9620 26582
rect 9676 26526 9744 26582
rect 9800 26526 9810 26582
rect 7874 26458 9810 26526
rect 7874 26402 7884 26458
rect 7940 26402 8008 26458
rect 8064 26402 8132 26458
rect 8188 26402 8256 26458
rect 8312 26402 8380 26458
rect 8436 26402 8504 26458
rect 8560 26402 8628 26458
rect 8684 26402 8752 26458
rect 8808 26402 8876 26458
rect 8932 26402 9000 26458
rect 9056 26402 9124 26458
rect 9180 26402 9248 26458
rect 9304 26402 9372 26458
rect 9428 26402 9496 26458
rect 9552 26402 9620 26458
rect 9676 26402 9744 26458
rect 9800 26402 9810 26458
rect 7874 26334 9810 26402
rect 7874 26278 7884 26334
rect 7940 26278 8008 26334
rect 8064 26278 8132 26334
rect 8188 26278 8256 26334
rect 8312 26278 8380 26334
rect 8436 26278 8504 26334
rect 8560 26278 8628 26334
rect 8684 26278 8752 26334
rect 8808 26278 8876 26334
rect 8932 26278 9000 26334
rect 9056 26278 9124 26334
rect 9180 26278 9248 26334
rect 9304 26278 9372 26334
rect 9428 26278 9496 26334
rect 9552 26278 9620 26334
rect 9676 26278 9744 26334
rect 9800 26278 9810 26334
rect 7874 26210 9810 26278
rect 7874 26154 7884 26210
rect 7940 26154 8008 26210
rect 8064 26154 8132 26210
rect 8188 26154 8256 26210
rect 8312 26154 8380 26210
rect 8436 26154 8504 26210
rect 8560 26154 8628 26210
rect 8684 26154 8752 26210
rect 8808 26154 8876 26210
rect 8932 26154 9000 26210
rect 9056 26154 9124 26210
rect 9180 26154 9248 26210
rect 9304 26154 9372 26210
rect 9428 26154 9496 26210
rect 9552 26154 9620 26210
rect 9676 26154 9744 26210
rect 9800 26154 9810 26210
rect 7874 26086 9810 26154
rect 7874 26030 7884 26086
rect 7940 26030 8008 26086
rect 8064 26030 8132 26086
rect 8188 26030 8256 26086
rect 8312 26030 8380 26086
rect 8436 26030 8504 26086
rect 8560 26030 8628 26086
rect 8684 26030 8752 26086
rect 8808 26030 8876 26086
rect 8932 26030 9000 26086
rect 9056 26030 9124 26086
rect 9180 26030 9248 26086
rect 9304 26030 9372 26086
rect 9428 26030 9496 26086
rect 9552 26030 9620 26086
rect 9676 26030 9744 26086
rect 9800 26030 9810 26086
rect 7874 25962 9810 26030
rect 7874 25906 7884 25962
rect 7940 25906 8008 25962
rect 8064 25906 8132 25962
rect 8188 25906 8256 25962
rect 8312 25906 8380 25962
rect 8436 25906 8504 25962
rect 8560 25906 8628 25962
rect 8684 25906 8752 25962
rect 8808 25906 8876 25962
rect 8932 25906 9000 25962
rect 9056 25906 9124 25962
rect 9180 25906 9248 25962
rect 9304 25906 9372 25962
rect 9428 25906 9496 25962
rect 9552 25906 9620 25962
rect 9676 25906 9744 25962
rect 9800 25906 9810 25962
rect 7874 25838 9810 25906
rect 7874 25782 7884 25838
rect 7940 25782 8008 25838
rect 8064 25782 8132 25838
rect 8188 25782 8256 25838
rect 8312 25782 8380 25838
rect 8436 25782 8504 25838
rect 8560 25782 8628 25838
rect 8684 25782 8752 25838
rect 8808 25782 8876 25838
rect 8932 25782 9000 25838
rect 9056 25782 9124 25838
rect 9180 25782 9248 25838
rect 9304 25782 9372 25838
rect 9428 25782 9496 25838
rect 9552 25782 9620 25838
rect 9676 25782 9744 25838
rect 9800 25782 9810 25838
rect 7874 25714 9810 25782
rect 7874 25658 7884 25714
rect 7940 25658 8008 25714
rect 8064 25658 8132 25714
rect 8188 25658 8256 25714
rect 8312 25658 8380 25714
rect 8436 25658 8504 25714
rect 8560 25658 8628 25714
rect 8684 25658 8752 25714
rect 8808 25658 8876 25714
rect 8932 25658 9000 25714
rect 9056 25658 9124 25714
rect 9180 25658 9248 25714
rect 9304 25658 9372 25714
rect 9428 25658 9496 25714
rect 9552 25658 9620 25714
rect 9676 25658 9744 25714
rect 9800 25658 9810 25714
rect 7874 25590 9810 25658
rect 7874 25534 7884 25590
rect 7940 25534 8008 25590
rect 8064 25534 8132 25590
rect 8188 25534 8256 25590
rect 8312 25534 8380 25590
rect 8436 25534 8504 25590
rect 8560 25534 8628 25590
rect 8684 25534 8752 25590
rect 8808 25534 8876 25590
rect 8932 25534 9000 25590
rect 9056 25534 9124 25590
rect 9180 25534 9248 25590
rect 9304 25534 9372 25590
rect 9428 25534 9496 25590
rect 9552 25534 9620 25590
rect 9676 25534 9744 25590
rect 9800 25534 9810 25590
rect 7874 25466 9810 25534
rect 7874 25410 7884 25466
rect 7940 25410 8008 25466
rect 8064 25410 8132 25466
rect 8188 25410 8256 25466
rect 8312 25410 8380 25466
rect 8436 25410 8504 25466
rect 8560 25410 8628 25466
rect 8684 25410 8752 25466
rect 8808 25410 8876 25466
rect 8932 25410 9000 25466
rect 9056 25410 9124 25466
rect 9180 25410 9248 25466
rect 9304 25410 9372 25466
rect 9428 25410 9496 25466
rect 9552 25410 9620 25466
rect 9676 25410 9744 25466
rect 9800 25410 9810 25466
rect 7874 25342 9810 25410
rect 7874 25286 7884 25342
rect 7940 25286 8008 25342
rect 8064 25286 8132 25342
rect 8188 25286 8256 25342
rect 8312 25286 8380 25342
rect 8436 25286 8504 25342
rect 8560 25286 8628 25342
rect 8684 25286 8752 25342
rect 8808 25286 8876 25342
rect 8932 25286 9000 25342
rect 9056 25286 9124 25342
rect 9180 25286 9248 25342
rect 9304 25286 9372 25342
rect 9428 25286 9496 25342
rect 9552 25286 9620 25342
rect 9676 25286 9744 25342
rect 9800 25286 9810 25342
rect 7874 25218 9810 25286
rect 7874 25162 7884 25218
rect 7940 25162 8008 25218
rect 8064 25162 8132 25218
rect 8188 25162 8256 25218
rect 8312 25162 8380 25218
rect 8436 25162 8504 25218
rect 8560 25162 8628 25218
rect 8684 25162 8752 25218
rect 8808 25162 8876 25218
rect 8932 25162 9000 25218
rect 9056 25162 9124 25218
rect 9180 25162 9248 25218
rect 9304 25162 9372 25218
rect 9428 25162 9496 25218
rect 9552 25162 9620 25218
rect 9676 25162 9744 25218
rect 9800 25162 9810 25218
rect 7874 25094 9810 25162
rect 7874 25038 7884 25094
rect 7940 25038 8008 25094
rect 8064 25038 8132 25094
rect 8188 25038 8256 25094
rect 8312 25038 8380 25094
rect 8436 25038 8504 25094
rect 8560 25038 8628 25094
rect 8684 25038 8752 25094
rect 8808 25038 8876 25094
rect 8932 25038 9000 25094
rect 9056 25038 9124 25094
rect 9180 25038 9248 25094
rect 9304 25038 9372 25094
rect 9428 25038 9496 25094
rect 9552 25038 9620 25094
rect 9676 25038 9744 25094
rect 9800 25038 9810 25094
rect 7874 24970 9810 25038
rect 7874 24914 7884 24970
rect 7940 24914 8008 24970
rect 8064 24914 8132 24970
rect 8188 24914 8256 24970
rect 8312 24914 8380 24970
rect 8436 24914 8504 24970
rect 8560 24914 8628 24970
rect 8684 24914 8752 24970
rect 8808 24914 8876 24970
rect 8932 24914 9000 24970
rect 9056 24914 9124 24970
rect 9180 24914 9248 24970
rect 9304 24914 9372 24970
rect 9428 24914 9496 24970
rect 9552 24914 9620 24970
rect 9676 24914 9744 24970
rect 9800 24914 9810 24970
rect 7874 24846 9810 24914
rect 7874 24790 7884 24846
rect 7940 24790 8008 24846
rect 8064 24790 8132 24846
rect 8188 24790 8256 24846
rect 8312 24790 8380 24846
rect 8436 24790 8504 24846
rect 8560 24790 8628 24846
rect 8684 24790 8752 24846
rect 8808 24790 8876 24846
rect 8932 24790 9000 24846
rect 9056 24790 9124 24846
rect 9180 24790 9248 24846
rect 9304 24790 9372 24846
rect 9428 24790 9496 24846
rect 9552 24790 9620 24846
rect 9676 24790 9744 24846
rect 9800 24790 9810 24846
rect 7874 24722 9810 24790
rect 7874 24666 7884 24722
rect 7940 24666 8008 24722
rect 8064 24666 8132 24722
rect 8188 24666 8256 24722
rect 8312 24666 8380 24722
rect 8436 24666 8504 24722
rect 8560 24666 8628 24722
rect 8684 24666 8752 24722
rect 8808 24666 8876 24722
rect 8932 24666 9000 24722
rect 9056 24666 9124 24722
rect 9180 24666 9248 24722
rect 9304 24666 9372 24722
rect 9428 24666 9496 24722
rect 9552 24666 9620 24722
rect 9676 24666 9744 24722
rect 9800 24666 9810 24722
rect 7874 24598 9810 24666
rect 7874 24542 7884 24598
rect 7940 24542 8008 24598
rect 8064 24542 8132 24598
rect 8188 24542 8256 24598
rect 8312 24542 8380 24598
rect 8436 24542 8504 24598
rect 8560 24542 8628 24598
rect 8684 24542 8752 24598
rect 8808 24542 8876 24598
rect 8932 24542 9000 24598
rect 9056 24542 9124 24598
rect 9180 24542 9248 24598
rect 9304 24542 9372 24598
rect 9428 24542 9496 24598
rect 9552 24542 9620 24598
rect 9676 24542 9744 24598
rect 9800 24542 9810 24598
rect 7874 24474 9810 24542
rect 7874 24418 7884 24474
rect 7940 24418 8008 24474
rect 8064 24418 8132 24474
rect 8188 24418 8256 24474
rect 8312 24418 8380 24474
rect 8436 24418 8504 24474
rect 8560 24418 8628 24474
rect 8684 24418 8752 24474
rect 8808 24418 8876 24474
rect 8932 24418 9000 24474
rect 9056 24418 9124 24474
rect 9180 24418 9248 24474
rect 9304 24418 9372 24474
rect 9428 24418 9496 24474
rect 9552 24418 9620 24474
rect 9676 24418 9744 24474
rect 9800 24418 9810 24474
rect 7874 24350 9810 24418
rect 7874 24294 7884 24350
rect 7940 24294 8008 24350
rect 8064 24294 8132 24350
rect 8188 24294 8256 24350
rect 8312 24294 8380 24350
rect 8436 24294 8504 24350
rect 8560 24294 8628 24350
rect 8684 24294 8752 24350
rect 8808 24294 8876 24350
rect 8932 24294 9000 24350
rect 9056 24294 9124 24350
rect 9180 24294 9248 24350
rect 9304 24294 9372 24350
rect 9428 24294 9496 24350
rect 9552 24294 9620 24350
rect 9676 24294 9744 24350
rect 9800 24294 9810 24350
rect 7874 24226 9810 24294
rect 7874 24170 7884 24226
rect 7940 24170 8008 24226
rect 8064 24170 8132 24226
rect 8188 24170 8256 24226
rect 8312 24170 8380 24226
rect 8436 24170 8504 24226
rect 8560 24170 8628 24226
rect 8684 24170 8752 24226
rect 8808 24170 8876 24226
rect 8932 24170 9000 24226
rect 9056 24170 9124 24226
rect 9180 24170 9248 24226
rect 9304 24170 9372 24226
rect 9428 24170 9496 24226
rect 9552 24170 9620 24226
rect 9676 24170 9744 24226
rect 9800 24170 9810 24226
rect 7874 24102 9810 24170
rect 7874 24046 7884 24102
rect 7940 24046 8008 24102
rect 8064 24046 8132 24102
rect 8188 24046 8256 24102
rect 8312 24046 8380 24102
rect 8436 24046 8504 24102
rect 8560 24046 8628 24102
rect 8684 24046 8752 24102
rect 8808 24046 8876 24102
rect 8932 24046 9000 24102
rect 9056 24046 9124 24102
rect 9180 24046 9248 24102
rect 9304 24046 9372 24102
rect 9428 24046 9496 24102
rect 9552 24046 9620 24102
rect 9676 24046 9744 24102
rect 9800 24046 9810 24102
rect 7874 24036 9810 24046
rect 10244 26954 12180 26964
rect 10244 26898 10254 26954
rect 10310 26898 10378 26954
rect 10434 26898 10502 26954
rect 10558 26898 10626 26954
rect 10682 26898 10750 26954
rect 10806 26898 10874 26954
rect 10930 26898 10998 26954
rect 11054 26898 11122 26954
rect 11178 26898 11246 26954
rect 11302 26898 11370 26954
rect 11426 26898 11494 26954
rect 11550 26898 11618 26954
rect 11674 26898 11742 26954
rect 11798 26898 11866 26954
rect 11922 26898 11990 26954
rect 12046 26898 12114 26954
rect 12170 26898 12180 26954
rect 10244 26830 12180 26898
rect 10244 26774 10254 26830
rect 10310 26774 10378 26830
rect 10434 26774 10502 26830
rect 10558 26774 10626 26830
rect 10682 26774 10750 26830
rect 10806 26774 10874 26830
rect 10930 26774 10998 26830
rect 11054 26774 11122 26830
rect 11178 26774 11246 26830
rect 11302 26774 11370 26830
rect 11426 26774 11494 26830
rect 11550 26774 11618 26830
rect 11674 26774 11742 26830
rect 11798 26774 11866 26830
rect 11922 26774 11990 26830
rect 12046 26774 12114 26830
rect 12170 26774 12180 26830
rect 10244 26706 12180 26774
rect 10244 26650 10254 26706
rect 10310 26650 10378 26706
rect 10434 26650 10502 26706
rect 10558 26650 10626 26706
rect 10682 26650 10750 26706
rect 10806 26650 10874 26706
rect 10930 26650 10998 26706
rect 11054 26650 11122 26706
rect 11178 26650 11246 26706
rect 11302 26650 11370 26706
rect 11426 26650 11494 26706
rect 11550 26650 11618 26706
rect 11674 26650 11742 26706
rect 11798 26650 11866 26706
rect 11922 26650 11990 26706
rect 12046 26650 12114 26706
rect 12170 26650 12180 26706
rect 10244 26582 12180 26650
rect 10244 26526 10254 26582
rect 10310 26526 10378 26582
rect 10434 26526 10502 26582
rect 10558 26526 10626 26582
rect 10682 26526 10750 26582
rect 10806 26526 10874 26582
rect 10930 26526 10998 26582
rect 11054 26526 11122 26582
rect 11178 26526 11246 26582
rect 11302 26526 11370 26582
rect 11426 26526 11494 26582
rect 11550 26526 11618 26582
rect 11674 26526 11742 26582
rect 11798 26526 11866 26582
rect 11922 26526 11990 26582
rect 12046 26526 12114 26582
rect 12170 26526 12180 26582
rect 10244 26458 12180 26526
rect 10244 26402 10254 26458
rect 10310 26402 10378 26458
rect 10434 26402 10502 26458
rect 10558 26402 10626 26458
rect 10682 26402 10750 26458
rect 10806 26402 10874 26458
rect 10930 26402 10998 26458
rect 11054 26402 11122 26458
rect 11178 26402 11246 26458
rect 11302 26402 11370 26458
rect 11426 26402 11494 26458
rect 11550 26402 11618 26458
rect 11674 26402 11742 26458
rect 11798 26402 11866 26458
rect 11922 26402 11990 26458
rect 12046 26402 12114 26458
rect 12170 26402 12180 26458
rect 10244 26334 12180 26402
rect 10244 26278 10254 26334
rect 10310 26278 10378 26334
rect 10434 26278 10502 26334
rect 10558 26278 10626 26334
rect 10682 26278 10750 26334
rect 10806 26278 10874 26334
rect 10930 26278 10998 26334
rect 11054 26278 11122 26334
rect 11178 26278 11246 26334
rect 11302 26278 11370 26334
rect 11426 26278 11494 26334
rect 11550 26278 11618 26334
rect 11674 26278 11742 26334
rect 11798 26278 11866 26334
rect 11922 26278 11990 26334
rect 12046 26278 12114 26334
rect 12170 26278 12180 26334
rect 10244 26210 12180 26278
rect 10244 26154 10254 26210
rect 10310 26154 10378 26210
rect 10434 26154 10502 26210
rect 10558 26154 10626 26210
rect 10682 26154 10750 26210
rect 10806 26154 10874 26210
rect 10930 26154 10998 26210
rect 11054 26154 11122 26210
rect 11178 26154 11246 26210
rect 11302 26154 11370 26210
rect 11426 26154 11494 26210
rect 11550 26154 11618 26210
rect 11674 26154 11742 26210
rect 11798 26154 11866 26210
rect 11922 26154 11990 26210
rect 12046 26154 12114 26210
rect 12170 26154 12180 26210
rect 10244 26086 12180 26154
rect 10244 26030 10254 26086
rect 10310 26030 10378 26086
rect 10434 26030 10502 26086
rect 10558 26030 10626 26086
rect 10682 26030 10750 26086
rect 10806 26030 10874 26086
rect 10930 26030 10998 26086
rect 11054 26030 11122 26086
rect 11178 26030 11246 26086
rect 11302 26030 11370 26086
rect 11426 26030 11494 26086
rect 11550 26030 11618 26086
rect 11674 26030 11742 26086
rect 11798 26030 11866 26086
rect 11922 26030 11990 26086
rect 12046 26030 12114 26086
rect 12170 26030 12180 26086
rect 10244 25962 12180 26030
rect 10244 25906 10254 25962
rect 10310 25906 10378 25962
rect 10434 25906 10502 25962
rect 10558 25906 10626 25962
rect 10682 25906 10750 25962
rect 10806 25906 10874 25962
rect 10930 25906 10998 25962
rect 11054 25906 11122 25962
rect 11178 25906 11246 25962
rect 11302 25906 11370 25962
rect 11426 25906 11494 25962
rect 11550 25906 11618 25962
rect 11674 25906 11742 25962
rect 11798 25906 11866 25962
rect 11922 25906 11990 25962
rect 12046 25906 12114 25962
rect 12170 25906 12180 25962
rect 10244 25838 12180 25906
rect 10244 25782 10254 25838
rect 10310 25782 10378 25838
rect 10434 25782 10502 25838
rect 10558 25782 10626 25838
rect 10682 25782 10750 25838
rect 10806 25782 10874 25838
rect 10930 25782 10998 25838
rect 11054 25782 11122 25838
rect 11178 25782 11246 25838
rect 11302 25782 11370 25838
rect 11426 25782 11494 25838
rect 11550 25782 11618 25838
rect 11674 25782 11742 25838
rect 11798 25782 11866 25838
rect 11922 25782 11990 25838
rect 12046 25782 12114 25838
rect 12170 25782 12180 25838
rect 10244 25714 12180 25782
rect 10244 25658 10254 25714
rect 10310 25658 10378 25714
rect 10434 25658 10502 25714
rect 10558 25658 10626 25714
rect 10682 25658 10750 25714
rect 10806 25658 10874 25714
rect 10930 25658 10998 25714
rect 11054 25658 11122 25714
rect 11178 25658 11246 25714
rect 11302 25658 11370 25714
rect 11426 25658 11494 25714
rect 11550 25658 11618 25714
rect 11674 25658 11742 25714
rect 11798 25658 11866 25714
rect 11922 25658 11990 25714
rect 12046 25658 12114 25714
rect 12170 25658 12180 25714
rect 10244 25590 12180 25658
rect 10244 25534 10254 25590
rect 10310 25534 10378 25590
rect 10434 25534 10502 25590
rect 10558 25534 10626 25590
rect 10682 25534 10750 25590
rect 10806 25534 10874 25590
rect 10930 25534 10998 25590
rect 11054 25534 11122 25590
rect 11178 25534 11246 25590
rect 11302 25534 11370 25590
rect 11426 25534 11494 25590
rect 11550 25534 11618 25590
rect 11674 25534 11742 25590
rect 11798 25534 11866 25590
rect 11922 25534 11990 25590
rect 12046 25534 12114 25590
rect 12170 25534 12180 25590
rect 10244 25466 12180 25534
rect 10244 25410 10254 25466
rect 10310 25410 10378 25466
rect 10434 25410 10502 25466
rect 10558 25410 10626 25466
rect 10682 25410 10750 25466
rect 10806 25410 10874 25466
rect 10930 25410 10998 25466
rect 11054 25410 11122 25466
rect 11178 25410 11246 25466
rect 11302 25410 11370 25466
rect 11426 25410 11494 25466
rect 11550 25410 11618 25466
rect 11674 25410 11742 25466
rect 11798 25410 11866 25466
rect 11922 25410 11990 25466
rect 12046 25410 12114 25466
rect 12170 25410 12180 25466
rect 10244 25342 12180 25410
rect 10244 25286 10254 25342
rect 10310 25286 10378 25342
rect 10434 25286 10502 25342
rect 10558 25286 10626 25342
rect 10682 25286 10750 25342
rect 10806 25286 10874 25342
rect 10930 25286 10998 25342
rect 11054 25286 11122 25342
rect 11178 25286 11246 25342
rect 11302 25286 11370 25342
rect 11426 25286 11494 25342
rect 11550 25286 11618 25342
rect 11674 25286 11742 25342
rect 11798 25286 11866 25342
rect 11922 25286 11990 25342
rect 12046 25286 12114 25342
rect 12170 25286 12180 25342
rect 10244 25218 12180 25286
rect 10244 25162 10254 25218
rect 10310 25162 10378 25218
rect 10434 25162 10502 25218
rect 10558 25162 10626 25218
rect 10682 25162 10750 25218
rect 10806 25162 10874 25218
rect 10930 25162 10998 25218
rect 11054 25162 11122 25218
rect 11178 25162 11246 25218
rect 11302 25162 11370 25218
rect 11426 25162 11494 25218
rect 11550 25162 11618 25218
rect 11674 25162 11742 25218
rect 11798 25162 11866 25218
rect 11922 25162 11990 25218
rect 12046 25162 12114 25218
rect 12170 25162 12180 25218
rect 10244 25094 12180 25162
rect 10244 25038 10254 25094
rect 10310 25038 10378 25094
rect 10434 25038 10502 25094
rect 10558 25038 10626 25094
rect 10682 25038 10750 25094
rect 10806 25038 10874 25094
rect 10930 25038 10998 25094
rect 11054 25038 11122 25094
rect 11178 25038 11246 25094
rect 11302 25038 11370 25094
rect 11426 25038 11494 25094
rect 11550 25038 11618 25094
rect 11674 25038 11742 25094
rect 11798 25038 11866 25094
rect 11922 25038 11990 25094
rect 12046 25038 12114 25094
rect 12170 25038 12180 25094
rect 10244 24970 12180 25038
rect 10244 24914 10254 24970
rect 10310 24914 10378 24970
rect 10434 24914 10502 24970
rect 10558 24914 10626 24970
rect 10682 24914 10750 24970
rect 10806 24914 10874 24970
rect 10930 24914 10998 24970
rect 11054 24914 11122 24970
rect 11178 24914 11246 24970
rect 11302 24914 11370 24970
rect 11426 24914 11494 24970
rect 11550 24914 11618 24970
rect 11674 24914 11742 24970
rect 11798 24914 11866 24970
rect 11922 24914 11990 24970
rect 12046 24914 12114 24970
rect 12170 24914 12180 24970
rect 10244 24846 12180 24914
rect 10244 24790 10254 24846
rect 10310 24790 10378 24846
rect 10434 24790 10502 24846
rect 10558 24790 10626 24846
rect 10682 24790 10750 24846
rect 10806 24790 10874 24846
rect 10930 24790 10998 24846
rect 11054 24790 11122 24846
rect 11178 24790 11246 24846
rect 11302 24790 11370 24846
rect 11426 24790 11494 24846
rect 11550 24790 11618 24846
rect 11674 24790 11742 24846
rect 11798 24790 11866 24846
rect 11922 24790 11990 24846
rect 12046 24790 12114 24846
rect 12170 24790 12180 24846
rect 10244 24722 12180 24790
rect 10244 24666 10254 24722
rect 10310 24666 10378 24722
rect 10434 24666 10502 24722
rect 10558 24666 10626 24722
rect 10682 24666 10750 24722
rect 10806 24666 10874 24722
rect 10930 24666 10998 24722
rect 11054 24666 11122 24722
rect 11178 24666 11246 24722
rect 11302 24666 11370 24722
rect 11426 24666 11494 24722
rect 11550 24666 11618 24722
rect 11674 24666 11742 24722
rect 11798 24666 11866 24722
rect 11922 24666 11990 24722
rect 12046 24666 12114 24722
rect 12170 24666 12180 24722
rect 10244 24598 12180 24666
rect 10244 24542 10254 24598
rect 10310 24542 10378 24598
rect 10434 24542 10502 24598
rect 10558 24542 10626 24598
rect 10682 24542 10750 24598
rect 10806 24542 10874 24598
rect 10930 24542 10998 24598
rect 11054 24542 11122 24598
rect 11178 24542 11246 24598
rect 11302 24542 11370 24598
rect 11426 24542 11494 24598
rect 11550 24542 11618 24598
rect 11674 24542 11742 24598
rect 11798 24542 11866 24598
rect 11922 24542 11990 24598
rect 12046 24542 12114 24598
rect 12170 24542 12180 24598
rect 10244 24474 12180 24542
rect 10244 24418 10254 24474
rect 10310 24418 10378 24474
rect 10434 24418 10502 24474
rect 10558 24418 10626 24474
rect 10682 24418 10750 24474
rect 10806 24418 10874 24474
rect 10930 24418 10998 24474
rect 11054 24418 11122 24474
rect 11178 24418 11246 24474
rect 11302 24418 11370 24474
rect 11426 24418 11494 24474
rect 11550 24418 11618 24474
rect 11674 24418 11742 24474
rect 11798 24418 11866 24474
rect 11922 24418 11990 24474
rect 12046 24418 12114 24474
rect 12170 24418 12180 24474
rect 10244 24350 12180 24418
rect 10244 24294 10254 24350
rect 10310 24294 10378 24350
rect 10434 24294 10502 24350
rect 10558 24294 10626 24350
rect 10682 24294 10750 24350
rect 10806 24294 10874 24350
rect 10930 24294 10998 24350
rect 11054 24294 11122 24350
rect 11178 24294 11246 24350
rect 11302 24294 11370 24350
rect 11426 24294 11494 24350
rect 11550 24294 11618 24350
rect 11674 24294 11742 24350
rect 11798 24294 11866 24350
rect 11922 24294 11990 24350
rect 12046 24294 12114 24350
rect 12170 24294 12180 24350
rect 10244 24226 12180 24294
rect 10244 24170 10254 24226
rect 10310 24170 10378 24226
rect 10434 24170 10502 24226
rect 10558 24170 10626 24226
rect 10682 24170 10750 24226
rect 10806 24170 10874 24226
rect 10930 24170 10998 24226
rect 11054 24170 11122 24226
rect 11178 24170 11246 24226
rect 11302 24170 11370 24226
rect 11426 24170 11494 24226
rect 11550 24170 11618 24226
rect 11674 24170 11742 24226
rect 11798 24170 11866 24226
rect 11922 24170 11990 24226
rect 12046 24170 12114 24226
rect 12170 24170 12180 24226
rect 10244 24102 12180 24170
rect 10244 24046 10254 24102
rect 10310 24046 10378 24102
rect 10434 24046 10502 24102
rect 10558 24046 10626 24102
rect 10682 24046 10750 24102
rect 10806 24046 10874 24102
rect 10930 24046 10998 24102
rect 11054 24046 11122 24102
rect 11178 24046 11246 24102
rect 11302 24046 11370 24102
rect 11426 24046 11494 24102
rect 11550 24046 11618 24102
rect 11674 24046 11742 24102
rect 11798 24046 11866 24102
rect 11922 24046 11990 24102
rect 12046 24046 12114 24102
rect 12170 24046 12180 24102
rect 10244 24036 12180 24046
rect 12861 26954 14673 26964
rect 12861 26898 12871 26954
rect 12927 26898 12995 26954
rect 13051 26898 13119 26954
rect 13175 26898 13243 26954
rect 13299 26898 13367 26954
rect 13423 26898 13491 26954
rect 13547 26898 13615 26954
rect 13671 26898 13739 26954
rect 13795 26898 13863 26954
rect 13919 26898 13987 26954
rect 14043 26898 14111 26954
rect 14167 26898 14235 26954
rect 14291 26898 14359 26954
rect 14415 26898 14483 26954
rect 14539 26898 14607 26954
rect 14663 26898 14673 26954
rect 12861 26830 14673 26898
rect 12861 26774 12871 26830
rect 12927 26774 12995 26830
rect 13051 26774 13119 26830
rect 13175 26774 13243 26830
rect 13299 26774 13367 26830
rect 13423 26774 13491 26830
rect 13547 26774 13615 26830
rect 13671 26774 13739 26830
rect 13795 26774 13863 26830
rect 13919 26774 13987 26830
rect 14043 26774 14111 26830
rect 14167 26774 14235 26830
rect 14291 26774 14359 26830
rect 14415 26774 14483 26830
rect 14539 26774 14607 26830
rect 14663 26774 14673 26830
rect 12861 26706 14673 26774
rect 12861 26650 12871 26706
rect 12927 26650 12995 26706
rect 13051 26650 13119 26706
rect 13175 26650 13243 26706
rect 13299 26650 13367 26706
rect 13423 26650 13491 26706
rect 13547 26650 13615 26706
rect 13671 26650 13739 26706
rect 13795 26650 13863 26706
rect 13919 26650 13987 26706
rect 14043 26650 14111 26706
rect 14167 26650 14235 26706
rect 14291 26650 14359 26706
rect 14415 26650 14483 26706
rect 14539 26650 14607 26706
rect 14663 26650 14673 26706
rect 12861 26582 14673 26650
rect 12861 26526 12871 26582
rect 12927 26526 12995 26582
rect 13051 26526 13119 26582
rect 13175 26526 13243 26582
rect 13299 26526 13367 26582
rect 13423 26526 13491 26582
rect 13547 26526 13615 26582
rect 13671 26526 13739 26582
rect 13795 26526 13863 26582
rect 13919 26526 13987 26582
rect 14043 26526 14111 26582
rect 14167 26526 14235 26582
rect 14291 26526 14359 26582
rect 14415 26526 14483 26582
rect 14539 26526 14607 26582
rect 14663 26526 14673 26582
rect 12861 26458 14673 26526
rect 12861 26402 12871 26458
rect 12927 26402 12995 26458
rect 13051 26402 13119 26458
rect 13175 26402 13243 26458
rect 13299 26402 13367 26458
rect 13423 26402 13491 26458
rect 13547 26402 13615 26458
rect 13671 26402 13739 26458
rect 13795 26402 13863 26458
rect 13919 26402 13987 26458
rect 14043 26402 14111 26458
rect 14167 26402 14235 26458
rect 14291 26402 14359 26458
rect 14415 26402 14483 26458
rect 14539 26402 14607 26458
rect 14663 26402 14673 26458
rect 12861 26334 14673 26402
rect 12861 26278 12871 26334
rect 12927 26278 12995 26334
rect 13051 26278 13119 26334
rect 13175 26278 13243 26334
rect 13299 26278 13367 26334
rect 13423 26278 13491 26334
rect 13547 26278 13615 26334
rect 13671 26278 13739 26334
rect 13795 26278 13863 26334
rect 13919 26278 13987 26334
rect 14043 26278 14111 26334
rect 14167 26278 14235 26334
rect 14291 26278 14359 26334
rect 14415 26278 14483 26334
rect 14539 26278 14607 26334
rect 14663 26278 14673 26334
rect 12861 26210 14673 26278
rect 12861 26154 12871 26210
rect 12927 26154 12995 26210
rect 13051 26154 13119 26210
rect 13175 26154 13243 26210
rect 13299 26154 13367 26210
rect 13423 26154 13491 26210
rect 13547 26154 13615 26210
rect 13671 26154 13739 26210
rect 13795 26154 13863 26210
rect 13919 26154 13987 26210
rect 14043 26154 14111 26210
rect 14167 26154 14235 26210
rect 14291 26154 14359 26210
rect 14415 26154 14483 26210
rect 14539 26154 14607 26210
rect 14663 26154 14673 26210
rect 12861 26086 14673 26154
rect 12861 26030 12871 26086
rect 12927 26030 12995 26086
rect 13051 26030 13119 26086
rect 13175 26030 13243 26086
rect 13299 26030 13367 26086
rect 13423 26030 13491 26086
rect 13547 26030 13615 26086
rect 13671 26030 13739 26086
rect 13795 26030 13863 26086
rect 13919 26030 13987 26086
rect 14043 26030 14111 26086
rect 14167 26030 14235 26086
rect 14291 26030 14359 26086
rect 14415 26030 14483 26086
rect 14539 26030 14607 26086
rect 14663 26030 14673 26086
rect 12861 25962 14673 26030
rect 12861 25906 12871 25962
rect 12927 25906 12995 25962
rect 13051 25906 13119 25962
rect 13175 25906 13243 25962
rect 13299 25906 13367 25962
rect 13423 25906 13491 25962
rect 13547 25906 13615 25962
rect 13671 25906 13739 25962
rect 13795 25906 13863 25962
rect 13919 25906 13987 25962
rect 14043 25906 14111 25962
rect 14167 25906 14235 25962
rect 14291 25906 14359 25962
rect 14415 25906 14483 25962
rect 14539 25906 14607 25962
rect 14663 25906 14673 25962
rect 12861 25838 14673 25906
rect 12861 25782 12871 25838
rect 12927 25782 12995 25838
rect 13051 25782 13119 25838
rect 13175 25782 13243 25838
rect 13299 25782 13367 25838
rect 13423 25782 13491 25838
rect 13547 25782 13615 25838
rect 13671 25782 13739 25838
rect 13795 25782 13863 25838
rect 13919 25782 13987 25838
rect 14043 25782 14111 25838
rect 14167 25782 14235 25838
rect 14291 25782 14359 25838
rect 14415 25782 14483 25838
rect 14539 25782 14607 25838
rect 14663 25782 14673 25838
rect 12861 25714 14673 25782
rect 12861 25658 12871 25714
rect 12927 25658 12995 25714
rect 13051 25658 13119 25714
rect 13175 25658 13243 25714
rect 13299 25658 13367 25714
rect 13423 25658 13491 25714
rect 13547 25658 13615 25714
rect 13671 25658 13739 25714
rect 13795 25658 13863 25714
rect 13919 25658 13987 25714
rect 14043 25658 14111 25714
rect 14167 25658 14235 25714
rect 14291 25658 14359 25714
rect 14415 25658 14483 25714
rect 14539 25658 14607 25714
rect 14663 25658 14673 25714
rect 12861 25590 14673 25658
rect 12861 25534 12871 25590
rect 12927 25534 12995 25590
rect 13051 25534 13119 25590
rect 13175 25534 13243 25590
rect 13299 25534 13367 25590
rect 13423 25534 13491 25590
rect 13547 25534 13615 25590
rect 13671 25534 13739 25590
rect 13795 25534 13863 25590
rect 13919 25534 13987 25590
rect 14043 25534 14111 25590
rect 14167 25534 14235 25590
rect 14291 25534 14359 25590
rect 14415 25534 14483 25590
rect 14539 25534 14607 25590
rect 14663 25534 14673 25590
rect 12861 25466 14673 25534
rect 12861 25410 12871 25466
rect 12927 25410 12995 25466
rect 13051 25410 13119 25466
rect 13175 25410 13243 25466
rect 13299 25410 13367 25466
rect 13423 25410 13491 25466
rect 13547 25410 13615 25466
rect 13671 25410 13739 25466
rect 13795 25410 13863 25466
rect 13919 25410 13987 25466
rect 14043 25410 14111 25466
rect 14167 25410 14235 25466
rect 14291 25410 14359 25466
rect 14415 25410 14483 25466
rect 14539 25410 14607 25466
rect 14663 25410 14673 25466
rect 12861 25342 14673 25410
rect 12861 25286 12871 25342
rect 12927 25286 12995 25342
rect 13051 25286 13119 25342
rect 13175 25286 13243 25342
rect 13299 25286 13367 25342
rect 13423 25286 13491 25342
rect 13547 25286 13615 25342
rect 13671 25286 13739 25342
rect 13795 25286 13863 25342
rect 13919 25286 13987 25342
rect 14043 25286 14111 25342
rect 14167 25286 14235 25342
rect 14291 25286 14359 25342
rect 14415 25286 14483 25342
rect 14539 25286 14607 25342
rect 14663 25286 14673 25342
rect 12861 25218 14673 25286
rect 12861 25162 12871 25218
rect 12927 25162 12995 25218
rect 13051 25162 13119 25218
rect 13175 25162 13243 25218
rect 13299 25162 13367 25218
rect 13423 25162 13491 25218
rect 13547 25162 13615 25218
rect 13671 25162 13739 25218
rect 13795 25162 13863 25218
rect 13919 25162 13987 25218
rect 14043 25162 14111 25218
rect 14167 25162 14235 25218
rect 14291 25162 14359 25218
rect 14415 25162 14483 25218
rect 14539 25162 14607 25218
rect 14663 25162 14673 25218
rect 12861 25094 14673 25162
rect 12861 25038 12871 25094
rect 12927 25038 12995 25094
rect 13051 25038 13119 25094
rect 13175 25038 13243 25094
rect 13299 25038 13367 25094
rect 13423 25038 13491 25094
rect 13547 25038 13615 25094
rect 13671 25038 13739 25094
rect 13795 25038 13863 25094
rect 13919 25038 13987 25094
rect 14043 25038 14111 25094
rect 14167 25038 14235 25094
rect 14291 25038 14359 25094
rect 14415 25038 14483 25094
rect 14539 25038 14607 25094
rect 14663 25038 14673 25094
rect 12861 24970 14673 25038
rect 12861 24914 12871 24970
rect 12927 24914 12995 24970
rect 13051 24914 13119 24970
rect 13175 24914 13243 24970
rect 13299 24914 13367 24970
rect 13423 24914 13491 24970
rect 13547 24914 13615 24970
rect 13671 24914 13739 24970
rect 13795 24914 13863 24970
rect 13919 24914 13987 24970
rect 14043 24914 14111 24970
rect 14167 24914 14235 24970
rect 14291 24914 14359 24970
rect 14415 24914 14483 24970
rect 14539 24914 14607 24970
rect 14663 24914 14673 24970
rect 12861 24846 14673 24914
rect 12861 24790 12871 24846
rect 12927 24790 12995 24846
rect 13051 24790 13119 24846
rect 13175 24790 13243 24846
rect 13299 24790 13367 24846
rect 13423 24790 13491 24846
rect 13547 24790 13615 24846
rect 13671 24790 13739 24846
rect 13795 24790 13863 24846
rect 13919 24790 13987 24846
rect 14043 24790 14111 24846
rect 14167 24790 14235 24846
rect 14291 24790 14359 24846
rect 14415 24790 14483 24846
rect 14539 24790 14607 24846
rect 14663 24790 14673 24846
rect 12861 24722 14673 24790
rect 12861 24666 12871 24722
rect 12927 24666 12995 24722
rect 13051 24666 13119 24722
rect 13175 24666 13243 24722
rect 13299 24666 13367 24722
rect 13423 24666 13491 24722
rect 13547 24666 13615 24722
rect 13671 24666 13739 24722
rect 13795 24666 13863 24722
rect 13919 24666 13987 24722
rect 14043 24666 14111 24722
rect 14167 24666 14235 24722
rect 14291 24666 14359 24722
rect 14415 24666 14483 24722
rect 14539 24666 14607 24722
rect 14663 24666 14673 24722
rect 12861 24598 14673 24666
rect 12861 24542 12871 24598
rect 12927 24542 12995 24598
rect 13051 24542 13119 24598
rect 13175 24542 13243 24598
rect 13299 24542 13367 24598
rect 13423 24542 13491 24598
rect 13547 24542 13615 24598
rect 13671 24542 13739 24598
rect 13795 24542 13863 24598
rect 13919 24542 13987 24598
rect 14043 24542 14111 24598
rect 14167 24542 14235 24598
rect 14291 24542 14359 24598
rect 14415 24542 14483 24598
rect 14539 24542 14607 24598
rect 14663 24542 14673 24598
rect 12861 24474 14673 24542
rect 12861 24418 12871 24474
rect 12927 24418 12995 24474
rect 13051 24418 13119 24474
rect 13175 24418 13243 24474
rect 13299 24418 13367 24474
rect 13423 24418 13491 24474
rect 13547 24418 13615 24474
rect 13671 24418 13739 24474
rect 13795 24418 13863 24474
rect 13919 24418 13987 24474
rect 14043 24418 14111 24474
rect 14167 24418 14235 24474
rect 14291 24418 14359 24474
rect 14415 24418 14483 24474
rect 14539 24418 14607 24474
rect 14663 24418 14673 24474
rect 12861 24350 14673 24418
rect 12861 24294 12871 24350
rect 12927 24294 12995 24350
rect 13051 24294 13119 24350
rect 13175 24294 13243 24350
rect 13299 24294 13367 24350
rect 13423 24294 13491 24350
rect 13547 24294 13615 24350
rect 13671 24294 13739 24350
rect 13795 24294 13863 24350
rect 13919 24294 13987 24350
rect 14043 24294 14111 24350
rect 14167 24294 14235 24350
rect 14291 24294 14359 24350
rect 14415 24294 14483 24350
rect 14539 24294 14607 24350
rect 14663 24294 14673 24350
rect 12861 24226 14673 24294
rect 12861 24170 12871 24226
rect 12927 24170 12995 24226
rect 13051 24170 13119 24226
rect 13175 24170 13243 24226
rect 13299 24170 13367 24226
rect 13423 24170 13491 24226
rect 13547 24170 13615 24226
rect 13671 24170 13739 24226
rect 13795 24170 13863 24226
rect 13919 24170 13987 24226
rect 14043 24170 14111 24226
rect 14167 24170 14235 24226
rect 14291 24170 14359 24226
rect 14415 24170 14483 24226
rect 14539 24170 14607 24226
rect 14663 24170 14673 24226
rect 12861 24102 14673 24170
rect 12861 24046 12871 24102
rect 12927 24046 12995 24102
rect 13051 24046 13119 24102
rect 13175 24046 13243 24102
rect 13299 24046 13367 24102
rect 13423 24046 13491 24102
rect 13547 24046 13615 24102
rect 13671 24046 13739 24102
rect 13795 24046 13863 24102
rect 13919 24046 13987 24102
rect 14043 24046 14111 24102
rect 14167 24046 14235 24102
rect 14291 24046 14359 24102
rect 14415 24046 14483 24102
rect 14539 24046 14607 24102
rect 14663 24046 14673 24102
rect 12861 24036 14673 24046
rect 305 23754 2117 23764
rect 305 23698 315 23754
rect 371 23698 439 23754
rect 495 23698 563 23754
rect 619 23698 687 23754
rect 743 23698 811 23754
rect 867 23698 935 23754
rect 991 23698 1059 23754
rect 1115 23698 1183 23754
rect 1239 23698 1307 23754
rect 1363 23698 1431 23754
rect 1487 23698 1555 23754
rect 1611 23698 1679 23754
rect 1735 23698 1803 23754
rect 1859 23698 1927 23754
rect 1983 23698 2051 23754
rect 2107 23698 2117 23754
rect 305 23630 2117 23698
rect 305 23574 315 23630
rect 371 23574 439 23630
rect 495 23574 563 23630
rect 619 23574 687 23630
rect 743 23574 811 23630
rect 867 23574 935 23630
rect 991 23574 1059 23630
rect 1115 23574 1183 23630
rect 1239 23574 1307 23630
rect 1363 23574 1431 23630
rect 1487 23574 1555 23630
rect 1611 23574 1679 23630
rect 1735 23574 1803 23630
rect 1859 23574 1927 23630
rect 1983 23574 2051 23630
rect 2107 23574 2117 23630
rect 305 23506 2117 23574
rect 305 23450 315 23506
rect 371 23450 439 23506
rect 495 23450 563 23506
rect 619 23450 687 23506
rect 743 23450 811 23506
rect 867 23450 935 23506
rect 991 23450 1059 23506
rect 1115 23450 1183 23506
rect 1239 23450 1307 23506
rect 1363 23450 1431 23506
rect 1487 23450 1555 23506
rect 1611 23450 1679 23506
rect 1735 23450 1803 23506
rect 1859 23450 1927 23506
rect 1983 23450 2051 23506
rect 2107 23450 2117 23506
rect 305 23382 2117 23450
rect 305 23326 315 23382
rect 371 23326 439 23382
rect 495 23326 563 23382
rect 619 23326 687 23382
rect 743 23326 811 23382
rect 867 23326 935 23382
rect 991 23326 1059 23382
rect 1115 23326 1183 23382
rect 1239 23326 1307 23382
rect 1363 23326 1431 23382
rect 1487 23326 1555 23382
rect 1611 23326 1679 23382
rect 1735 23326 1803 23382
rect 1859 23326 1927 23382
rect 1983 23326 2051 23382
rect 2107 23326 2117 23382
rect 305 23258 2117 23326
rect 305 23202 315 23258
rect 371 23202 439 23258
rect 495 23202 563 23258
rect 619 23202 687 23258
rect 743 23202 811 23258
rect 867 23202 935 23258
rect 991 23202 1059 23258
rect 1115 23202 1183 23258
rect 1239 23202 1307 23258
rect 1363 23202 1431 23258
rect 1487 23202 1555 23258
rect 1611 23202 1679 23258
rect 1735 23202 1803 23258
rect 1859 23202 1927 23258
rect 1983 23202 2051 23258
rect 2107 23202 2117 23258
rect 305 23134 2117 23202
rect 305 23078 315 23134
rect 371 23078 439 23134
rect 495 23078 563 23134
rect 619 23078 687 23134
rect 743 23078 811 23134
rect 867 23078 935 23134
rect 991 23078 1059 23134
rect 1115 23078 1183 23134
rect 1239 23078 1307 23134
rect 1363 23078 1431 23134
rect 1487 23078 1555 23134
rect 1611 23078 1679 23134
rect 1735 23078 1803 23134
rect 1859 23078 1927 23134
rect 1983 23078 2051 23134
rect 2107 23078 2117 23134
rect 305 23010 2117 23078
rect 305 22954 315 23010
rect 371 22954 439 23010
rect 495 22954 563 23010
rect 619 22954 687 23010
rect 743 22954 811 23010
rect 867 22954 935 23010
rect 991 22954 1059 23010
rect 1115 22954 1183 23010
rect 1239 22954 1307 23010
rect 1363 22954 1431 23010
rect 1487 22954 1555 23010
rect 1611 22954 1679 23010
rect 1735 22954 1803 23010
rect 1859 22954 1927 23010
rect 1983 22954 2051 23010
rect 2107 22954 2117 23010
rect 305 22886 2117 22954
rect 305 22830 315 22886
rect 371 22830 439 22886
rect 495 22830 563 22886
rect 619 22830 687 22886
rect 743 22830 811 22886
rect 867 22830 935 22886
rect 991 22830 1059 22886
rect 1115 22830 1183 22886
rect 1239 22830 1307 22886
rect 1363 22830 1431 22886
rect 1487 22830 1555 22886
rect 1611 22830 1679 22886
rect 1735 22830 1803 22886
rect 1859 22830 1927 22886
rect 1983 22830 2051 22886
rect 2107 22830 2117 22886
rect 305 22762 2117 22830
rect 305 22706 315 22762
rect 371 22706 439 22762
rect 495 22706 563 22762
rect 619 22706 687 22762
rect 743 22706 811 22762
rect 867 22706 935 22762
rect 991 22706 1059 22762
rect 1115 22706 1183 22762
rect 1239 22706 1307 22762
rect 1363 22706 1431 22762
rect 1487 22706 1555 22762
rect 1611 22706 1679 22762
rect 1735 22706 1803 22762
rect 1859 22706 1927 22762
rect 1983 22706 2051 22762
rect 2107 22706 2117 22762
rect 305 22638 2117 22706
rect 305 22582 315 22638
rect 371 22582 439 22638
rect 495 22582 563 22638
rect 619 22582 687 22638
rect 743 22582 811 22638
rect 867 22582 935 22638
rect 991 22582 1059 22638
rect 1115 22582 1183 22638
rect 1239 22582 1307 22638
rect 1363 22582 1431 22638
rect 1487 22582 1555 22638
rect 1611 22582 1679 22638
rect 1735 22582 1803 22638
rect 1859 22582 1927 22638
rect 1983 22582 2051 22638
rect 2107 22582 2117 22638
rect 305 22514 2117 22582
rect 305 22458 315 22514
rect 371 22458 439 22514
rect 495 22458 563 22514
rect 619 22458 687 22514
rect 743 22458 811 22514
rect 867 22458 935 22514
rect 991 22458 1059 22514
rect 1115 22458 1183 22514
rect 1239 22458 1307 22514
rect 1363 22458 1431 22514
rect 1487 22458 1555 22514
rect 1611 22458 1679 22514
rect 1735 22458 1803 22514
rect 1859 22458 1927 22514
rect 1983 22458 2051 22514
rect 2107 22458 2117 22514
rect 305 22390 2117 22458
rect 305 22334 315 22390
rect 371 22334 439 22390
rect 495 22334 563 22390
rect 619 22334 687 22390
rect 743 22334 811 22390
rect 867 22334 935 22390
rect 991 22334 1059 22390
rect 1115 22334 1183 22390
rect 1239 22334 1307 22390
rect 1363 22334 1431 22390
rect 1487 22334 1555 22390
rect 1611 22334 1679 22390
rect 1735 22334 1803 22390
rect 1859 22334 1927 22390
rect 1983 22334 2051 22390
rect 2107 22334 2117 22390
rect 305 22266 2117 22334
rect 305 22210 315 22266
rect 371 22210 439 22266
rect 495 22210 563 22266
rect 619 22210 687 22266
rect 743 22210 811 22266
rect 867 22210 935 22266
rect 991 22210 1059 22266
rect 1115 22210 1183 22266
rect 1239 22210 1307 22266
rect 1363 22210 1431 22266
rect 1487 22210 1555 22266
rect 1611 22210 1679 22266
rect 1735 22210 1803 22266
rect 1859 22210 1927 22266
rect 1983 22210 2051 22266
rect 2107 22210 2117 22266
rect 305 22142 2117 22210
rect 305 22086 315 22142
rect 371 22086 439 22142
rect 495 22086 563 22142
rect 619 22086 687 22142
rect 743 22086 811 22142
rect 867 22086 935 22142
rect 991 22086 1059 22142
rect 1115 22086 1183 22142
rect 1239 22086 1307 22142
rect 1363 22086 1431 22142
rect 1487 22086 1555 22142
rect 1611 22086 1679 22142
rect 1735 22086 1803 22142
rect 1859 22086 1927 22142
rect 1983 22086 2051 22142
rect 2107 22086 2117 22142
rect 305 22018 2117 22086
rect 305 21962 315 22018
rect 371 21962 439 22018
rect 495 21962 563 22018
rect 619 21962 687 22018
rect 743 21962 811 22018
rect 867 21962 935 22018
rect 991 21962 1059 22018
rect 1115 21962 1183 22018
rect 1239 21962 1307 22018
rect 1363 21962 1431 22018
rect 1487 21962 1555 22018
rect 1611 21962 1679 22018
rect 1735 21962 1803 22018
rect 1859 21962 1927 22018
rect 1983 21962 2051 22018
rect 2107 21962 2117 22018
rect 305 21894 2117 21962
rect 305 21838 315 21894
rect 371 21838 439 21894
rect 495 21838 563 21894
rect 619 21838 687 21894
rect 743 21838 811 21894
rect 867 21838 935 21894
rect 991 21838 1059 21894
rect 1115 21838 1183 21894
rect 1239 21838 1307 21894
rect 1363 21838 1431 21894
rect 1487 21838 1555 21894
rect 1611 21838 1679 21894
rect 1735 21838 1803 21894
rect 1859 21838 1927 21894
rect 1983 21838 2051 21894
rect 2107 21838 2117 21894
rect 305 21770 2117 21838
rect 305 21714 315 21770
rect 371 21714 439 21770
rect 495 21714 563 21770
rect 619 21714 687 21770
rect 743 21714 811 21770
rect 867 21714 935 21770
rect 991 21714 1059 21770
rect 1115 21714 1183 21770
rect 1239 21714 1307 21770
rect 1363 21714 1431 21770
rect 1487 21714 1555 21770
rect 1611 21714 1679 21770
rect 1735 21714 1803 21770
rect 1859 21714 1927 21770
rect 1983 21714 2051 21770
rect 2107 21714 2117 21770
rect 305 21646 2117 21714
rect 305 21590 315 21646
rect 371 21590 439 21646
rect 495 21590 563 21646
rect 619 21590 687 21646
rect 743 21590 811 21646
rect 867 21590 935 21646
rect 991 21590 1059 21646
rect 1115 21590 1183 21646
rect 1239 21590 1307 21646
rect 1363 21590 1431 21646
rect 1487 21590 1555 21646
rect 1611 21590 1679 21646
rect 1735 21590 1803 21646
rect 1859 21590 1927 21646
rect 1983 21590 2051 21646
rect 2107 21590 2117 21646
rect 305 21522 2117 21590
rect 305 21466 315 21522
rect 371 21466 439 21522
rect 495 21466 563 21522
rect 619 21466 687 21522
rect 743 21466 811 21522
rect 867 21466 935 21522
rect 991 21466 1059 21522
rect 1115 21466 1183 21522
rect 1239 21466 1307 21522
rect 1363 21466 1431 21522
rect 1487 21466 1555 21522
rect 1611 21466 1679 21522
rect 1735 21466 1803 21522
rect 1859 21466 1927 21522
rect 1983 21466 2051 21522
rect 2107 21466 2117 21522
rect 305 21398 2117 21466
rect 305 21342 315 21398
rect 371 21342 439 21398
rect 495 21342 563 21398
rect 619 21342 687 21398
rect 743 21342 811 21398
rect 867 21342 935 21398
rect 991 21342 1059 21398
rect 1115 21342 1183 21398
rect 1239 21342 1307 21398
rect 1363 21342 1431 21398
rect 1487 21342 1555 21398
rect 1611 21342 1679 21398
rect 1735 21342 1803 21398
rect 1859 21342 1927 21398
rect 1983 21342 2051 21398
rect 2107 21342 2117 21398
rect 305 21274 2117 21342
rect 305 21218 315 21274
rect 371 21218 439 21274
rect 495 21218 563 21274
rect 619 21218 687 21274
rect 743 21218 811 21274
rect 867 21218 935 21274
rect 991 21218 1059 21274
rect 1115 21218 1183 21274
rect 1239 21218 1307 21274
rect 1363 21218 1431 21274
rect 1487 21218 1555 21274
rect 1611 21218 1679 21274
rect 1735 21218 1803 21274
rect 1859 21218 1927 21274
rect 1983 21218 2051 21274
rect 2107 21218 2117 21274
rect 305 21150 2117 21218
rect 305 21094 315 21150
rect 371 21094 439 21150
rect 495 21094 563 21150
rect 619 21094 687 21150
rect 743 21094 811 21150
rect 867 21094 935 21150
rect 991 21094 1059 21150
rect 1115 21094 1183 21150
rect 1239 21094 1307 21150
rect 1363 21094 1431 21150
rect 1487 21094 1555 21150
rect 1611 21094 1679 21150
rect 1735 21094 1803 21150
rect 1859 21094 1927 21150
rect 1983 21094 2051 21150
rect 2107 21094 2117 21150
rect 305 21026 2117 21094
rect 305 20970 315 21026
rect 371 20970 439 21026
rect 495 20970 563 21026
rect 619 20970 687 21026
rect 743 20970 811 21026
rect 867 20970 935 21026
rect 991 20970 1059 21026
rect 1115 20970 1183 21026
rect 1239 20970 1307 21026
rect 1363 20970 1431 21026
rect 1487 20970 1555 21026
rect 1611 20970 1679 21026
rect 1735 20970 1803 21026
rect 1859 20970 1927 21026
rect 1983 20970 2051 21026
rect 2107 20970 2117 21026
rect 305 20902 2117 20970
rect 305 20846 315 20902
rect 371 20846 439 20902
rect 495 20846 563 20902
rect 619 20846 687 20902
rect 743 20846 811 20902
rect 867 20846 935 20902
rect 991 20846 1059 20902
rect 1115 20846 1183 20902
rect 1239 20846 1307 20902
rect 1363 20846 1431 20902
rect 1487 20846 1555 20902
rect 1611 20846 1679 20902
rect 1735 20846 1803 20902
rect 1859 20846 1927 20902
rect 1983 20846 2051 20902
rect 2107 20846 2117 20902
rect 305 20836 2117 20846
rect 2798 23754 4734 23764
rect 2798 23698 2808 23754
rect 2864 23698 2932 23754
rect 2988 23698 3056 23754
rect 3112 23698 3180 23754
rect 3236 23698 3304 23754
rect 3360 23698 3428 23754
rect 3484 23698 3552 23754
rect 3608 23698 3676 23754
rect 3732 23698 3800 23754
rect 3856 23698 3924 23754
rect 3980 23698 4048 23754
rect 4104 23698 4172 23754
rect 4228 23698 4296 23754
rect 4352 23698 4420 23754
rect 4476 23698 4544 23754
rect 4600 23698 4668 23754
rect 4724 23698 4734 23754
rect 2798 23630 4734 23698
rect 2798 23574 2808 23630
rect 2864 23574 2932 23630
rect 2988 23574 3056 23630
rect 3112 23574 3180 23630
rect 3236 23574 3304 23630
rect 3360 23574 3428 23630
rect 3484 23574 3552 23630
rect 3608 23574 3676 23630
rect 3732 23574 3800 23630
rect 3856 23574 3924 23630
rect 3980 23574 4048 23630
rect 4104 23574 4172 23630
rect 4228 23574 4296 23630
rect 4352 23574 4420 23630
rect 4476 23574 4544 23630
rect 4600 23574 4668 23630
rect 4724 23574 4734 23630
rect 2798 23506 4734 23574
rect 2798 23450 2808 23506
rect 2864 23450 2932 23506
rect 2988 23450 3056 23506
rect 3112 23450 3180 23506
rect 3236 23450 3304 23506
rect 3360 23450 3428 23506
rect 3484 23450 3552 23506
rect 3608 23450 3676 23506
rect 3732 23450 3800 23506
rect 3856 23450 3924 23506
rect 3980 23450 4048 23506
rect 4104 23450 4172 23506
rect 4228 23450 4296 23506
rect 4352 23450 4420 23506
rect 4476 23450 4544 23506
rect 4600 23450 4668 23506
rect 4724 23450 4734 23506
rect 2798 23382 4734 23450
rect 2798 23326 2808 23382
rect 2864 23326 2932 23382
rect 2988 23326 3056 23382
rect 3112 23326 3180 23382
rect 3236 23326 3304 23382
rect 3360 23326 3428 23382
rect 3484 23326 3552 23382
rect 3608 23326 3676 23382
rect 3732 23326 3800 23382
rect 3856 23326 3924 23382
rect 3980 23326 4048 23382
rect 4104 23326 4172 23382
rect 4228 23326 4296 23382
rect 4352 23326 4420 23382
rect 4476 23326 4544 23382
rect 4600 23326 4668 23382
rect 4724 23326 4734 23382
rect 2798 23258 4734 23326
rect 2798 23202 2808 23258
rect 2864 23202 2932 23258
rect 2988 23202 3056 23258
rect 3112 23202 3180 23258
rect 3236 23202 3304 23258
rect 3360 23202 3428 23258
rect 3484 23202 3552 23258
rect 3608 23202 3676 23258
rect 3732 23202 3800 23258
rect 3856 23202 3924 23258
rect 3980 23202 4048 23258
rect 4104 23202 4172 23258
rect 4228 23202 4296 23258
rect 4352 23202 4420 23258
rect 4476 23202 4544 23258
rect 4600 23202 4668 23258
rect 4724 23202 4734 23258
rect 2798 23134 4734 23202
rect 2798 23078 2808 23134
rect 2864 23078 2932 23134
rect 2988 23078 3056 23134
rect 3112 23078 3180 23134
rect 3236 23078 3304 23134
rect 3360 23078 3428 23134
rect 3484 23078 3552 23134
rect 3608 23078 3676 23134
rect 3732 23078 3800 23134
rect 3856 23078 3924 23134
rect 3980 23078 4048 23134
rect 4104 23078 4172 23134
rect 4228 23078 4296 23134
rect 4352 23078 4420 23134
rect 4476 23078 4544 23134
rect 4600 23078 4668 23134
rect 4724 23078 4734 23134
rect 2798 23010 4734 23078
rect 2798 22954 2808 23010
rect 2864 22954 2932 23010
rect 2988 22954 3056 23010
rect 3112 22954 3180 23010
rect 3236 22954 3304 23010
rect 3360 22954 3428 23010
rect 3484 22954 3552 23010
rect 3608 22954 3676 23010
rect 3732 22954 3800 23010
rect 3856 22954 3924 23010
rect 3980 22954 4048 23010
rect 4104 22954 4172 23010
rect 4228 22954 4296 23010
rect 4352 22954 4420 23010
rect 4476 22954 4544 23010
rect 4600 22954 4668 23010
rect 4724 22954 4734 23010
rect 2798 22886 4734 22954
rect 2798 22830 2808 22886
rect 2864 22830 2932 22886
rect 2988 22830 3056 22886
rect 3112 22830 3180 22886
rect 3236 22830 3304 22886
rect 3360 22830 3428 22886
rect 3484 22830 3552 22886
rect 3608 22830 3676 22886
rect 3732 22830 3800 22886
rect 3856 22830 3924 22886
rect 3980 22830 4048 22886
rect 4104 22830 4172 22886
rect 4228 22830 4296 22886
rect 4352 22830 4420 22886
rect 4476 22830 4544 22886
rect 4600 22830 4668 22886
rect 4724 22830 4734 22886
rect 2798 22762 4734 22830
rect 2798 22706 2808 22762
rect 2864 22706 2932 22762
rect 2988 22706 3056 22762
rect 3112 22706 3180 22762
rect 3236 22706 3304 22762
rect 3360 22706 3428 22762
rect 3484 22706 3552 22762
rect 3608 22706 3676 22762
rect 3732 22706 3800 22762
rect 3856 22706 3924 22762
rect 3980 22706 4048 22762
rect 4104 22706 4172 22762
rect 4228 22706 4296 22762
rect 4352 22706 4420 22762
rect 4476 22706 4544 22762
rect 4600 22706 4668 22762
rect 4724 22706 4734 22762
rect 2798 22638 4734 22706
rect 2798 22582 2808 22638
rect 2864 22582 2932 22638
rect 2988 22582 3056 22638
rect 3112 22582 3180 22638
rect 3236 22582 3304 22638
rect 3360 22582 3428 22638
rect 3484 22582 3552 22638
rect 3608 22582 3676 22638
rect 3732 22582 3800 22638
rect 3856 22582 3924 22638
rect 3980 22582 4048 22638
rect 4104 22582 4172 22638
rect 4228 22582 4296 22638
rect 4352 22582 4420 22638
rect 4476 22582 4544 22638
rect 4600 22582 4668 22638
rect 4724 22582 4734 22638
rect 2798 22514 4734 22582
rect 2798 22458 2808 22514
rect 2864 22458 2932 22514
rect 2988 22458 3056 22514
rect 3112 22458 3180 22514
rect 3236 22458 3304 22514
rect 3360 22458 3428 22514
rect 3484 22458 3552 22514
rect 3608 22458 3676 22514
rect 3732 22458 3800 22514
rect 3856 22458 3924 22514
rect 3980 22458 4048 22514
rect 4104 22458 4172 22514
rect 4228 22458 4296 22514
rect 4352 22458 4420 22514
rect 4476 22458 4544 22514
rect 4600 22458 4668 22514
rect 4724 22458 4734 22514
rect 2798 22390 4734 22458
rect 2798 22334 2808 22390
rect 2864 22334 2932 22390
rect 2988 22334 3056 22390
rect 3112 22334 3180 22390
rect 3236 22334 3304 22390
rect 3360 22334 3428 22390
rect 3484 22334 3552 22390
rect 3608 22334 3676 22390
rect 3732 22334 3800 22390
rect 3856 22334 3924 22390
rect 3980 22334 4048 22390
rect 4104 22334 4172 22390
rect 4228 22334 4296 22390
rect 4352 22334 4420 22390
rect 4476 22334 4544 22390
rect 4600 22334 4668 22390
rect 4724 22334 4734 22390
rect 2798 22266 4734 22334
rect 2798 22210 2808 22266
rect 2864 22210 2932 22266
rect 2988 22210 3056 22266
rect 3112 22210 3180 22266
rect 3236 22210 3304 22266
rect 3360 22210 3428 22266
rect 3484 22210 3552 22266
rect 3608 22210 3676 22266
rect 3732 22210 3800 22266
rect 3856 22210 3924 22266
rect 3980 22210 4048 22266
rect 4104 22210 4172 22266
rect 4228 22210 4296 22266
rect 4352 22210 4420 22266
rect 4476 22210 4544 22266
rect 4600 22210 4668 22266
rect 4724 22210 4734 22266
rect 2798 22142 4734 22210
rect 2798 22086 2808 22142
rect 2864 22086 2932 22142
rect 2988 22086 3056 22142
rect 3112 22086 3180 22142
rect 3236 22086 3304 22142
rect 3360 22086 3428 22142
rect 3484 22086 3552 22142
rect 3608 22086 3676 22142
rect 3732 22086 3800 22142
rect 3856 22086 3924 22142
rect 3980 22086 4048 22142
rect 4104 22086 4172 22142
rect 4228 22086 4296 22142
rect 4352 22086 4420 22142
rect 4476 22086 4544 22142
rect 4600 22086 4668 22142
rect 4724 22086 4734 22142
rect 2798 22018 4734 22086
rect 2798 21962 2808 22018
rect 2864 21962 2932 22018
rect 2988 21962 3056 22018
rect 3112 21962 3180 22018
rect 3236 21962 3304 22018
rect 3360 21962 3428 22018
rect 3484 21962 3552 22018
rect 3608 21962 3676 22018
rect 3732 21962 3800 22018
rect 3856 21962 3924 22018
rect 3980 21962 4048 22018
rect 4104 21962 4172 22018
rect 4228 21962 4296 22018
rect 4352 21962 4420 22018
rect 4476 21962 4544 22018
rect 4600 21962 4668 22018
rect 4724 21962 4734 22018
rect 2798 21894 4734 21962
rect 2798 21838 2808 21894
rect 2864 21838 2932 21894
rect 2988 21838 3056 21894
rect 3112 21838 3180 21894
rect 3236 21838 3304 21894
rect 3360 21838 3428 21894
rect 3484 21838 3552 21894
rect 3608 21838 3676 21894
rect 3732 21838 3800 21894
rect 3856 21838 3924 21894
rect 3980 21838 4048 21894
rect 4104 21838 4172 21894
rect 4228 21838 4296 21894
rect 4352 21838 4420 21894
rect 4476 21838 4544 21894
rect 4600 21838 4668 21894
rect 4724 21838 4734 21894
rect 2798 21770 4734 21838
rect 2798 21714 2808 21770
rect 2864 21714 2932 21770
rect 2988 21714 3056 21770
rect 3112 21714 3180 21770
rect 3236 21714 3304 21770
rect 3360 21714 3428 21770
rect 3484 21714 3552 21770
rect 3608 21714 3676 21770
rect 3732 21714 3800 21770
rect 3856 21714 3924 21770
rect 3980 21714 4048 21770
rect 4104 21714 4172 21770
rect 4228 21714 4296 21770
rect 4352 21714 4420 21770
rect 4476 21714 4544 21770
rect 4600 21714 4668 21770
rect 4724 21714 4734 21770
rect 2798 21646 4734 21714
rect 2798 21590 2808 21646
rect 2864 21590 2932 21646
rect 2988 21590 3056 21646
rect 3112 21590 3180 21646
rect 3236 21590 3304 21646
rect 3360 21590 3428 21646
rect 3484 21590 3552 21646
rect 3608 21590 3676 21646
rect 3732 21590 3800 21646
rect 3856 21590 3924 21646
rect 3980 21590 4048 21646
rect 4104 21590 4172 21646
rect 4228 21590 4296 21646
rect 4352 21590 4420 21646
rect 4476 21590 4544 21646
rect 4600 21590 4668 21646
rect 4724 21590 4734 21646
rect 2798 21522 4734 21590
rect 2798 21466 2808 21522
rect 2864 21466 2932 21522
rect 2988 21466 3056 21522
rect 3112 21466 3180 21522
rect 3236 21466 3304 21522
rect 3360 21466 3428 21522
rect 3484 21466 3552 21522
rect 3608 21466 3676 21522
rect 3732 21466 3800 21522
rect 3856 21466 3924 21522
rect 3980 21466 4048 21522
rect 4104 21466 4172 21522
rect 4228 21466 4296 21522
rect 4352 21466 4420 21522
rect 4476 21466 4544 21522
rect 4600 21466 4668 21522
rect 4724 21466 4734 21522
rect 2798 21398 4734 21466
rect 2798 21342 2808 21398
rect 2864 21342 2932 21398
rect 2988 21342 3056 21398
rect 3112 21342 3180 21398
rect 3236 21342 3304 21398
rect 3360 21342 3428 21398
rect 3484 21342 3552 21398
rect 3608 21342 3676 21398
rect 3732 21342 3800 21398
rect 3856 21342 3924 21398
rect 3980 21342 4048 21398
rect 4104 21342 4172 21398
rect 4228 21342 4296 21398
rect 4352 21342 4420 21398
rect 4476 21342 4544 21398
rect 4600 21342 4668 21398
rect 4724 21342 4734 21398
rect 2798 21274 4734 21342
rect 2798 21218 2808 21274
rect 2864 21218 2932 21274
rect 2988 21218 3056 21274
rect 3112 21218 3180 21274
rect 3236 21218 3304 21274
rect 3360 21218 3428 21274
rect 3484 21218 3552 21274
rect 3608 21218 3676 21274
rect 3732 21218 3800 21274
rect 3856 21218 3924 21274
rect 3980 21218 4048 21274
rect 4104 21218 4172 21274
rect 4228 21218 4296 21274
rect 4352 21218 4420 21274
rect 4476 21218 4544 21274
rect 4600 21218 4668 21274
rect 4724 21218 4734 21274
rect 2798 21150 4734 21218
rect 2798 21094 2808 21150
rect 2864 21094 2932 21150
rect 2988 21094 3056 21150
rect 3112 21094 3180 21150
rect 3236 21094 3304 21150
rect 3360 21094 3428 21150
rect 3484 21094 3552 21150
rect 3608 21094 3676 21150
rect 3732 21094 3800 21150
rect 3856 21094 3924 21150
rect 3980 21094 4048 21150
rect 4104 21094 4172 21150
rect 4228 21094 4296 21150
rect 4352 21094 4420 21150
rect 4476 21094 4544 21150
rect 4600 21094 4668 21150
rect 4724 21094 4734 21150
rect 2798 21026 4734 21094
rect 2798 20970 2808 21026
rect 2864 20970 2932 21026
rect 2988 20970 3056 21026
rect 3112 20970 3180 21026
rect 3236 20970 3304 21026
rect 3360 20970 3428 21026
rect 3484 20970 3552 21026
rect 3608 20970 3676 21026
rect 3732 20970 3800 21026
rect 3856 20970 3924 21026
rect 3980 20970 4048 21026
rect 4104 20970 4172 21026
rect 4228 20970 4296 21026
rect 4352 20970 4420 21026
rect 4476 20970 4544 21026
rect 4600 20970 4668 21026
rect 4724 20970 4734 21026
rect 2798 20902 4734 20970
rect 2798 20846 2808 20902
rect 2864 20846 2932 20902
rect 2988 20846 3056 20902
rect 3112 20846 3180 20902
rect 3236 20846 3304 20902
rect 3360 20846 3428 20902
rect 3484 20846 3552 20902
rect 3608 20846 3676 20902
rect 3732 20846 3800 20902
rect 3856 20846 3924 20902
rect 3980 20846 4048 20902
rect 4104 20846 4172 20902
rect 4228 20846 4296 20902
rect 4352 20846 4420 20902
rect 4476 20846 4544 20902
rect 4600 20846 4668 20902
rect 4724 20846 4734 20902
rect 2798 20836 4734 20846
rect 5168 23754 7104 23764
rect 5168 23698 5178 23754
rect 5234 23698 5302 23754
rect 5358 23698 5426 23754
rect 5482 23698 5550 23754
rect 5606 23698 5674 23754
rect 5730 23698 5798 23754
rect 5854 23698 5922 23754
rect 5978 23698 6046 23754
rect 6102 23698 6170 23754
rect 6226 23698 6294 23754
rect 6350 23698 6418 23754
rect 6474 23698 6542 23754
rect 6598 23698 6666 23754
rect 6722 23698 6790 23754
rect 6846 23698 6914 23754
rect 6970 23698 7038 23754
rect 7094 23698 7104 23754
rect 5168 23630 7104 23698
rect 5168 23574 5178 23630
rect 5234 23574 5302 23630
rect 5358 23574 5426 23630
rect 5482 23574 5550 23630
rect 5606 23574 5674 23630
rect 5730 23574 5798 23630
rect 5854 23574 5922 23630
rect 5978 23574 6046 23630
rect 6102 23574 6170 23630
rect 6226 23574 6294 23630
rect 6350 23574 6418 23630
rect 6474 23574 6542 23630
rect 6598 23574 6666 23630
rect 6722 23574 6790 23630
rect 6846 23574 6914 23630
rect 6970 23574 7038 23630
rect 7094 23574 7104 23630
rect 5168 23506 7104 23574
rect 5168 23450 5178 23506
rect 5234 23450 5302 23506
rect 5358 23450 5426 23506
rect 5482 23450 5550 23506
rect 5606 23450 5674 23506
rect 5730 23450 5798 23506
rect 5854 23450 5922 23506
rect 5978 23450 6046 23506
rect 6102 23450 6170 23506
rect 6226 23450 6294 23506
rect 6350 23450 6418 23506
rect 6474 23450 6542 23506
rect 6598 23450 6666 23506
rect 6722 23450 6790 23506
rect 6846 23450 6914 23506
rect 6970 23450 7038 23506
rect 7094 23450 7104 23506
rect 5168 23382 7104 23450
rect 5168 23326 5178 23382
rect 5234 23326 5302 23382
rect 5358 23326 5426 23382
rect 5482 23326 5550 23382
rect 5606 23326 5674 23382
rect 5730 23326 5798 23382
rect 5854 23326 5922 23382
rect 5978 23326 6046 23382
rect 6102 23326 6170 23382
rect 6226 23326 6294 23382
rect 6350 23326 6418 23382
rect 6474 23326 6542 23382
rect 6598 23326 6666 23382
rect 6722 23326 6790 23382
rect 6846 23326 6914 23382
rect 6970 23326 7038 23382
rect 7094 23326 7104 23382
rect 5168 23258 7104 23326
rect 5168 23202 5178 23258
rect 5234 23202 5302 23258
rect 5358 23202 5426 23258
rect 5482 23202 5550 23258
rect 5606 23202 5674 23258
rect 5730 23202 5798 23258
rect 5854 23202 5922 23258
rect 5978 23202 6046 23258
rect 6102 23202 6170 23258
rect 6226 23202 6294 23258
rect 6350 23202 6418 23258
rect 6474 23202 6542 23258
rect 6598 23202 6666 23258
rect 6722 23202 6790 23258
rect 6846 23202 6914 23258
rect 6970 23202 7038 23258
rect 7094 23202 7104 23258
rect 5168 23134 7104 23202
rect 5168 23078 5178 23134
rect 5234 23078 5302 23134
rect 5358 23078 5426 23134
rect 5482 23078 5550 23134
rect 5606 23078 5674 23134
rect 5730 23078 5798 23134
rect 5854 23078 5922 23134
rect 5978 23078 6046 23134
rect 6102 23078 6170 23134
rect 6226 23078 6294 23134
rect 6350 23078 6418 23134
rect 6474 23078 6542 23134
rect 6598 23078 6666 23134
rect 6722 23078 6790 23134
rect 6846 23078 6914 23134
rect 6970 23078 7038 23134
rect 7094 23078 7104 23134
rect 5168 23010 7104 23078
rect 5168 22954 5178 23010
rect 5234 22954 5302 23010
rect 5358 22954 5426 23010
rect 5482 22954 5550 23010
rect 5606 22954 5674 23010
rect 5730 22954 5798 23010
rect 5854 22954 5922 23010
rect 5978 22954 6046 23010
rect 6102 22954 6170 23010
rect 6226 22954 6294 23010
rect 6350 22954 6418 23010
rect 6474 22954 6542 23010
rect 6598 22954 6666 23010
rect 6722 22954 6790 23010
rect 6846 22954 6914 23010
rect 6970 22954 7038 23010
rect 7094 22954 7104 23010
rect 5168 22886 7104 22954
rect 5168 22830 5178 22886
rect 5234 22830 5302 22886
rect 5358 22830 5426 22886
rect 5482 22830 5550 22886
rect 5606 22830 5674 22886
rect 5730 22830 5798 22886
rect 5854 22830 5922 22886
rect 5978 22830 6046 22886
rect 6102 22830 6170 22886
rect 6226 22830 6294 22886
rect 6350 22830 6418 22886
rect 6474 22830 6542 22886
rect 6598 22830 6666 22886
rect 6722 22830 6790 22886
rect 6846 22830 6914 22886
rect 6970 22830 7038 22886
rect 7094 22830 7104 22886
rect 5168 22762 7104 22830
rect 5168 22706 5178 22762
rect 5234 22706 5302 22762
rect 5358 22706 5426 22762
rect 5482 22706 5550 22762
rect 5606 22706 5674 22762
rect 5730 22706 5798 22762
rect 5854 22706 5922 22762
rect 5978 22706 6046 22762
rect 6102 22706 6170 22762
rect 6226 22706 6294 22762
rect 6350 22706 6418 22762
rect 6474 22706 6542 22762
rect 6598 22706 6666 22762
rect 6722 22706 6790 22762
rect 6846 22706 6914 22762
rect 6970 22706 7038 22762
rect 7094 22706 7104 22762
rect 5168 22638 7104 22706
rect 5168 22582 5178 22638
rect 5234 22582 5302 22638
rect 5358 22582 5426 22638
rect 5482 22582 5550 22638
rect 5606 22582 5674 22638
rect 5730 22582 5798 22638
rect 5854 22582 5922 22638
rect 5978 22582 6046 22638
rect 6102 22582 6170 22638
rect 6226 22582 6294 22638
rect 6350 22582 6418 22638
rect 6474 22582 6542 22638
rect 6598 22582 6666 22638
rect 6722 22582 6790 22638
rect 6846 22582 6914 22638
rect 6970 22582 7038 22638
rect 7094 22582 7104 22638
rect 5168 22514 7104 22582
rect 5168 22458 5178 22514
rect 5234 22458 5302 22514
rect 5358 22458 5426 22514
rect 5482 22458 5550 22514
rect 5606 22458 5674 22514
rect 5730 22458 5798 22514
rect 5854 22458 5922 22514
rect 5978 22458 6046 22514
rect 6102 22458 6170 22514
rect 6226 22458 6294 22514
rect 6350 22458 6418 22514
rect 6474 22458 6542 22514
rect 6598 22458 6666 22514
rect 6722 22458 6790 22514
rect 6846 22458 6914 22514
rect 6970 22458 7038 22514
rect 7094 22458 7104 22514
rect 5168 22390 7104 22458
rect 5168 22334 5178 22390
rect 5234 22334 5302 22390
rect 5358 22334 5426 22390
rect 5482 22334 5550 22390
rect 5606 22334 5674 22390
rect 5730 22334 5798 22390
rect 5854 22334 5922 22390
rect 5978 22334 6046 22390
rect 6102 22334 6170 22390
rect 6226 22334 6294 22390
rect 6350 22334 6418 22390
rect 6474 22334 6542 22390
rect 6598 22334 6666 22390
rect 6722 22334 6790 22390
rect 6846 22334 6914 22390
rect 6970 22334 7038 22390
rect 7094 22334 7104 22390
rect 5168 22266 7104 22334
rect 5168 22210 5178 22266
rect 5234 22210 5302 22266
rect 5358 22210 5426 22266
rect 5482 22210 5550 22266
rect 5606 22210 5674 22266
rect 5730 22210 5798 22266
rect 5854 22210 5922 22266
rect 5978 22210 6046 22266
rect 6102 22210 6170 22266
rect 6226 22210 6294 22266
rect 6350 22210 6418 22266
rect 6474 22210 6542 22266
rect 6598 22210 6666 22266
rect 6722 22210 6790 22266
rect 6846 22210 6914 22266
rect 6970 22210 7038 22266
rect 7094 22210 7104 22266
rect 5168 22142 7104 22210
rect 5168 22086 5178 22142
rect 5234 22086 5302 22142
rect 5358 22086 5426 22142
rect 5482 22086 5550 22142
rect 5606 22086 5674 22142
rect 5730 22086 5798 22142
rect 5854 22086 5922 22142
rect 5978 22086 6046 22142
rect 6102 22086 6170 22142
rect 6226 22086 6294 22142
rect 6350 22086 6418 22142
rect 6474 22086 6542 22142
rect 6598 22086 6666 22142
rect 6722 22086 6790 22142
rect 6846 22086 6914 22142
rect 6970 22086 7038 22142
rect 7094 22086 7104 22142
rect 5168 22018 7104 22086
rect 5168 21962 5178 22018
rect 5234 21962 5302 22018
rect 5358 21962 5426 22018
rect 5482 21962 5550 22018
rect 5606 21962 5674 22018
rect 5730 21962 5798 22018
rect 5854 21962 5922 22018
rect 5978 21962 6046 22018
rect 6102 21962 6170 22018
rect 6226 21962 6294 22018
rect 6350 21962 6418 22018
rect 6474 21962 6542 22018
rect 6598 21962 6666 22018
rect 6722 21962 6790 22018
rect 6846 21962 6914 22018
rect 6970 21962 7038 22018
rect 7094 21962 7104 22018
rect 5168 21894 7104 21962
rect 5168 21838 5178 21894
rect 5234 21838 5302 21894
rect 5358 21838 5426 21894
rect 5482 21838 5550 21894
rect 5606 21838 5674 21894
rect 5730 21838 5798 21894
rect 5854 21838 5922 21894
rect 5978 21838 6046 21894
rect 6102 21838 6170 21894
rect 6226 21838 6294 21894
rect 6350 21838 6418 21894
rect 6474 21838 6542 21894
rect 6598 21838 6666 21894
rect 6722 21838 6790 21894
rect 6846 21838 6914 21894
rect 6970 21838 7038 21894
rect 7094 21838 7104 21894
rect 5168 21770 7104 21838
rect 5168 21714 5178 21770
rect 5234 21714 5302 21770
rect 5358 21714 5426 21770
rect 5482 21714 5550 21770
rect 5606 21714 5674 21770
rect 5730 21714 5798 21770
rect 5854 21714 5922 21770
rect 5978 21714 6046 21770
rect 6102 21714 6170 21770
rect 6226 21714 6294 21770
rect 6350 21714 6418 21770
rect 6474 21714 6542 21770
rect 6598 21714 6666 21770
rect 6722 21714 6790 21770
rect 6846 21714 6914 21770
rect 6970 21714 7038 21770
rect 7094 21714 7104 21770
rect 5168 21646 7104 21714
rect 5168 21590 5178 21646
rect 5234 21590 5302 21646
rect 5358 21590 5426 21646
rect 5482 21590 5550 21646
rect 5606 21590 5674 21646
rect 5730 21590 5798 21646
rect 5854 21590 5922 21646
rect 5978 21590 6046 21646
rect 6102 21590 6170 21646
rect 6226 21590 6294 21646
rect 6350 21590 6418 21646
rect 6474 21590 6542 21646
rect 6598 21590 6666 21646
rect 6722 21590 6790 21646
rect 6846 21590 6914 21646
rect 6970 21590 7038 21646
rect 7094 21590 7104 21646
rect 5168 21522 7104 21590
rect 5168 21466 5178 21522
rect 5234 21466 5302 21522
rect 5358 21466 5426 21522
rect 5482 21466 5550 21522
rect 5606 21466 5674 21522
rect 5730 21466 5798 21522
rect 5854 21466 5922 21522
rect 5978 21466 6046 21522
rect 6102 21466 6170 21522
rect 6226 21466 6294 21522
rect 6350 21466 6418 21522
rect 6474 21466 6542 21522
rect 6598 21466 6666 21522
rect 6722 21466 6790 21522
rect 6846 21466 6914 21522
rect 6970 21466 7038 21522
rect 7094 21466 7104 21522
rect 5168 21398 7104 21466
rect 5168 21342 5178 21398
rect 5234 21342 5302 21398
rect 5358 21342 5426 21398
rect 5482 21342 5550 21398
rect 5606 21342 5674 21398
rect 5730 21342 5798 21398
rect 5854 21342 5922 21398
rect 5978 21342 6046 21398
rect 6102 21342 6170 21398
rect 6226 21342 6294 21398
rect 6350 21342 6418 21398
rect 6474 21342 6542 21398
rect 6598 21342 6666 21398
rect 6722 21342 6790 21398
rect 6846 21342 6914 21398
rect 6970 21342 7038 21398
rect 7094 21342 7104 21398
rect 5168 21274 7104 21342
rect 5168 21218 5178 21274
rect 5234 21218 5302 21274
rect 5358 21218 5426 21274
rect 5482 21218 5550 21274
rect 5606 21218 5674 21274
rect 5730 21218 5798 21274
rect 5854 21218 5922 21274
rect 5978 21218 6046 21274
rect 6102 21218 6170 21274
rect 6226 21218 6294 21274
rect 6350 21218 6418 21274
rect 6474 21218 6542 21274
rect 6598 21218 6666 21274
rect 6722 21218 6790 21274
rect 6846 21218 6914 21274
rect 6970 21218 7038 21274
rect 7094 21218 7104 21274
rect 5168 21150 7104 21218
rect 5168 21094 5178 21150
rect 5234 21094 5302 21150
rect 5358 21094 5426 21150
rect 5482 21094 5550 21150
rect 5606 21094 5674 21150
rect 5730 21094 5798 21150
rect 5854 21094 5922 21150
rect 5978 21094 6046 21150
rect 6102 21094 6170 21150
rect 6226 21094 6294 21150
rect 6350 21094 6418 21150
rect 6474 21094 6542 21150
rect 6598 21094 6666 21150
rect 6722 21094 6790 21150
rect 6846 21094 6914 21150
rect 6970 21094 7038 21150
rect 7094 21094 7104 21150
rect 5168 21026 7104 21094
rect 5168 20970 5178 21026
rect 5234 20970 5302 21026
rect 5358 20970 5426 21026
rect 5482 20970 5550 21026
rect 5606 20970 5674 21026
rect 5730 20970 5798 21026
rect 5854 20970 5922 21026
rect 5978 20970 6046 21026
rect 6102 20970 6170 21026
rect 6226 20970 6294 21026
rect 6350 20970 6418 21026
rect 6474 20970 6542 21026
rect 6598 20970 6666 21026
rect 6722 20970 6790 21026
rect 6846 20970 6914 21026
rect 6970 20970 7038 21026
rect 7094 20970 7104 21026
rect 5168 20902 7104 20970
rect 5168 20846 5178 20902
rect 5234 20846 5302 20902
rect 5358 20846 5426 20902
rect 5482 20846 5550 20902
rect 5606 20846 5674 20902
rect 5730 20846 5798 20902
rect 5854 20846 5922 20902
rect 5978 20846 6046 20902
rect 6102 20846 6170 20902
rect 6226 20846 6294 20902
rect 6350 20846 6418 20902
rect 6474 20846 6542 20902
rect 6598 20846 6666 20902
rect 6722 20846 6790 20902
rect 6846 20846 6914 20902
rect 6970 20846 7038 20902
rect 7094 20846 7104 20902
rect 5168 20836 7104 20846
rect 7874 23754 9810 23764
rect 7874 23698 7884 23754
rect 7940 23698 8008 23754
rect 8064 23698 8132 23754
rect 8188 23698 8256 23754
rect 8312 23698 8380 23754
rect 8436 23698 8504 23754
rect 8560 23698 8628 23754
rect 8684 23698 8752 23754
rect 8808 23698 8876 23754
rect 8932 23698 9000 23754
rect 9056 23698 9124 23754
rect 9180 23698 9248 23754
rect 9304 23698 9372 23754
rect 9428 23698 9496 23754
rect 9552 23698 9620 23754
rect 9676 23698 9744 23754
rect 9800 23698 9810 23754
rect 7874 23630 9810 23698
rect 7874 23574 7884 23630
rect 7940 23574 8008 23630
rect 8064 23574 8132 23630
rect 8188 23574 8256 23630
rect 8312 23574 8380 23630
rect 8436 23574 8504 23630
rect 8560 23574 8628 23630
rect 8684 23574 8752 23630
rect 8808 23574 8876 23630
rect 8932 23574 9000 23630
rect 9056 23574 9124 23630
rect 9180 23574 9248 23630
rect 9304 23574 9372 23630
rect 9428 23574 9496 23630
rect 9552 23574 9620 23630
rect 9676 23574 9744 23630
rect 9800 23574 9810 23630
rect 7874 23506 9810 23574
rect 7874 23450 7884 23506
rect 7940 23450 8008 23506
rect 8064 23450 8132 23506
rect 8188 23450 8256 23506
rect 8312 23450 8380 23506
rect 8436 23450 8504 23506
rect 8560 23450 8628 23506
rect 8684 23450 8752 23506
rect 8808 23450 8876 23506
rect 8932 23450 9000 23506
rect 9056 23450 9124 23506
rect 9180 23450 9248 23506
rect 9304 23450 9372 23506
rect 9428 23450 9496 23506
rect 9552 23450 9620 23506
rect 9676 23450 9744 23506
rect 9800 23450 9810 23506
rect 7874 23382 9810 23450
rect 7874 23326 7884 23382
rect 7940 23326 8008 23382
rect 8064 23326 8132 23382
rect 8188 23326 8256 23382
rect 8312 23326 8380 23382
rect 8436 23326 8504 23382
rect 8560 23326 8628 23382
rect 8684 23326 8752 23382
rect 8808 23326 8876 23382
rect 8932 23326 9000 23382
rect 9056 23326 9124 23382
rect 9180 23326 9248 23382
rect 9304 23326 9372 23382
rect 9428 23326 9496 23382
rect 9552 23326 9620 23382
rect 9676 23326 9744 23382
rect 9800 23326 9810 23382
rect 7874 23258 9810 23326
rect 7874 23202 7884 23258
rect 7940 23202 8008 23258
rect 8064 23202 8132 23258
rect 8188 23202 8256 23258
rect 8312 23202 8380 23258
rect 8436 23202 8504 23258
rect 8560 23202 8628 23258
rect 8684 23202 8752 23258
rect 8808 23202 8876 23258
rect 8932 23202 9000 23258
rect 9056 23202 9124 23258
rect 9180 23202 9248 23258
rect 9304 23202 9372 23258
rect 9428 23202 9496 23258
rect 9552 23202 9620 23258
rect 9676 23202 9744 23258
rect 9800 23202 9810 23258
rect 7874 23134 9810 23202
rect 7874 23078 7884 23134
rect 7940 23078 8008 23134
rect 8064 23078 8132 23134
rect 8188 23078 8256 23134
rect 8312 23078 8380 23134
rect 8436 23078 8504 23134
rect 8560 23078 8628 23134
rect 8684 23078 8752 23134
rect 8808 23078 8876 23134
rect 8932 23078 9000 23134
rect 9056 23078 9124 23134
rect 9180 23078 9248 23134
rect 9304 23078 9372 23134
rect 9428 23078 9496 23134
rect 9552 23078 9620 23134
rect 9676 23078 9744 23134
rect 9800 23078 9810 23134
rect 7874 23010 9810 23078
rect 7874 22954 7884 23010
rect 7940 22954 8008 23010
rect 8064 22954 8132 23010
rect 8188 22954 8256 23010
rect 8312 22954 8380 23010
rect 8436 22954 8504 23010
rect 8560 22954 8628 23010
rect 8684 22954 8752 23010
rect 8808 22954 8876 23010
rect 8932 22954 9000 23010
rect 9056 22954 9124 23010
rect 9180 22954 9248 23010
rect 9304 22954 9372 23010
rect 9428 22954 9496 23010
rect 9552 22954 9620 23010
rect 9676 22954 9744 23010
rect 9800 22954 9810 23010
rect 7874 22886 9810 22954
rect 7874 22830 7884 22886
rect 7940 22830 8008 22886
rect 8064 22830 8132 22886
rect 8188 22830 8256 22886
rect 8312 22830 8380 22886
rect 8436 22830 8504 22886
rect 8560 22830 8628 22886
rect 8684 22830 8752 22886
rect 8808 22830 8876 22886
rect 8932 22830 9000 22886
rect 9056 22830 9124 22886
rect 9180 22830 9248 22886
rect 9304 22830 9372 22886
rect 9428 22830 9496 22886
rect 9552 22830 9620 22886
rect 9676 22830 9744 22886
rect 9800 22830 9810 22886
rect 7874 22762 9810 22830
rect 7874 22706 7884 22762
rect 7940 22706 8008 22762
rect 8064 22706 8132 22762
rect 8188 22706 8256 22762
rect 8312 22706 8380 22762
rect 8436 22706 8504 22762
rect 8560 22706 8628 22762
rect 8684 22706 8752 22762
rect 8808 22706 8876 22762
rect 8932 22706 9000 22762
rect 9056 22706 9124 22762
rect 9180 22706 9248 22762
rect 9304 22706 9372 22762
rect 9428 22706 9496 22762
rect 9552 22706 9620 22762
rect 9676 22706 9744 22762
rect 9800 22706 9810 22762
rect 7874 22638 9810 22706
rect 7874 22582 7884 22638
rect 7940 22582 8008 22638
rect 8064 22582 8132 22638
rect 8188 22582 8256 22638
rect 8312 22582 8380 22638
rect 8436 22582 8504 22638
rect 8560 22582 8628 22638
rect 8684 22582 8752 22638
rect 8808 22582 8876 22638
rect 8932 22582 9000 22638
rect 9056 22582 9124 22638
rect 9180 22582 9248 22638
rect 9304 22582 9372 22638
rect 9428 22582 9496 22638
rect 9552 22582 9620 22638
rect 9676 22582 9744 22638
rect 9800 22582 9810 22638
rect 7874 22514 9810 22582
rect 7874 22458 7884 22514
rect 7940 22458 8008 22514
rect 8064 22458 8132 22514
rect 8188 22458 8256 22514
rect 8312 22458 8380 22514
rect 8436 22458 8504 22514
rect 8560 22458 8628 22514
rect 8684 22458 8752 22514
rect 8808 22458 8876 22514
rect 8932 22458 9000 22514
rect 9056 22458 9124 22514
rect 9180 22458 9248 22514
rect 9304 22458 9372 22514
rect 9428 22458 9496 22514
rect 9552 22458 9620 22514
rect 9676 22458 9744 22514
rect 9800 22458 9810 22514
rect 7874 22390 9810 22458
rect 7874 22334 7884 22390
rect 7940 22334 8008 22390
rect 8064 22334 8132 22390
rect 8188 22334 8256 22390
rect 8312 22334 8380 22390
rect 8436 22334 8504 22390
rect 8560 22334 8628 22390
rect 8684 22334 8752 22390
rect 8808 22334 8876 22390
rect 8932 22334 9000 22390
rect 9056 22334 9124 22390
rect 9180 22334 9248 22390
rect 9304 22334 9372 22390
rect 9428 22334 9496 22390
rect 9552 22334 9620 22390
rect 9676 22334 9744 22390
rect 9800 22334 9810 22390
rect 7874 22266 9810 22334
rect 7874 22210 7884 22266
rect 7940 22210 8008 22266
rect 8064 22210 8132 22266
rect 8188 22210 8256 22266
rect 8312 22210 8380 22266
rect 8436 22210 8504 22266
rect 8560 22210 8628 22266
rect 8684 22210 8752 22266
rect 8808 22210 8876 22266
rect 8932 22210 9000 22266
rect 9056 22210 9124 22266
rect 9180 22210 9248 22266
rect 9304 22210 9372 22266
rect 9428 22210 9496 22266
rect 9552 22210 9620 22266
rect 9676 22210 9744 22266
rect 9800 22210 9810 22266
rect 7874 22142 9810 22210
rect 7874 22086 7884 22142
rect 7940 22086 8008 22142
rect 8064 22086 8132 22142
rect 8188 22086 8256 22142
rect 8312 22086 8380 22142
rect 8436 22086 8504 22142
rect 8560 22086 8628 22142
rect 8684 22086 8752 22142
rect 8808 22086 8876 22142
rect 8932 22086 9000 22142
rect 9056 22086 9124 22142
rect 9180 22086 9248 22142
rect 9304 22086 9372 22142
rect 9428 22086 9496 22142
rect 9552 22086 9620 22142
rect 9676 22086 9744 22142
rect 9800 22086 9810 22142
rect 7874 22018 9810 22086
rect 7874 21962 7884 22018
rect 7940 21962 8008 22018
rect 8064 21962 8132 22018
rect 8188 21962 8256 22018
rect 8312 21962 8380 22018
rect 8436 21962 8504 22018
rect 8560 21962 8628 22018
rect 8684 21962 8752 22018
rect 8808 21962 8876 22018
rect 8932 21962 9000 22018
rect 9056 21962 9124 22018
rect 9180 21962 9248 22018
rect 9304 21962 9372 22018
rect 9428 21962 9496 22018
rect 9552 21962 9620 22018
rect 9676 21962 9744 22018
rect 9800 21962 9810 22018
rect 7874 21894 9810 21962
rect 7874 21838 7884 21894
rect 7940 21838 8008 21894
rect 8064 21838 8132 21894
rect 8188 21838 8256 21894
rect 8312 21838 8380 21894
rect 8436 21838 8504 21894
rect 8560 21838 8628 21894
rect 8684 21838 8752 21894
rect 8808 21838 8876 21894
rect 8932 21838 9000 21894
rect 9056 21838 9124 21894
rect 9180 21838 9248 21894
rect 9304 21838 9372 21894
rect 9428 21838 9496 21894
rect 9552 21838 9620 21894
rect 9676 21838 9744 21894
rect 9800 21838 9810 21894
rect 7874 21770 9810 21838
rect 7874 21714 7884 21770
rect 7940 21714 8008 21770
rect 8064 21714 8132 21770
rect 8188 21714 8256 21770
rect 8312 21714 8380 21770
rect 8436 21714 8504 21770
rect 8560 21714 8628 21770
rect 8684 21714 8752 21770
rect 8808 21714 8876 21770
rect 8932 21714 9000 21770
rect 9056 21714 9124 21770
rect 9180 21714 9248 21770
rect 9304 21714 9372 21770
rect 9428 21714 9496 21770
rect 9552 21714 9620 21770
rect 9676 21714 9744 21770
rect 9800 21714 9810 21770
rect 7874 21646 9810 21714
rect 7874 21590 7884 21646
rect 7940 21590 8008 21646
rect 8064 21590 8132 21646
rect 8188 21590 8256 21646
rect 8312 21590 8380 21646
rect 8436 21590 8504 21646
rect 8560 21590 8628 21646
rect 8684 21590 8752 21646
rect 8808 21590 8876 21646
rect 8932 21590 9000 21646
rect 9056 21590 9124 21646
rect 9180 21590 9248 21646
rect 9304 21590 9372 21646
rect 9428 21590 9496 21646
rect 9552 21590 9620 21646
rect 9676 21590 9744 21646
rect 9800 21590 9810 21646
rect 7874 21522 9810 21590
rect 7874 21466 7884 21522
rect 7940 21466 8008 21522
rect 8064 21466 8132 21522
rect 8188 21466 8256 21522
rect 8312 21466 8380 21522
rect 8436 21466 8504 21522
rect 8560 21466 8628 21522
rect 8684 21466 8752 21522
rect 8808 21466 8876 21522
rect 8932 21466 9000 21522
rect 9056 21466 9124 21522
rect 9180 21466 9248 21522
rect 9304 21466 9372 21522
rect 9428 21466 9496 21522
rect 9552 21466 9620 21522
rect 9676 21466 9744 21522
rect 9800 21466 9810 21522
rect 7874 21398 9810 21466
rect 7874 21342 7884 21398
rect 7940 21342 8008 21398
rect 8064 21342 8132 21398
rect 8188 21342 8256 21398
rect 8312 21342 8380 21398
rect 8436 21342 8504 21398
rect 8560 21342 8628 21398
rect 8684 21342 8752 21398
rect 8808 21342 8876 21398
rect 8932 21342 9000 21398
rect 9056 21342 9124 21398
rect 9180 21342 9248 21398
rect 9304 21342 9372 21398
rect 9428 21342 9496 21398
rect 9552 21342 9620 21398
rect 9676 21342 9744 21398
rect 9800 21342 9810 21398
rect 7874 21274 9810 21342
rect 7874 21218 7884 21274
rect 7940 21218 8008 21274
rect 8064 21218 8132 21274
rect 8188 21218 8256 21274
rect 8312 21218 8380 21274
rect 8436 21218 8504 21274
rect 8560 21218 8628 21274
rect 8684 21218 8752 21274
rect 8808 21218 8876 21274
rect 8932 21218 9000 21274
rect 9056 21218 9124 21274
rect 9180 21218 9248 21274
rect 9304 21218 9372 21274
rect 9428 21218 9496 21274
rect 9552 21218 9620 21274
rect 9676 21218 9744 21274
rect 9800 21218 9810 21274
rect 7874 21150 9810 21218
rect 7874 21094 7884 21150
rect 7940 21094 8008 21150
rect 8064 21094 8132 21150
rect 8188 21094 8256 21150
rect 8312 21094 8380 21150
rect 8436 21094 8504 21150
rect 8560 21094 8628 21150
rect 8684 21094 8752 21150
rect 8808 21094 8876 21150
rect 8932 21094 9000 21150
rect 9056 21094 9124 21150
rect 9180 21094 9248 21150
rect 9304 21094 9372 21150
rect 9428 21094 9496 21150
rect 9552 21094 9620 21150
rect 9676 21094 9744 21150
rect 9800 21094 9810 21150
rect 7874 21026 9810 21094
rect 7874 20970 7884 21026
rect 7940 20970 8008 21026
rect 8064 20970 8132 21026
rect 8188 20970 8256 21026
rect 8312 20970 8380 21026
rect 8436 20970 8504 21026
rect 8560 20970 8628 21026
rect 8684 20970 8752 21026
rect 8808 20970 8876 21026
rect 8932 20970 9000 21026
rect 9056 20970 9124 21026
rect 9180 20970 9248 21026
rect 9304 20970 9372 21026
rect 9428 20970 9496 21026
rect 9552 20970 9620 21026
rect 9676 20970 9744 21026
rect 9800 20970 9810 21026
rect 7874 20902 9810 20970
rect 7874 20846 7884 20902
rect 7940 20846 8008 20902
rect 8064 20846 8132 20902
rect 8188 20846 8256 20902
rect 8312 20846 8380 20902
rect 8436 20846 8504 20902
rect 8560 20846 8628 20902
rect 8684 20846 8752 20902
rect 8808 20846 8876 20902
rect 8932 20846 9000 20902
rect 9056 20846 9124 20902
rect 9180 20846 9248 20902
rect 9304 20846 9372 20902
rect 9428 20846 9496 20902
rect 9552 20846 9620 20902
rect 9676 20846 9744 20902
rect 9800 20846 9810 20902
rect 7874 20836 9810 20846
rect 10244 23754 12180 23764
rect 10244 23698 10254 23754
rect 10310 23698 10378 23754
rect 10434 23698 10502 23754
rect 10558 23698 10626 23754
rect 10682 23698 10750 23754
rect 10806 23698 10874 23754
rect 10930 23698 10998 23754
rect 11054 23698 11122 23754
rect 11178 23698 11246 23754
rect 11302 23698 11370 23754
rect 11426 23698 11494 23754
rect 11550 23698 11618 23754
rect 11674 23698 11742 23754
rect 11798 23698 11866 23754
rect 11922 23698 11990 23754
rect 12046 23698 12114 23754
rect 12170 23698 12180 23754
rect 10244 23630 12180 23698
rect 10244 23574 10254 23630
rect 10310 23574 10378 23630
rect 10434 23574 10502 23630
rect 10558 23574 10626 23630
rect 10682 23574 10750 23630
rect 10806 23574 10874 23630
rect 10930 23574 10998 23630
rect 11054 23574 11122 23630
rect 11178 23574 11246 23630
rect 11302 23574 11370 23630
rect 11426 23574 11494 23630
rect 11550 23574 11618 23630
rect 11674 23574 11742 23630
rect 11798 23574 11866 23630
rect 11922 23574 11990 23630
rect 12046 23574 12114 23630
rect 12170 23574 12180 23630
rect 10244 23506 12180 23574
rect 10244 23450 10254 23506
rect 10310 23450 10378 23506
rect 10434 23450 10502 23506
rect 10558 23450 10626 23506
rect 10682 23450 10750 23506
rect 10806 23450 10874 23506
rect 10930 23450 10998 23506
rect 11054 23450 11122 23506
rect 11178 23450 11246 23506
rect 11302 23450 11370 23506
rect 11426 23450 11494 23506
rect 11550 23450 11618 23506
rect 11674 23450 11742 23506
rect 11798 23450 11866 23506
rect 11922 23450 11990 23506
rect 12046 23450 12114 23506
rect 12170 23450 12180 23506
rect 10244 23382 12180 23450
rect 10244 23326 10254 23382
rect 10310 23326 10378 23382
rect 10434 23326 10502 23382
rect 10558 23326 10626 23382
rect 10682 23326 10750 23382
rect 10806 23326 10874 23382
rect 10930 23326 10998 23382
rect 11054 23326 11122 23382
rect 11178 23326 11246 23382
rect 11302 23326 11370 23382
rect 11426 23326 11494 23382
rect 11550 23326 11618 23382
rect 11674 23326 11742 23382
rect 11798 23326 11866 23382
rect 11922 23326 11990 23382
rect 12046 23326 12114 23382
rect 12170 23326 12180 23382
rect 10244 23258 12180 23326
rect 10244 23202 10254 23258
rect 10310 23202 10378 23258
rect 10434 23202 10502 23258
rect 10558 23202 10626 23258
rect 10682 23202 10750 23258
rect 10806 23202 10874 23258
rect 10930 23202 10998 23258
rect 11054 23202 11122 23258
rect 11178 23202 11246 23258
rect 11302 23202 11370 23258
rect 11426 23202 11494 23258
rect 11550 23202 11618 23258
rect 11674 23202 11742 23258
rect 11798 23202 11866 23258
rect 11922 23202 11990 23258
rect 12046 23202 12114 23258
rect 12170 23202 12180 23258
rect 10244 23134 12180 23202
rect 10244 23078 10254 23134
rect 10310 23078 10378 23134
rect 10434 23078 10502 23134
rect 10558 23078 10626 23134
rect 10682 23078 10750 23134
rect 10806 23078 10874 23134
rect 10930 23078 10998 23134
rect 11054 23078 11122 23134
rect 11178 23078 11246 23134
rect 11302 23078 11370 23134
rect 11426 23078 11494 23134
rect 11550 23078 11618 23134
rect 11674 23078 11742 23134
rect 11798 23078 11866 23134
rect 11922 23078 11990 23134
rect 12046 23078 12114 23134
rect 12170 23078 12180 23134
rect 10244 23010 12180 23078
rect 10244 22954 10254 23010
rect 10310 22954 10378 23010
rect 10434 22954 10502 23010
rect 10558 22954 10626 23010
rect 10682 22954 10750 23010
rect 10806 22954 10874 23010
rect 10930 22954 10998 23010
rect 11054 22954 11122 23010
rect 11178 22954 11246 23010
rect 11302 22954 11370 23010
rect 11426 22954 11494 23010
rect 11550 22954 11618 23010
rect 11674 22954 11742 23010
rect 11798 22954 11866 23010
rect 11922 22954 11990 23010
rect 12046 22954 12114 23010
rect 12170 22954 12180 23010
rect 10244 22886 12180 22954
rect 10244 22830 10254 22886
rect 10310 22830 10378 22886
rect 10434 22830 10502 22886
rect 10558 22830 10626 22886
rect 10682 22830 10750 22886
rect 10806 22830 10874 22886
rect 10930 22830 10998 22886
rect 11054 22830 11122 22886
rect 11178 22830 11246 22886
rect 11302 22830 11370 22886
rect 11426 22830 11494 22886
rect 11550 22830 11618 22886
rect 11674 22830 11742 22886
rect 11798 22830 11866 22886
rect 11922 22830 11990 22886
rect 12046 22830 12114 22886
rect 12170 22830 12180 22886
rect 10244 22762 12180 22830
rect 10244 22706 10254 22762
rect 10310 22706 10378 22762
rect 10434 22706 10502 22762
rect 10558 22706 10626 22762
rect 10682 22706 10750 22762
rect 10806 22706 10874 22762
rect 10930 22706 10998 22762
rect 11054 22706 11122 22762
rect 11178 22706 11246 22762
rect 11302 22706 11370 22762
rect 11426 22706 11494 22762
rect 11550 22706 11618 22762
rect 11674 22706 11742 22762
rect 11798 22706 11866 22762
rect 11922 22706 11990 22762
rect 12046 22706 12114 22762
rect 12170 22706 12180 22762
rect 10244 22638 12180 22706
rect 10244 22582 10254 22638
rect 10310 22582 10378 22638
rect 10434 22582 10502 22638
rect 10558 22582 10626 22638
rect 10682 22582 10750 22638
rect 10806 22582 10874 22638
rect 10930 22582 10998 22638
rect 11054 22582 11122 22638
rect 11178 22582 11246 22638
rect 11302 22582 11370 22638
rect 11426 22582 11494 22638
rect 11550 22582 11618 22638
rect 11674 22582 11742 22638
rect 11798 22582 11866 22638
rect 11922 22582 11990 22638
rect 12046 22582 12114 22638
rect 12170 22582 12180 22638
rect 10244 22514 12180 22582
rect 10244 22458 10254 22514
rect 10310 22458 10378 22514
rect 10434 22458 10502 22514
rect 10558 22458 10626 22514
rect 10682 22458 10750 22514
rect 10806 22458 10874 22514
rect 10930 22458 10998 22514
rect 11054 22458 11122 22514
rect 11178 22458 11246 22514
rect 11302 22458 11370 22514
rect 11426 22458 11494 22514
rect 11550 22458 11618 22514
rect 11674 22458 11742 22514
rect 11798 22458 11866 22514
rect 11922 22458 11990 22514
rect 12046 22458 12114 22514
rect 12170 22458 12180 22514
rect 10244 22390 12180 22458
rect 10244 22334 10254 22390
rect 10310 22334 10378 22390
rect 10434 22334 10502 22390
rect 10558 22334 10626 22390
rect 10682 22334 10750 22390
rect 10806 22334 10874 22390
rect 10930 22334 10998 22390
rect 11054 22334 11122 22390
rect 11178 22334 11246 22390
rect 11302 22334 11370 22390
rect 11426 22334 11494 22390
rect 11550 22334 11618 22390
rect 11674 22334 11742 22390
rect 11798 22334 11866 22390
rect 11922 22334 11990 22390
rect 12046 22334 12114 22390
rect 12170 22334 12180 22390
rect 10244 22266 12180 22334
rect 10244 22210 10254 22266
rect 10310 22210 10378 22266
rect 10434 22210 10502 22266
rect 10558 22210 10626 22266
rect 10682 22210 10750 22266
rect 10806 22210 10874 22266
rect 10930 22210 10998 22266
rect 11054 22210 11122 22266
rect 11178 22210 11246 22266
rect 11302 22210 11370 22266
rect 11426 22210 11494 22266
rect 11550 22210 11618 22266
rect 11674 22210 11742 22266
rect 11798 22210 11866 22266
rect 11922 22210 11990 22266
rect 12046 22210 12114 22266
rect 12170 22210 12180 22266
rect 10244 22142 12180 22210
rect 10244 22086 10254 22142
rect 10310 22086 10378 22142
rect 10434 22086 10502 22142
rect 10558 22086 10626 22142
rect 10682 22086 10750 22142
rect 10806 22086 10874 22142
rect 10930 22086 10998 22142
rect 11054 22086 11122 22142
rect 11178 22086 11246 22142
rect 11302 22086 11370 22142
rect 11426 22086 11494 22142
rect 11550 22086 11618 22142
rect 11674 22086 11742 22142
rect 11798 22086 11866 22142
rect 11922 22086 11990 22142
rect 12046 22086 12114 22142
rect 12170 22086 12180 22142
rect 10244 22018 12180 22086
rect 10244 21962 10254 22018
rect 10310 21962 10378 22018
rect 10434 21962 10502 22018
rect 10558 21962 10626 22018
rect 10682 21962 10750 22018
rect 10806 21962 10874 22018
rect 10930 21962 10998 22018
rect 11054 21962 11122 22018
rect 11178 21962 11246 22018
rect 11302 21962 11370 22018
rect 11426 21962 11494 22018
rect 11550 21962 11618 22018
rect 11674 21962 11742 22018
rect 11798 21962 11866 22018
rect 11922 21962 11990 22018
rect 12046 21962 12114 22018
rect 12170 21962 12180 22018
rect 10244 21894 12180 21962
rect 10244 21838 10254 21894
rect 10310 21838 10378 21894
rect 10434 21838 10502 21894
rect 10558 21838 10626 21894
rect 10682 21838 10750 21894
rect 10806 21838 10874 21894
rect 10930 21838 10998 21894
rect 11054 21838 11122 21894
rect 11178 21838 11246 21894
rect 11302 21838 11370 21894
rect 11426 21838 11494 21894
rect 11550 21838 11618 21894
rect 11674 21838 11742 21894
rect 11798 21838 11866 21894
rect 11922 21838 11990 21894
rect 12046 21838 12114 21894
rect 12170 21838 12180 21894
rect 10244 21770 12180 21838
rect 10244 21714 10254 21770
rect 10310 21714 10378 21770
rect 10434 21714 10502 21770
rect 10558 21714 10626 21770
rect 10682 21714 10750 21770
rect 10806 21714 10874 21770
rect 10930 21714 10998 21770
rect 11054 21714 11122 21770
rect 11178 21714 11246 21770
rect 11302 21714 11370 21770
rect 11426 21714 11494 21770
rect 11550 21714 11618 21770
rect 11674 21714 11742 21770
rect 11798 21714 11866 21770
rect 11922 21714 11990 21770
rect 12046 21714 12114 21770
rect 12170 21714 12180 21770
rect 10244 21646 12180 21714
rect 10244 21590 10254 21646
rect 10310 21590 10378 21646
rect 10434 21590 10502 21646
rect 10558 21590 10626 21646
rect 10682 21590 10750 21646
rect 10806 21590 10874 21646
rect 10930 21590 10998 21646
rect 11054 21590 11122 21646
rect 11178 21590 11246 21646
rect 11302 21590 11370 21646
rect 11426 21590 11494 21646
rect 11550 21590 11618 21646
rect 11674 21590 11742 21646
rect 11798 21590 11866 21646
rect 11922 21590 11990 21646
rect 12046 21590 12114 21646
rect 12170 21590 12180 21646
rect 10244 21522 12180 21590
rect 10244 21466 10254 21522
rect 10310 21466 10378 21522
rect 10434 21466 10502 21522
rect 10558 21466 10626 21522
rect 10682 21466 10750 21522
rect 10806 21466 10874 21522
rect 10930 21466 10998 21522
rect 11054 21466 11122 21522
rect 11178 21466 11246 21522
rect 11302 21466 11370 21522
rect 11426 21466 11494 21522
rect 11550 21466 11618 21522
rect 11674 21466 11742 21522
rect 11798 21466 11866 21522
rect 11922 21466 11990 21522
rect 12046 21466 12114 21522
rect 12170 21466 12180 21522
rect 10244 21398 12180 21466
rect 10244 21342 10254 21398
rect 10310 21342 10378 21398
rect 10434 21342 10502 21398
rect 10558 21342 10626 21398
rect 10682 21342 10750 21398
rect 10806 21342 10874 21398
rect 10930 21342 10998 21398
rect 11054 21342 11122 21398
rect 11178 21342 11246 21398
rect 11302 21342 11370 21398
rect 11426 21342 11494 21398
rect 11550 21342 11618 21398
rect 11674 21342 11742 21398
rect 11798 21342 11866 21398
rect 11922 21342 11990 21398
rect 12046 21342 12114 21398
rect 12170 21342 12180 21398
rect 10244 21274 12180 21342
rect 10244 21218 10254 21274
rect 10310 21218 10378 21274
rect 10434 21218 10502 21274
rect 10558 21218 10626 21274
rect 10682 21218 10750 21274
rect 10806 21218 10874 21274
rect 10930 21218 10998 21274
rect 11054 21218 11122 21274
rect 11178 21218 11246 21274
rect 11302 21218 11370 21274
rect 11426 21218 11494 21274
rect 11550 21218 11618 21274
rect 11674 21218 11742 21274
rect 11798 21218 11866 21274
rect 11922 21218 11990 21274
rect 12046 21218 12114 21274
rect 12170 21218 12180 21274
rect 10244 21150 12180 21218
rect 10244 21094 10254 21150
rect 10310 21094 10378 21150
rect 10434 21094 10502 21150
rect 10558 21094 10626 21150
rect 10682 21094 10750 21150
rect 10806 21094 10874 21150
rect 10930 21094 10998 21150
rect 11054 21094 11122 21150
rect 11178 21094 11246 21150
rect 11302 21094 11370 21150
rect 11426 21094 11494 21150
rect 11550 21094 11618 21150
rect 11674 21094 11742 21150
rect 11798 21094 11866 21150
rect 11922 21094 11990 21150
rect 12046 21094 12114 21150
rect 12170 21094 12180 21150
rect 10244 21026 12180 21094
rect 10244 20970 10254 21026
rect 10310 20970 10378 21026
rect 10434 20970 10502 21026
rect 10558 20970 10626 21026
rect 10682 20970 10750 21026
rect 10806 20970 10874 21026
rect 10930 20970 10998 21026
rect 11054 20970 11122 21026
rect 11178 20970 11246 21026
rect 11302 20970 11370 21026
rect 11426 20970 11494 21026
rect 11550 20970 11618 21026
rect 11674 20970 11742 21026
rect 11798 20970 11866 21026
rect 11922 20970 11990 21026
rect 12046 20970 12114 21026
rect 12170 20970 12180 21026
rect 10244 20902 12180 20970
rect 10244 20846 10254 20902
rect 10310 20846 10378 20902
rect 10434 20846 10502 20902
rect 10558 20846 10626 20902
rect 10682 20846 10750 20902
rect 10806 20846 10874 20902
rect 10930 20846 10998 20902
rect 11054 20846 11122 20902
rect 11178 20846 11246 20902
rect 11302 20846 11370 20902
rect 11426 20846 11494 20902
rect 11550 20846 11618 20902
rect 11674 20846 11742 20902
rect 11798 20846 11866 20902
rect 11922 20846 11990 20902
rect 12046 20846 12114 20902
rect 12170 20846 12180 20902
rect 10244 20836 12180 20846
rect 12861 23754 14673 23764
rect 12861 23698 12871 23754
rect 12927 23698 12995 23754
rect 13051 23698 13119 23754
rect 13175 23698 13243 23754
rect 13299 23698 13367 23754
rect 13423 23698 13491 23754
rect 13547 23698 13615 23754
rect 13671 23698 13739 23754
rect 13795 23698 13863 23754
rect 13919 23698 13987 23754
rect 14043 23698 14111 23754
rect 14167 23698 14235 23754
rect 14291 23698 14359 23754
rect 14415 23698 14483 23754
rect 14539 23698 14607 23754
rect 14663 23698 14673 23754
rect 12861 23630 14673 23698
rect 12861 23574 12871 23630
rect 12927 23574 12995 23630
rect 13051 23574 13119 23630
rect 13175 23574 13243 23630
rect 13299 23574 13367 23630
rect 13423 23574 13491 23630
rect 13547 23574 13615 23630
rect 13671 23574 13739 23630
rect 13795 23574 13863 23630
rect 13919 23574 13987 23630
rect 14043 23574 14111 23630
rect 14167 23574 14235 23630
rect 14291 23574 14359 23630
rect 14415 23574 14483 23630
rect 14539 23574 14607 23630
rect 14663 23574 14673 23630
rect 12861 23506 14673 23574
rect 12861 23450 12871 23506
rect 12927 23450 12995 23506
rect 13051 23450 13119 23506
rect 13175 23450 13243 23506
rect 13299 23450 13367 23506
rect 13423 23450 13491 23506
rect 13547 23450 13615 23506
rect 13671 23450 13739 23506
rect 13795 23450 13863 23506
rect 13919 23450 13987 23506
rect 14043 23450 14111 23506
rect 14167 23450 14235 23506
rect 14291 23450 14359 23506
rect 14415 23450 14483 23506
rect 14539 23450 14607 23506
rect 14663 23450 14673 23506
rect 12861 23382 14673 23450
rect 12861 23326 12871 23382
rect 12927 23326 12995 23382
rect 13051 23326 13119 23382
rect 13175 23326 13243 23382
rect 13299 23326 13367 23382
rect 13423 23326 13491 23382
rect 13547 23326 13615 23382
rect 13671 23326 13739 23382
rect 13795 23326 13863 23382
rect 13919 23326 13987 23382
rect 14043 23326 14111 23382
rect 14167 23326 14235 23382
rect 14291 23326 14359 23382
rect 14415 23326 14483 23382
rect 14539 23326 14607 23382
rect 14663 23326 14673 23382
rect 12861 23258 14673 23326
rect 12861 23202 12871 23258
rect 12927 23202 12995 23258
rect 13051 23202 13119 23258
rect 13175 23202 13243 23258
rect 13299 23202 13367 23258
rect 13423 23202 13491 23258
rect 13547 23202 13615 23258
rect 13671 23202 13739 23258
rect 13795 23202 13863 23258
rect 13919 23202 13987 23258
rect 14043 23202 14111 23258
rect 14167 23202 14235 23258
rect 14291 23202 14359 23258
rect 14415 23202 14483 23258
rect 14539 23202 14607 23258
rect 14663 23202 14673 23258
rect 12861 23134 14673 23202
rect 12861 23078 12871 23134
rect 12927 23078 12995 23134
rect 13051 23078 13119 23134
rect 13175 23078 13243 23134
rect 13299 23078 13367 23134
rect 13423 23078 13491 23134
rect 13547 23078 13615 23134
rect 13671 23078 13739 23134
rect 13795 23078 13863 23134
rect 13919 23078 13987 23134
rect 14043 23078 14111 23134
rect 14167 23078 14235 23134
rect 14291 23078 14359 23134
rect 14415 23078 14483 23134
rect 14539 23078 14607 23134
rect 14663 23078 14673 23134
rect 12861 23010 14673 23078
rect 12861 22954 12871 23010
rect 12927 22954 12995 23010
rect 13051 22954 13119 23010
rect 13175 22954 13243 23010
rect 13299 22954 13367 23010
rect 13423 22954 13491 23010
rect 13547 22954 13615 23010
rect 13671 22954 13739 23010
rect 13795 22954 13863 23010
rect 13919 22954 13987 23010
rect 14043 22954 14111 23010
rect 14167 22954 14235 23010
rect 14291 22954 14359 23010
rect 14415 22954 14483 23010
rect 14539 22954 14607 23010
rect 14663 22954 14673 23010
rect 12861 22886 14673 22954
rect 12861 22830 12871 22886
rect 12927 22830 12995 22886
rect 13051 22830 13119 22886
rect 13175 22830 13243 22886
rect 13299 22830 13367 22886
rect 13423 22830 13491 22886
rect 13547 22830 13615 22886
rect 13671 22830 13739 22886
rect 13795 22830 13863 22886
rect 13919 22830 13987 22886
rect 14043 22830 14111 22886
rect 14167 22830 14235 22886
rect 14291 22830 14359 22886
rect 14415 22830 14483 22886
rect 14539 22830 14607 22886
rect 14663 22830 14673 22886
rect 12861 22762 14673 22830
rect 12861 22706 12871 22762
rect 12927 22706 12995 22762
rect 13051 22706 13119 22762
rect 13175 22706 13243 22762
rect 13299 22706 13367 22762
rect 13423 22706 13491 22762
rect 13547 22706 13615 22762
rect 13671 22706 13739 22762
rect 13795 22706 13863 22762
rect 13919 22706 13987 22762
rect 14043 22706 14111 22762
rect 14167 22706 14235 22762
rect 14291 22706 14359 22762
rect 14415 22706 14483 22762
rect 14539 22706 14607 22762
rect 14663 22706 14673 22762
rect 12861 22638 14673 22706
rect 12861 22582 12871 22638
rect 12927 22582 12995 22638
rect 13051 22582 13119 22638
rect 13175 22582 13243 22638
rect 13299 22582 13367 22638
rect 13423 22582 13491 22638
rect 13547 22582 13615 22638
rect 13671 22582 13739 22638
rect 13795 22582 13863 22638
rect 13919 22582 13987 22638
rect 14043 22582 14111 22638
rect 14167 22582 14235 22638
rect 14291 22582 14359 22638
rect 14415 22582 14483 22638
rect 14539 22582 14607 22638
rect 14663 22582 14673 22638
rect 12861 22514 14673 22582
rect 12861 22458 12871 22514
rect 12927 22458 12995 22514
rect 13051 22458 13119 22514
rect 13175 22458 13243 22514
rect 13299 22458 13367 22514
rect 13423 22458 13491 22514
rect 13547 22458 13615 22514
rect 13671 22458 13739 22514
rect 13795 22458 13863 22514
rect 13919 22458 13987 22514
rect 14043 22458 14111 22514
rect 14167 22458 14235 22514
rect 14291 22458 14359 22514
rect 14415 22458 14483 22514
rect 14539 22458 14607 22514
rect 14663 22458 14673 22514
rect 12861 22390 14673 22458
rect 12861 22334 12871 22390
rect 12927 22334 12995 22390
rect 13051 22334 13119 22390
rect 13175 22334 13243 22390
rect 13299 22334 13367 22390
rect 13423 22334 13491 22390
rect 13547 22334 13615 22390
rect 13671 22334 13739 22390
rect 13795 22334 13863 22390
rect 13919 22334 13987 22390
rect 14043 22334 14111 22390
rect 14167 22334 14235 22390
rect 14291 22334 14359 22390
rect 14415 22334 14483 22390
rect 14539 22334 14607 22390
rect 14663 22334 14673 22390
rect 12861 22266 14673 22334
rect 12861 22210 12871 22266
rect 12927 22210 12995 22266
rect 13051 22210 13119 22266
rect 13175 22210 13243 22266
rect 13299 22210 13367 22266
rect 13423 22210 13491 22266
rect 13547 22210 13615 22266
rect 13671 22210 13739 22266
rect 13795 22210 13863 22266
rect 13919 22210 13987 22266
rect 14043 22210 14111 22266
rect 14167 22210 14235 22266
rect 14291 22210 14359 22266
rect 14415 22210 14483 22266
rect 14539 22210 14607 22266
rect 14663 22210 14673 22266
rect 12861 22142 14673 22210
rect 12861 22086 12871 22142
rect 12927 22086 12995 22142
rect 13051 22086 13119 22142
rect 13175 22086 13243 22142
rect 13299 22086 13367 22142
rect 13423 22086 13491 22142
rect 13547 22086 13615 22142
rect 13671 22086 13739 22142
rect 13795 22086 13863 22142
rect 13919 22086 13987 22142
rect 14043 22086 14111 22142
rect 14167 22086 14235 22142
rect 14291 22086 14359 22142
rect 14415 22086 14483 22142
rect 14539 22086 14607 22142
rect 14663 22086 14673 22142
rect 12861 22018 14673 22086
rect 12861 21962 12871 22018
rect 12927 21962 12995 22018
rect 13051 21962 13119 22018
rect 13175 21962 13243 22018
rect 13299 21962 13367 22018
rect 13423 21962 13491 22018
rect 13547 21962 13615 22018
rect 13671 21962 13739 22018
rect 13795 21962 13863 22018
rect 13919 21962 13987 22018
rect 14043 21962 14111 22018
rect 14167 21962 14235 22018
rect 14291 21962 14359 22018
rect 14415 21962 14483 22018
rect 14539 21962 14607 22018
rect 14663 21962 14673 22018
rect 12861 21894 14673 21962
rect 12861 21838 12871 21894
rect 12927 21838 12995 21894
rect 13051 21838 13119 21894
rect 13175 21838 13243 21894
rect 13299 21838 13367 21894
rect 13423 21838 13491 21894
rect 13547 21838 13615 21894
rect 13671 21838 13739 21894
rect 13795 21838 13863 21894
rect 13919 21838 13987 21894
rect 14043 21838 14111 21894
rect 14167 21838 14235 21894
rect 14291 21838 14359 21894
rect 14415 21838 14483 21894
rect 14539 21838 14607 21894
rect 14663 21838 14673 21894
rect 12861 21770 14673 21838
rect 12861 21714 12871 21770
rect 12927 21714 12995 21770
rect 13051 21714 13119 21770
rect 13175 21714 13243 21770
rect 13299 21714 13367 21770
rect 13423 21714 13491 21770
rect 13547 21714 13615 21770
rect 13671 21714 13739 21770
rect 13795 21714 13863 21770
rect 13919 21714 13987 21770
rect 14043 21714 14111 21770
rect 14167 21714 14235 21770
rect 14291 21714 14359 21770
rect 14415 21714 14483 21770
rect 14539 21714 14607 21770
rect 14663 21714 14673 21770
rect 12861 21646 14673 21714
rect 12861 21590 12871 21646
rect 12927 21590 12995 21646
rect 13051 21590 13119 21646
rect 13175 21590 13243 21646
rect 13299 21590 13367 21646
rect 13423 21590 13491 21646
rect 13547 21590 13615 21646
rect 13671 21590 13739 21646
rect 13795 21590 13863 21646
rect 13919 21590 13987 21646
rect 14043 21590 14111 21646
rect 14167 21590 14235 21646
rect 14291 21590 14359 21646
rect 14415 21590 14483 21646
rect 14539 21590 14607 21646
rect 14663 21590 14673 21646
rect 12861 21522 14673 21590
rect 12861 21466 12871 21522
rect 12927 21466 12995 21522
rect 13051 21466 13119 21522
rect 13175 21466 13243 21522
rect 13299 21466 13367 21522
rect 13423 21466 13491 21522
rect 13547 21466 13615 21522
rect 13671 21466 13739 21522
rect 13795 21466 13863 21522
rect 13919 21466 13987 21522
rect 14043 21466 14111 21522
rect 14167 21466 14235 21522
rect 14291 21466 14359 21522
rect 14415 21466 14483 21522
rect 14539 21466 14607 21522
rect 14663 21466 14673 21522
rect 12861 21398 14673 21466
rect 12861 21342 12871 21398
rect 12927 21342 12995 21398
rect 13051 21342 13119 21398
rect 13175 21342 13243 21398
rect 13299 21342 13367 21398
rect 13423 21342 13491 21398
rect 13547 21342 13615 21398
rect 13671 21342 13739 21398
rect 13795 21342 13863 21398
rect 13919 21342 13987 21398
rect 14043 21342 14111 21398
rect 14167 21342 14235 21398
rect 14291 21342 14359 21398
rect 14415 21342 14483 21398
rect 14539 21342 14607 21398
rect 14663 21342 14673 21398
rect 12861 21274 14673 21342
rect 12861 21218 12871 21274
rect 12927 21218 12995 21274
rect 13051 21218 13119 21274
rect 13175 21218 13243 21274
rect 13299 21218 13367 21274
rect 13423 21218 13491 21274
rect 13547 21218 13615 21274
rect 13671 21218 13739 21274
rect 13795 21218 13863 21274
rect 13919 21218 13987 21274
rect 14043 21218 14111 21274
rect 14167 21218 14235 21274
rect 14291 21218 14359 21274
rect 14415 21218 14483 21274
rect 14539 21218 14607 21274
rect 14663 21218 14673 21274
rect 12861 21150 14673 21218
rect 12861 21094 12871 21150
rect 12927 21094 12995 21150
rect 13051 21094 13119 21150
rect 13175 21094 13243 21150
rect 13299 21094 13367 21150
rect 13423 21094 13491 21150
rect 13547 21094 13615 21150
rect 13671 21094 13739 21150
rect 13795 21094 13863 21150
rect 13919 21094 13987 21150
rect 14043 21094 14111 21150
rect 14167 21094 14235 21150
rect 14291 21094 14359 21150
rect 14415 21094 14483 21150
rect 14539 21094 14607 21150
rect 14663 21094 14673 21150
rect 12861 21026 14673 21094
rect 12861 20970 12871 21026
rect 12927 20970 12995 21026
rect 13051 20970 13119 21026
rect 13175 20970 13243 21026
rect 13299 20970 13367 21026
rect 13423 20970 13491 21026
rect 13547 20970 13615 21026
rect 13671 20970 13739 21026
rect 13795 20970 13863 21026
rect 13919 20970 13987 21026
rect 14043 20970 14111 21026
rect 14167 20970 14235 21026
rect 14291 20970 14359 21026
rect 14415 20970 14483 21026
rect 14539 20970 14607 21026
rect 14663 20970 14673 21026
rect 12861 20902 14673 20970
rect 12861 20846 12871 20902
rect 12927 20846 12995 20902
rect 13051 20846 13119 20902
rect 13175 20846 13243 20902
rect 13299 20846 13367 20902
rect 13423 20846 13491 20902
rect 13547 20846 13615 20902
rect 13671 20846 13739 20902
rect 13795 20846 13863 20902
rect 13919 20846 13987 20902
rect 14043 20846 14111 20902
rect 14167 20846 14235 20902
rect 14291 20846 14359 20902
rect 14415 20846 14483 20902
rect 14539 20846 14607 20902
rect 14663 20846 14673 20902
rect 12861 20836 14673 20846
rect 305 20554 2117 20564
rect 305 20498 315 20554
rect 371 20498 439 20554
rect 495 20498 563 20554
rect 619 20498 687 20554
rect 743 20498 811 20554
rect 867 20498 935 20554
rect 991 20498 1059 20554
rect 1115 20498 1183 20554
rect 1239 20498 1307 20554
rect 1363 20498 1431 20554
rect 1487 20498 1555 20554
rect 1611 20498 1679 20554
rect 1735 20498 1803 20554
rect 1859 20498 1927 20554
rect 1983 20498 2051 20554
rect 2107 20498 2117 20554
rect 305 20430 2117 20498
rect 305 20374 315 20430
rect 371 20374 439 20430
rect 495 20374 563 20430
rect 619 20374 687 20430
rect 743 20374 811 20430
rect 867 20374 935 20430
rect 991 20374 1059 20430
rect 1115 20374 1183 20430
rect 1239 20374 1307 20430
rect 1363 20374 1431 20430
rect 1487 20374 1555 20430
rect 1611 20374 1679 20430
rect 1735 20374 1803 20430
rect 1859 20374 1927 20430
rect 1983 20374 2051 20430
rect 2107 20374 2117 20430
rect 305 20306 2117 20374
rect 305 20250 315 20306
rect 371 20250 439 20306
rect 495 20250 563 20306
rect 619 20250 687 20306
rect 743 20250 811 20306
rect 867 20250 935 20306
rect 991 20250 1059 20306
rect 1115 20250 1183 20306
rect 1239 20250 1307 20306
rect 1363 20250 1431 20306
rect 1487 20250 1555 20306
rect 1611 20250 1679 20306
rect 1735 20250 1803 20306
rect 1859 20250 1927 20306
rect 1983 20250 2051 20306
rect 2107 20250 2117 20306
rect 305 20182 2117 20250
rect 305 20126 315 20182
rect 371 20126 439 20182
rect 495 20126 563 20182
rect 619 20126 687 20182
rect 743 20126 811 20182
rect 867 20126 935 20182
rect 991 20126 1059 20182
rect 1115 20126 1183 20182
rect 1239 20126 1307 20182
rect 1363 20126 1431 20182
rect 1487 20126 1555 20182
rect 1611 20126 1679 20182
rect 1735 20126 1803 20182
rect 1859 20126 1927 20182
rect 1983 20126 2051 20182
rect 2107 20126 2117 20182
rect 305 20058 2117 20126
rect 305 20002 315 20058
rect 371 20002 439 20058
rect 495 20002 563 20058
rect 619 20002 687 20058
rect 743 20002 811 20058
rect 867 20002 935 20058
rect 991 20002 1059 20058
rect 1115 20002 1183 20058
rect 1239 20002 1307 20058
rect 1363 20002 1431 20058
rect 1487 20002 1555 20058
rect 1611 20002 1679 20058
rect 1735 20002 1803 20058
rect 1859 20002 1927 20058
rect 1983 20002 2051 20058
rect 2107 20002 2117 20058
rect 305 19934 2117 20002
rect 305 19878 315 19934
rect 371 19878 439 19934
rect 495 19878 563 19934
rect 619 19878 687 19934
rect 743 19878 811 19934
rect 867 19878 935 19934
rect 991 19878 1059 19934
rect 1115 19878 1183 19934
rect 1239 19878 1307 19934
rect 1363 19878 1431 19934
rect 1487 19878 1555 19934
rect 1611 19878 1679 19934
rect 1735 19878 1803 19934
rect 1859 19878 1927 19934
rect 1983 19878 2051 19934
rect 2107 19878 2117 19934
rect 305 19810 2117 19878
rect 305 19754 315 19810
rect 371 19754 439 19810
rect 495 19754 563 19810
rect 619 19754 687 19810
rect 743 19754 811 19810
rect 867 19754 935 19810
rect 991 19754 1059 19810
rect 1115 19754 1183 19810
rect 1239 19754 1307 19810
rect 1363 19754 1431 19810
rect 1487 19754 1555 19810
rect 1611 19754 1679 19810
rect 1735 19754 1803 19810
rect 1859 19754 1927 19810
rect 1983 19754 2051 19810
rect 2107 19754 2117 19810
rect 305 19686 2117 19754
rect 305 19630 315 19686
rect 371 19630 439 19686
rect 495 19630 563 19686
rect 619 19630 687 19686
rect 743 19630 811 19686
rect 867 19630 935 19686
rect 991 19630 1059 19686
rect 1115 19630 1183 19686
rect 1239 19630 1307 19686
rect 1363 19630 1431 19686
rect 1487 19630 1555 19686
rect 1611 19630 1679 19686
rect 1735 19630 1803 19686
rect 1859 19630 1927 19686
rect 1983 19630 2051 19686
rect 2107 19630 2117 19686
rect 305 19562 2117 19630
rect 305 19506 315 19562
rect 371 19506 439 19562
rect 495 19506 563 19562
rect 619 19506 687 19562
rect 743 19506 811 19562
rect 867 19506 935 19562
rect 991 19506 1059 19562
rect 1115 19506 1183 19562
rect 1239 19506 1307 19562
rect 1363 19506 1431 19562
rect 1487 19506 1555 19562
rect 1611 19506 1679 19562
rect 1735 19506 1803 19562
rect 1859 19506 1927 19562
rect 1983 19506 2051 19562
rect 2107 19506 2117 19562
rect 305 19438 2117 19506
rect 305 19382 315 19438
rect 371 19382 439 19438
rect 495 19382 563 19438
rect 619 19382 687 19438
rect 743 19382 811 19438
rect 867 19382 935 19438
rect 991 19382 1059 19438
rect 1115 19382 1183 19438
rect 1239 19382 1307 19438
rect 1363 19382 1431 19438
rect 1487 19382 1555 19438
rect 1611 19382 1679 19438
rect 1735 19382 1803 19438
rect 1859 19382 1927 19438
rect 1983 19382 2051 19438
rect 2107 19382 2117 19438
rect 305 19314 2117 19382
rect 305 19258 315 19314
rect 371 19258 439 19314
rect 495 19258 563 19314
rect 619 19258 687 19314
rect 743 19258 811 19314
rect 867 19258 935 19314
rect 991 19258 1059 19314
rect 1115 19258 1183 19314
rect 1239 19258 1307 19314
rect 1363 19258 1431 19314
rect 1487 19258 1555 19314
rect 1611 19258 1679 19314
rect 1735 19258 1803 19314
rect 1859 19258 1927 19314
rect 1983 19258 2051 19314
rect 2107 19258 2117 19314
rect 305 19190 2117 19258
rect 305 19134 315 19190
rect 371 19134 439 19190
rect 495 19134 563 19190
rect 619 19134 687 19190
rect 743 19134 811 19190
rect 867 19134 935 19190
rect 991 19134 1059 19190
rect 1115 19134 1183 19190
rect 1239 19134 1307 19190
rect 1363 19134 1431 19190
rect 1487 19134 1555 19190
rect 1611 19134 1679 19190
rect 1735 19134 1803 19190
rect 1859 19134 1927 19190
rect 1983 19134 2051 19190
rect 2107 19134 2117 19190
rect 305 19066 2117 19134
rect 305 19010 315 19066
rect 371 19010 439 19066
rect 495 19010 563 19066
rect 619 19010 687 19066
rect 743 19010 811 19066
rect 867 19010 935 19066
rect 991 19010 1059 19066
rect 1115 19010 1183 19066
rect 1239 19010 1307 19066
rect 1363 19010 1431 19066
rect 1487 19010 1555 19066
rect 1611 19010 1679 19066
rect 1735 19010 1803 19066
rect 1859 19010 1927 19066
rect 1983 19010 2051 19066
rect 2107 19010 2117 19066
rect 305 18942 2117 19010
rect 305 18886 315 18942
rect 371 18886 439 18942
rect 495 18886 563 18942
rect 619 18886 687 18942
rect 743 18886 811 18942
rect 867 18886 935 18942
rect 991 18886 1059 18942
rect 1115 18886 1183 18942
rect 1239 18886 1307 18942
rect 1363 18886 1431 18942
rect 1487 18886 1555 18942
rect 1611 18886 1679 18942
rect 1735 18886 1803 18942
rect 1859 18886 1927 18942
rect 1983 18886 2051 18942
rect 2107 18886 2117 18942
rect 305 18818 2117 18886
rect 305 18762 315 18818
rect 371 18762 439 18818
rect 495 18762 563 18818
rect 619 18762 687 18818
rect 743 18762 811 18818
rect 867 18762 935 18818
rect 991 18762 1059 18818
rect 1115 18762 1183 18818
rect 1239 18762 1307 18818
rect 1363 18762 1431 18818
rect 1487 18762 1555 18818
rect 1611 18762 1679 18818
rect 1735 18762 1803 18818
rect 1859 18762 1927 18818
rect 1983 18762 2051 18818
rect 2107 18762 2117 18818
rect 305 18694 2117 18762
rect 305 18638 315 18694
rect 371 18638 439 18694
rect 495 18638 563 18694
rect 619 18638 687 18694
rect 743 18638 811 18694
rect 867 18638 935 18694
rect 991 18638 1059 18694
rect 1115 18638 1183 18694
rect 1239 18638 1307 18694
rect 1363 18638 1431 18694
rect 1487 18638 1555 18694
rect 1611 18638 1679 18694
rect 1735 18638 1803 18694
rect 1859 18638 1927 18694
rect 1983 18638 2051 18694
rect 2107 18638 2117 18694
rect 305 18570 2117 18638
rect 305 18514 315 18570
rect 371 18514 439 18570
rect 495 18514 563 18570
rect 619 18514 687 18570
rect 743 18514 811 18570
rect 867 18514 935 18570
rect 991 18514 1059 18570
rect 1115 18514 1183 18570
rect 1239 18514 1307 18570
rect 1363 18514 1431 18570
rect 1487 18514 1555 18570
rect 1611 18514 1679 18570
rect 1735 18514 1803 18570
rect 1859 18514 1927 18570
rect 1983 18514 2051 18570
rect 2107 18514 2117 18570
rect 305 18446 2117 18514
rect 305 18390 315 18446
rect 371 18390 439 18446
rect 495 18390 563 18446
rect 619 18390 687 18446
rect 743 18390 811 18446
rect 867 18390 935 18446
rect 991 18390 1059 18446
rect 1115 18390 1183 18446
rect 1239 18390 1307 18446
rect 1363 18390 1431 18446
rect 1487 18390 1555 18446
rect 1611 18390 1679 18446
rect 1735 18390 1803 18446
rect 1859 18390 1927 18446
rect 1983 18390 2051 18446
rect 2107 18390 2117 18446
rect 305 18322 2117 18390
rect 305 18266 315 18322
rect 371 18266 439 18322
rect 495 18266 563 18322
rect 619 18266 687 18322
rect 743 18266 811 18322
rect 867 18266 935 18322
rect 991 18266 1059 18322
rect 1115 18266 1183 18322
rect 1239 18266 1307 18322
rect 1363 18266 1431 18322
rect 1487 18266 1555 18322
rect 1611 18266 1679 18322
rect 1735 18266 1803 18322
rect 1859 18266 1927 18322
rect 1983 18266 2051 18322
rect 2107 18266 2117 18322
rect 305 18198 2117 18266
rect 305 18142 315 18198
rect 371 18142 439 18198
rect 495 18142 563 18198
rect 619 18142 687 18198
rect 743 18142 811 18198
rect 867 18142 935 18198
rect 991 18142 1059 18198
rect 1115 18142 1183 18198
rect 1239 18142 1307 18198
rect 1363 18142 1431 18198
rect 1487 18142 1555 18198
rect 1611 18142 1679 18198
rect 1735 18142 1803 18198
rect 1859 18142 1927 18198
rect 1983 18142 2051 18198
rect 2107 18142 2117 18198
rect 305 18074 2117 18142
rect 305 18018 315 18074
rect 371 18018 439 18074
rect 495 18018 563 18074
rect 619 18018 687 18074
rect 743 18018 811 18074
rect 867 18018 935 18074
rect 991 18018 1059 18074
rect 1115 18018 1183 18074
rect 1239 18018 1307 18074
rect 1363 18018 1431 18074
rect 1487 18018 1555 18074
rect 1611 18018 1679 18074
rect 1735 18018 1803 18074
rect 1859 18018 1927 18074
rect 1983 18018 2051 18074
rect 2107 18018 2117 18074
rect 305 17950 2117 18018
rect 305 17894 315 17950
rect 371 17894 439 17950
rect 495 17894 563 17950
rect 619 17894 687 17950
rect 743 17894 811 17950
rect 867 17894 935 17950
rect 991 17894 1059 17950
rect 1115 17894 1183 17950
rect 1239 17894 1307 17950
rect 1363 17894 1431 17950
rect 1487 17894 1555 17950
rect 1611 17894 1679 17950
rect 1735 17894 1803 17950
rect 1859 17894 1927 17950
rect 1983 17894 2051 17950
rect 2107 17894 2117 17950
rect 305 17826 2117 17894
rect 305 17770 315 17826
rect 371 17770 439 17826
rect 495 17770 563 17826
rect 619 17770 687 17826
rect 743 17770 811 17826
rect 867 17770 935 17826
rect 991 17770 1059 17826
rect 1115 17770 1183 17826
rect 1239 17770 1307 17826
rect 1363 17770 1431 17826
rect 1487 17770 1555 17826
rect 1611 17770 1679 17826
rect 1735 17770 1803 17826
rect 1859 17770 1927 17826
rect 1983 17770 2051 17826
rect 2107 17770 2117 17826
rect 305 17702 2117 17770
rect 305 17646 315 17702
rect 371 17646 439 17702
rect 495 17646 563 17702
rect 619 17646 687 17702
rect 743 17646 811 17702
rect 867 17646 935 17702
rect 991 17646 1059 17702
rect 1115 17646 1183 17702
rect 1239 17646 1307 17702
rect 1363 17646 1431 17702
rect 1487 17646 1555 17702
rect 1611 17646 1679 17702
rect 1735 17646 1803 17702
rect 1859 17646 1927 17702
rect 1983 17646 2051 17702
rect 2107 17646 2117 17702
rect 305 17636 2117 17646
rect 2798 20554 4734 20564
rect 2798 20498 2808 20554
rect 2864 20498 2932 20554
rect 2988 20498 3056 20554
rect 3112 20498 3180 20554
rect 3236 20498 3304 20554
rect 3360 20498 3428 20554
rect 3484 20498 3552 20554
rect 3608 20498 3676 20554
rect 3732 20498 3800 20554
rect 3856 20498 3924 20554
rect 3980 20498 4048 20554
rect 4104 20498 4172 20554
rect 4228 20498 4296 20554
rect 4352 20498 4420 20554
rect 4476 20498 4544 20554
rect 4600 20498 4668 20554
rect 4724 20498 4734 20554
rect 2798 20430 4734 20498
rect 2798 20374 2808 20430
rect 2864 20374 2932 20430
rect 2988 20374 3056 20430
rect 3112 20374 3180 20430
rect 3236 20374 3304 20430
rect 3360 20374 3428 20430
rect 3484 20374 3552 20430
rect 3608 20374 3676 20430
rect 3732 20374 3800 20430
rect 3856 20374 3924 20430
rect 3980 20374 4048 20430
rect 4104 20374 4172 20430
rect 4228 20374 4296 20430
rect 4352 20374 4420 20430
rect 4476 20374 4544 20430
rect 4600 20374 4668 20430
rect 4724 20374 4734 20430
rect 2798 20306 4734 20374
rect 2798 20250 2808 20306
rect 2864 20250 2932 20306
rect 2988 20250 3056 20306
rect 3112 20250 3180 20306
rect 3236 20250 3304 20306
rect 3360 20250 3428 20306
rect 3484 20250 3552 20306
rect 3608 20250 3676 20306
rect 3732 20250 3800 20306
rect 3856 20250 3924 20306
rect 3980 20250 4048 20306
rect 4104 20250 4172 20306
rect 4228 20250 4296 20306
rect 4352 20250 4420 20306
rect 4476 20250 4544 20306
rect 4600 20250 4668 20306
rect 4724 20250 4734 20306
rect 2798 20182 4734 20250
rect 2798 20126 2808 20182
rect 2864 20126 2932 20182
rect 2988 20126 3056 20182
rect 3112 20126 3180 20182
rect 3236 20126 3304 20182
rect 3360 20126 3428 20182
rect 3484 20126 3552 20182
rect 3608 20126 3676 20182
rect 3732 20126 3800 20182
rect 3856 20126 3924 20182
rect 3980 20126 4048 20182
rect 4104 20126 4172 20182
rect 4228 20126 4296 20182
rect 4352 20126 4420 20182
rect 4476 20126 4544 20182
rect 4600 20126 4668 20182
rect 4724 20126 4734 20182
rect 2798 20058 4734 20126
rect 2798 20002 2808 20058
rect 2864 20002 2932 20058
rect 2988 20002 3056 20058
rect 3112 20002 3180 20058
rect 3236 20002 3304 20058
rect 3360 20002 3428 20058
rect 3484 20002 3552 20058
rect 3608 20002 3676 20058
rect 3732 20002 3800 20058
rect 3856 20002 3924 20058
rect 3980 20002 4048 20058
rect 4104 20002 4172 20058
rect 4228 20002 4296 20058
rect 4352 20002 4420 20058
rect 4476 20002 4544 20058
rect 4600 20002 4668 20058
rect 4724 20002 4734 20058
rect 2798 19934 4734 20002
rect 2798 19878 2808 19934
rect 2864 19878 2932 19934
rect 2988 19878 3056 19934
rect 3112 19878 3180 19934
rect 3236 19878 3304 19934
rect 3360 19878 3428 19934
rect 3484 19878 3552 19934
rect 3608 19878 3676 19934
rect 3732 19878 3800 19934
rect 3856 19878 3924 19934
rect 3980 19878 4048 19934
rect 4104 19878 4172 19934
rect 4228 19878 4296 19934
rect 4352 19878 4420 19934
rect 4476 19878 4544 19934
rect 4600 19878 4668 19934
rect 4724 19878 4734 19934
rect 2798 19810 4734 19878
rect 2798 19754 2808 19810
rect 2864 19754 2932 19810
rect 2988 19754 3056 19810
rect 3112 19754 3180 19810
rect 3236 19754 3304 19810
rect 3360 19754 3428 19810
rect 3484 19754 3552 19810
rect 3608 19754 3676 19810
rect 3732 19754 3800 19810
rect 3856 19754 3924 19810
rect 3980 19754 4048 19810
rect 4104 19754 4172 19810
rect 4228 19754 4296 19810
rect 4352 19754 4420 19810
rect 4476 19754 4544 19810
rect 4600 19754 4668 19810
rect 4724 19754 4734 19810
rect 2798 19686 4734 19754
rect 2798 19630 2808 19686
rect 2864 19630 2932 19686
rect 2988 19630 3056 19686
rect 3112 19630 3180 19686
rect 3236 19630 3304 19686
rect 3360 19630 3428 19686
rect 3484 19630 3552 19686
rect 3608 19630 3676 19686
rect 3732 19630 3800 19686
rect 3856 19630 3924 19686
rect 3980 19630 4048 19686
rect 4104 19630 4172 19686
rect 4228 19630 4296 19686
rect 4352 19630 4420 19686
rect 4476 19630 4544 19686
rect 4600 19630 4668 19686
rect 4724 19630 4734 19686
rect 2798 19562 4734 19630
rect 2798 19506 2808 19562
rect 2864 19506 2932 19562
rect 2988 19506 3056 19562
rect 3112 19506 3180 19562
rect 3236 19506 3304 19562
rect 3360 19506 3428 19562
rect 3484 19506 3552 19562
rect 3608 19506 3676 19562
rect 3732 19506 3800 19562
rect 3856 19506 3924 19562
rect 3980 19506 4048 19562
rect 4104 19506 4172 19562
rect 4228 19506 4296 19562
rect 4352 19506 4420 19562
rect 4476 19506 4544 19562
rect 4600 19506 4668 19562
rect 4724 19506 4734 19562
rect 2798 19438 4734 19506
rect 2798 19382 2808 19438
rect 2864 19382 2932 19438
rect 2988 19382 3056 19438
rect 3112 19382 3180 19438
rect 3236 19382 3304 19438
rect 3360 19382 3428 19438
rect 3484 19382 3552 19438
rect 3608 19382 3676 19438
rect 3732 19382 3800 19438
rect 3856 19382 3924 19438
rect 3980 19382 4048 19438
rect 4104 19382 4172 19438
rect 4228 19382 4296 19438
rect 4352 19382 4420 19438
rect 4476 19382 4544 19438
rect 4600 19382 4668 19438
rect 4724 19382 4734 19438
rect 2798 19314 4734 19382
rect 2798 19258 2808 19314
rect 2864 19258 2932 19314
rect 2988 19258 3056 19314
rect 3112 19258 3180 19314
rect 3236 19258 3304 19314
rect 3360 19258 3428 19314
rect 3484 19258 3552 19314
rect 3608 19258 3676 19314
rect 3732 19258 3800 19314
rect 3856 19258 3924 19314
rect 3980 19258 4048 19314
rect 4104 19258 4172 19314
rect 4228 19258 4296 19314
rect 4352 19258 4420 19314
rect 4476 19258 4544 19314
rect 4600 19258 4668 19314
rect 4724 19258 4734 19314
rect 2798 19190 4734 19258
rect 2798 19134 2808 19190
rect 2864 19134 2932 19190
rect 2988 19134 3056 19190
rect 3112 19134 3180 19190
rect 3236 19134 3304 19190
rect 3360 19134 3428 19190
rect 3484 19134 3552 19190
rect 3608 19134 3676 19190
rect 3732 19134 3800 19190
rect 3856 19134 3924 19190
rect 3980 19134 4048 19190
rect 4104 19134 4172 19190
rect 4228 19134 4296 19190
rect 4352 19134 4420 19190
rect 4476 19134 4544 19190
rect 4600 19134 4668 19190
rect 4724 19134 4734 19190
rect 2798 19066 4734 19134
rect 2798 19010 2808 19066
rect 2864 19010 2932 19066
rect 2988 19010 3056 19066
rect 3112 19010 3180 19066
rect 3236 19010 3304 19066
rect 3360 19010 3428 19066
rect 3484 19010 3552 19066
rect 3608 19010 3676 19066
rect 3732 19010 3800 19066
rect 3856 19010 3924 19066
rect 3980 19010 4048 19066
rect 4104 19010 4172 19066
rect 4228 19010 4296 19066
rect 4352 19010 4420 19066
rect 4476 19010 4544 19066
rect 4600 19010 4668 19066
rect 4724 19010 4734 19066
rect 2798 18942 4734 19010
rect 2798 18886 2808 18942
rect 2864 18886 2932 18942
rect 2988 18886 3056 18942
rect 3112 18886 3180 18942
rect 3236 18886 3304 18942
rect 3360 18886 3428 18942
rect 3484 18886 3552 18942
rect 3608 18886 3676 18942
rect 3732 18886 3800 18942
rect 3856 18886 3924 18942
rect 3980 18886 4048 18942
rect 4104 18886 4172 18942
rect 4228 18886 4296 18942
rect 4352 18886 4420 18942
rect 4476 18886 4544 18942
rect 4600 18886 4668 18942
rect 4724 18886 4734 18942
rect 2798 18818 4734 18886
rect 2798 18762 2808 18818
rect 2864 18762 2932 18818
rect 2988 18762 3056 18818
rect 3112 18762 3180 18818
rect 3236 18762 3304 18818
rect 3360 18762 3428 18818
rect 3484 18762 3552 18818
rect 3608 18762 3676 18818
rect 3732 18762 3800 18818
rect 3856 18762 3924 18818
rect 3980 18762 4048 18818
rect 4104 18762 4172 18818
rect 4228 18762 4296 18818
rect 4352 18762 4420 18818
rect 4476 18762 4544 18818
rect 4600 18762 4668 18818
rect 4724 18762 4734 18818
rect 2798 18694 4734 18762
rect 2798 18638 2808 18694
rect 2864 18638 2932 18694
rect 2988 18638 3056 18694
rect 3112 18638 3180 18694
rect 3236 18638 3304 18694
rect 3360 18638 3428 18694
rect 3484 18638 3552 18694
rect 3608 18638 3676 18694
rect 3732 18638 3800 18694
rect 3856 18638 3924 18694
rect 3980 18638 4048 18694
rect 4104 18638 4172 18694
rect 4228 18638 4296 18694
rect 4352 18638 4420 18694
rect 4476 18638 4544 18694
rect 4600 18638 4668 18694
rect 4724 18638 4734 18694
rect 2798 18570 4734 18638
rect 2798 18514 2808 18570
rect 2864 18514 2932 18570
rect 2988 18514 3056 18570
rect 3112 18514 3180 18570
rect 3236 18514 3304 18570
rect 3360 18514 3428 18570
rect 3484 18514 3552 18570
rect 3608 18514 3676 18570
rect 3732 18514 3800 18570
rect 3856 18514 3924 18570
rect 3980 18514 4048 18570
rect 4104 18514 4172 18570
rect 4228 18514 4296 18570
rect 4352 18514 4420 18570
rect 4476 18514 4544 18570
rect 4600 18514 4668 18570
rect 4724 18514 4734 18570
rect 2798 18446 4734 18514
rect 2798 18390 2808 18446
rect 2864 18390 2932 18446
rect 2988 18390 3056 18446
rect 3112 18390 3180 18446
rect 3236 18390 3304 18446
rect 3360 18390 3428 18446
rect 3484 18390 3552 18446
rect 3608 18390 3676 18446
rect 3732 18390 3800 18446
rect 3856 18390 3924 18446
rect 3980 18390 4048 18446
rect 4104 18390 4172 18446
rect 4228 18390 4296 18446
rect 4352 18390 4420 18446
rect 4476 18390 4544 18446
rect 4600 18390 4668 18446
rect 4724 18390 4734 18446
rect 2798 18322 4734 18390
rect 2798 18266 2808 18322
rect 2864 18266 2932 18322
rect 2988 18266 3056 18322
rect 3112 18266 3180 18322
rect 3236 18266 3304 18322
rect 3360 18266 3428 18322
rect 3484 18266 3552 18322
rect 3608 18266 3676 18322
rect 3732 18266 3800 18322
rect 3856 18266 3924 18322
rect 3980 18266 4048 18322
rect 4104 18266 4172 18322
rect 4228 18266 4296 18322
rect 4352 18266 4420 18322
rect 4476 18266 4544 18322
rect 4600 18266 4668 18322
rect 4724 18266 4734 18322
rect 2798 18198 4734 18266
rect 2798 18142 2808 18198
rect 2864 18142 2932 18198
rect 2988 18142 3056 18198
rect 3112 18142 3180 18198
rect 3236 18142 3304 18198
rect 3360 18142 3428 18198
rect 3484 18142 3552 18198
rect 3608 18142 3676 18198
rect 3732 18142 3800 18198
rect 3856 18142 3924 18198
rect 3980 18142 4048 18198
rect 4104 18142 4172 18198
rect 4228 18142 4296 18198
rect 4352 18142 4420 18198
rect 4476 18142 4544 18198
rect 4600 18142 4668 18198
rect 4724 18142 4734 18198
rect 2798 18074 4734 18142
rect 2798 18018 2808 18074
rect 2864 18018 2932 18074
rect 2988 18018 3056 18074
rect 3112 18018 3180 18074
rect 3236 18018 3304 18074
rect 3360 18018 3428 18074
rect 3484 18018 3552 18074
rect 3608 18018 3676 18074
rect 3732 18018 3800 18074
rect 3856 18018 3924 18074
rect 3980 18018 4048 18074
rect 4104 18018 4172 18074
rect 4228 18018 4296 18074
rect 4352 18018 4420 18074
rect 4476 18018 4544 18074
rect 4600 18018 4668 18074
rect 4724 18018 4734 18074
rect 2798 17950 4734 18018
rect 2798 17894 2808 17950
rect 2864 17894 2932 17950
rect 2988 17894 3056 17950
rect 3112 17894 3180 17950
rect 3236 17894 3304 17950
rect 3360 17894 3428 17950
rect 3484 17894 3552 17950
rect 3608 17894 3676 17950
rect 3732 17894 3800 17950
rect 3856 17894 3924 17950
rect 3980 17894 4048 17950
rect 4104 17894 4172 17950
rect 4228 17894 4296 17950
rect 4352 17894 4420 17950
rect 4476 17894 4544 17950
rect 4600 17894 4668 17950
rect 4724 17894 4734 17950
rect 2798 17826 4734 17894
rect 2798 17770 2808 17826
rect 2864 17770 2932 17826
rect 2988 17770 3056 17826
rect 3112 17770 3180 17826
rect 3236 17770 3304 17826
rect 3360 17770 3428 17826
rect 3484 17770 3552 17826
rect 3608 17770 3676 17826
rect 3732 17770 3800 17826
rect 3856 17770 3924 17826
rect 3980 17770 4048 17826
rect 4104 17770 4172 17826
rect 4228 17770 4296 17826
rect 4352 17770 4420 17826
rect 4476 17770 4544 17826
rect 4600 17770 4668 17826
rect 4724 17770 4734 17826
rect 2798 17702 4734 17770
rect 2798 17646 2808 17702
rect 2864 17646 2932 17702
rect 2988 17646 3056 17702
rect 3112 17646 3180 17702
rect 3236 17646 3304 17702
rect 3360 17646 3428 17702
rect 3484 17646 3552 17702
rect 3608 17646 3676 17702
rect 3732 17646 3800 17702
rect 3856 17646 3924 17702
rect 3980 17646 4048 17702
rect 4104 17646 4172 17702
rect 4228 17646 4296 17702
rect 4352 17646 4420 17702
rect 4476 17646 4544 17702
rect 4600 17646 4668 17702
rect 4724 17646 4734 17702
rect 2798 17636 4734 17646
rect 5168 20554 7104 20564
rect 5168 20498 5178 20554
rect 5234 20498 5302 20554
rect 5358 20498 5426 20554
rect 5482 20498 5550 20554
rect 5606 20498 5674 20554
rect 5730 20498 5798 20554
rect 5854 20498 5922 20554
rect 5978 20498 6046 20554
rect 6102 20498 6170 20554
rect 6226 20498 6294 20554
rect 6350 20498 6418 20554
rect 6474 20498 6542 20554
rect 6598 20498 6666 20554
rect 6722 20498 6790 20554
rect 6846 20498 6914 20554
rect 6970 20498 7038 20554
rect 7094 20498 7104 20554
rect 5168 20430 7104 20498
rect 5168 20374 5178 20430
rect 5234 20374 5302 20430
rect 5358 20374 5426 20430
rect 5482 20374 5550 20430
rect 5606 20374 5674 20430
rect 5730 20374 5798 20430
rect 5854 20374 5922 20430
rect 5978 20374 6046 20430
rect 6102 20374 6170 20430
rect 6226 20374 6294 20430
rect 6350 20374 6418 20430
rect 6474 20374 6542 20430
rect 6598 20374 6666 20430
rect 6722 20374 6790 20430
rect 6846 20374 6914 20430
rect 6970 20374 7038 20430
rect 7094 20374 7104 20430
rect 5168 20306 7104 20374
rect 5168 20250 5178 20306
rect 5234 20250 5302 20306
rect 5358 20250 5426 20306
rect 5482 20250 5550 20306
rect 5606 20250 5674 20306
rect 5730 20250 5798 20306
rect 5854 20250 5922 20306
rect 5978 20250 6046 20306
rect 6102 20250 6170 20306
rect 6226 20250 6294 20306
rect 6350 20250 6418 20306
rect 6474 20250 6542 20306
rect 6598 20250 6666 20306
rect 6722 20250 6790 20306
rect 6846 20250 6914 20306
rect 6970 20250 7038 20306
rect 7094 20250 7104 20306
rect 5168 20182 7104 20250
rect 5168 20126 5178 20182
rect 5234 20126 5302 20182
rect 5358 20126 5426 20182
rect 5482 20126 5550 20182
rect 5606 20126 5674 20182
rect 5730 20126 5798 20182
rect 5854 20126 5922 20182
rect 5978 20126 6046 20182
rect 6102 20126 6170 20182
rect 6226 20126 6294 20182
rect 6350 20126 6418 20182
rect 6474 20126 6542 20182
rect 6598 20126 6666 20182
rect 6722 20126 6790 20182
rect 6846 20126 6914 20182
rect 6970 20126 7038 20182
rect 7094 20126 7104 20182
rect 5168 20058 7104 20126
rect 5168 20002 5178 20058
rect 5234 20002 5302 20058
rect 5358 20002 5426 20058
rect 5482 20002 5550 20058
rect 5606 20002 5674 20058
rect 5730 20002 5798 20058
rect 5854 20002 5922 20058
rect 5978 20002 6046 20058
rect 6102 20002 6170 20058
rect 6226 20002 6294 20058
rect 6350 20002 6418 20058
rect 6474 20002 6542 20058
rect 6598 20002 6666 20058
rect 6722 20002 6790 20058
rect 6846 20002 6914 20058
rect 6970 20002 7038 20058
rect 7094 20002 7104 20058
rect 5168 19934 7104 20002
rect 5168 19878 5178 19934
rect 5234 19878 5302 19934
rect 5358 19878 5426 19934
rect 5482 19878 5550 19934
rect 5606 19878 5674 19934
rect 5730 19878 5798 19934
rect 5854 19878 5922 19934
rect 5978 19878 6046 19934
rect 6102 19878 6170 19934
rect 6226 19878 6294 19934
rect 6350 19878 6418 19934
rect 6474 19878 6542 19934
rect 6598 19878 6666 19934
rect 6722 19878 6790 19934
rect 6846 19878 6914 19934
rect 6970 19878 7038 19934
rect 7094 19878 7104 19934
rect 5168 19810 7104 19878
rect 5168 19754 5178 19810
rect 5234 19754 5302 19810
rect 5358 19754 5426 19810
rect 5482 19754 5550 19810
rect 5606 19754 5674 19810
rect 5730 19754 5798 19810
rect 5854 19754 5922 19810
rect 5978 19754 6046 19810
rect 6102 19754 6170 19810
rect 6226 19754 6294 19810
rect 6350 19754 6418 19810
rect 6474 19754 6542 19810
rect 6598 19754 6666 19810
rect 6722 19754 6790 19810
rect 6846 19754 6914 19810
rect 6970 19754 7038 19810
rect 7094 19754 7104 19810
rect 5168 19686 7104 19754
rect 5168 19630 5178 19686
rect 5234 19630 5302 19686
rect 5358 19630 5426 19686
rect 5482 19630 5550 19686
rect 5606 19630 5674 19686
rect 5730 19630 5798 19686
rect 5854 19630 5922 19686
rect 5978 19630 6046 19686
rect 6102 19630 6170 19686
rect 6226 19630 6294 19686
rect 6350 19630 6418 19686
rect 6474 19630 6542 19686
rect 6598 19630 6666 19686
rect 6722 19630 6790 19686
rect 6846 19630 6914 19686
rect 6970 19630 7038 19686
rect 7094 19630 7104 19686
rect 5168 19562 7104 19630
rect 5168 19506 5178 19562
rect 5234 19506 5302 19562
rect 5358 19506 5426 19562
rect 5482 19506 5550 19562
rect 5606 19506 5674 19562
rect 5730 19506 5798 19562
rect 5854 19506 5922 19562
rect 5978 19506 6046 19562
rect 6102 19506 6170 19562
rect 6226 19506 6294 19562
rect 6350 19506 6418 19562
rect 6474 19506 6542 19562
rect 6598 19506 6666 19562
rect 6722 19506 6790 19562
rect 6846 19506 6914 19562
rect 6970 19506 7038 19562
rect 7094 19506 7104 19562
rect 5168 19438 7104 19506
rect 5168 19382 5178 19438
rect 5234 19382 5302 19438
rect 5358 19382 5426 19438
rect 5482 19382 5550 19438
rect 5606 19382 5674 19438
rect 5730 19382 5798 19438
rect 5854 19382 5922 19438
rect 5978 19382 6046 19438
rect 6102 19382 6170 19438
rect 6226 19382 6294 19438
rect 6350 19382 6418 19438
rect 6474 19382 6542 19438
rect 6598 19382 6666 19438
rect 6722 19382 6790 19438
rect 6846 19382 6914 19438
rect 6970 19382 7038 19438
rect 7094 19382 7104 19438
rect 5168 19314 7104 19382
rect 5168 19258 5178 19314
rect 5234 19258 5302 19314
rect 5358 19258 5426 19314
rect 5482 19258 5550 19314
rect 5606 19258 5674 19314
rect 5730 19258 5798 19314
rect 5854 19258 5922 19314
rect 5978 19258 6046 19314
rect 6102 19258 6170 19314
rect 6226 19258 6294 19314
rect 6350 19258 6418 19314
rect 6474 19258 6542 19314
rect 6598 19258 6666 19314
rect 6722 19258 6790 19314
rect 6846 19258 6914 19314
rect 6970 19258 7038 19314
rect 7094 19258 7104 19314
rect 5168 19190 7104 19258
rect 5168 19134 5178 19190
rect 5234 19134 5302 19190
rect 5358 19134 5426 19190
rect 5482 19134 5550 19190
rect 5606 19134 5674 19190
rect 5730 19134 5798 19190
rect 5854 19134 5922 19190
rect 5978 19134 6046 19190
rect 6102 19134 6170 19190
rect 6226 19134 6294 19190
rect 6350 19134 6418 19190
rect 6474 19134 6542 19190
rect 6598 19134 6666 19190
rect 6722 19134 6790 19190
rect 6846 19134 6914 19190
rect 6970 19134 7038 19190
rect 7094 19134 7104 19190
rect 5168 19066 7104 19134
rect 5168 19010 5178 19066
rect 5234 19010 5302 19066
rect 5358 19010 5426 19066
rect 5482 19010 5550 19066
rect 5606 19010 5674 19066
rect 5730 19010 5798 19066
rect 5854 19010 5922 19066
rect 5978 19010 6046 19066
rect 6102 19010 6170 19066
rect 6226 19010 6294 19066
rect 6350 19010 6418 19066
rect 6474 19010 6542 19066
rect 6598 19010 6666 19066
rect 6722 19010 6790 19066
rect 6846 19010 6914 19066
rect 6970 19010 7038 19066
rect 7094 19010 7104 19066
rect 5168 18942 7104 19010
rect 5168 18886 5178 18942
rect 5234 18886 5302 18942
rect 5358 18886 5426 18942
rect 5482 18886 5550 18942
rect 5606 18886 5674 18942
rect 5730 18886 5798 18942
rect 5854 18886 5922 18942
rect 5978 18886 6046 18942
rect 6102 18886 6170 18942
rect 6226 18886 6294 18942
rect 6350 18886 6418 18942
rect 6474 18886 6542 18942
rect 6598 18886 6666 18942
rect 6722 18886 6790 18942
rect 6846 18886 6914 18942
rect 6970 18886 7038 18942
rect 7094 18886 7104 18942
rect 5168 18818 7104 18886
rect 5168 18762 5178 18818
rect 5234 18762 5302 18818
rect 5358 18762 5426 18818
rect 5482 18762 5550 18818
rect 5606 18762 5674 18818
rect 5730 18762 5798 18818
rect 5854 18762 5922 18818
rect 5978 18762 6046 18818
rect 6102 18762 6170 18818
rect 6226 18762 6294 18818
rect 6350 18762 6418 18818
rect 6474 18762 6542 18818
rect 6598 18762 6666 18818
rect 6722 18762 6790 18818
rect 6846 18762 6914 18818
rect 6970 18762 7038 18818
rect 7094 18762 7104 18818
rect 5168 18694 7104 18762
rect 5168 18638 5178 18694
rect 5234 18638 5302 18694
rect 5358 18638 5426 18694
rect 5482 18638 5550 18694
rect 5606 18638 5674 18694
rect 5730 18638 5798 18694
rect 5854 18638 5922 18694
rect 5978 18638 6046 18694
rect 6102 18638 6170 18694
rect 6226 18638 6294 18694
rect 6350 18638 6418 18694
rect 6474 18638 6542 18694
rect 6598 18638 6666 18694
rect 6722 18638 6790 18694
rect 6846 18638 6914 18694
rect 6970 18638 7038 18694
rect 7094 18638 7104 18694
rect 5168 18570 7104 18638
rect 5168 18514 5178 18570
rect 5234 18514 5302 18570
rect 5358 18514 5426 18570
rect 5482 18514 5550 18570
rect 5606 18514 5674 18570
rect 5730 18514 5798 18570
rect 5854 18514 5922 18570
rect 5978 18514 6046 18570
rect 6102 18514 6170 18570
rect 6226 18514 6294 18570
rect 6350 18514 6418 18570
rect 6474 18514 6542 18570
rect 6598 18514 6666 18570
rect 6722 18514 6790 18570
rect 6846 18514 6914 18570
rect 6970 18514 7038 18570
rect 7094 18514 7104 18570
rect 5168 18446 7104 18514
rect 5168 18390 5178 18446
rect 5234 18390 5302 18446
rect 5358 18390 5426 18446
rect 5482 18390 5550 18446
rect 5606 18390 5674 18446
rect 5730 18390 5798 18446
rect 5854 18390 5922 18446
rect 5978 18390 6046 18446
rect 6102 18390 6170 18446
rect 6226 18390 6294 18446
rect 6350 18390 6418 18446
rect 6474 18390 6542 18446
rect 6598 18390 6666 18446
rect 6722 18390 6790 18446
rect 6846 18390 6914 18446
rect 6970 18390 7038 18446
rect 7094 18390 7104 18446
rect 5168 18322 7104 18390
rect 5168 18266 5178 18322
rect 5234 18266 5302 18322
rect 5358 18266 5426 18322
rect 5482 18266 5550 18322
rect 5606 18266 5674 18322
rect 5730 18266 5798 18322
rect 5854 18266 5922 18322
rect 5978 18266 6046 18322
rect 6102 18266 6170 18322
rect 6226 18266 6294 18322
rect 6350 18266 6418 18322
rect 6474 18266 6542 18322
rect 6598 18266 6666 18322
rect 6722 18266 6790 18322
rect 6846 18266 6914 18322
rect 6970 18266 7038 18322
rect 7094 18266 7104 18322
rect 5168 18198 7104 18266
rect 5168 18142 5178 18198
rect 5234 18142 5302 18198
rect 5358 18142 5426 18198
rect 5482 18142 5550 18198
rect 5606 18142 5674 18198
rect 5730 18142 5798 18198
rect 5854 18142 5922 18198
rect 5978 18142 6046 18198
rect 6102 18142 6170 18198
rect 6226 18142 6294 18198
rect 6350 18142 6418 18198
rect 6474 18142 6542 18198
rect 6598 18142 6666 18198
rect 6722 18142 6790 18198
rect 6846 18142 6914 18198
rect 6970 18142 7038 18198
rect 7094 18142 7104 18198
rect 5168 18074 7104 18142
rect 5168 18018 5178 18074
rect 5234 18018 5302 18074
rect 5358 18018 5426 18074
rect 5482 18018 5550 18074
rect 5606 18018 5674 18074
rect 5730 18018 5798 18074
rect 5854 18018 5922 18074
rect 5978 18018 6046 18074
rect 6102 18018 6170 18074
rect 6226 18018 6294 18074
rect 6350 18018 6418 18074
rect 6474 18018 6542 18074
rect 6598 18018 6666 18074
rect 6722 18018 6790 18074
rect 6846 18018 6914 18074
rect 6970 18018 7038 18074
rect 7094 18018 7104 18074
rect 5168 17950 7104 18018
rect 5168 17894 5178 17950
rect 5234 17894 5302 17950
rect 5358 17894 5426 17950
rect 5482 17894 5550 17950
rect 5606 17894 5674 17950
rect 5730 17894 5798 17950
rect 5854 17894 5922 17950
rect 5978 17894 6046 17950
rect 6102 17894 6170 17950
rect 6226 17894 6294 17950
rect 6350 17894 6418 17950
rect 6474 17894 6542 17950
rect 6598 17894 6666 17950
rect 6722 17894 6790 17950
rect 6846 17894 6914 17950
rect 6970 17894 7038 17950
rect 7094 17894 7104 17950
rect 5168 17826 7104 17894
rect 5168 17770 5178 17826
rect 5234 17770 5302 17826
rect 5358 17770 5426 17826
rect 5482 17770 5550 17826
rect 5606 17770 5674 17826
rect 5730 17770 5798 17826
rect 5854 17770 5922 17826
rect 5978 17770 6046 17826
rect 6102 17770 6170 17826
rect 6226 17770 6294 17826
rect 6350 17770 6418 17826
rect 6474 17770 6542 17826
rect 6598 17770 6666 17826
rect 6722 17770 6790 17826
rect 6846 17770 6914 17826
rect 6970 17770 7038 17826
rect 7094 17770 7104 17826
rect 5168 17702 7104 17770
rect 5168 17646 5178 17702
rect 5234 17646 5302 17702
rect 5358 17646 5426 17702
rect 5482 17646 5550 17702
rect 5606 17646 5674 17702
rect 5730 17646 5798 17702
rect 5854 17646 5922 17702
rect 5978 17646 6046 17702
rect 6102 17646 6170 17702
rect 6226 17646 6294 17702
rect 6350 17646 6418 17702
rect 6474 17646 6542 17702
rect 6598 17646 6666 17702
rect 6722 17646 6790 17702
rect 6846 17646 6914 17702
rect 6970 17646 7038 17702
rect 7094 17646 7104 17702
rect 5168 17636 7104 17646
rect 7874 20554 9810 20564
rect 7874 20498 7884 20554
rect 7940 20498 8008 20554
rect 8064 20498 8132 20554
rect 8188 20498 8256 20554
rect 8312 20498 8380 20554
rect 8436 20498 8504 20554
rect 8560 20498 8628 20554
rect 8684 20498 8752 20554
rect 8808 20498 8876 20554
rect 8932 20498 9000 20554
rect 9056 20498 9124 20554
rect 9180 20498 9248 20554
rect 9304 20498 9372 20554
rect 9428 20498 9496 20554
rect 9552 20498 9620 20554
rect 9676 20498 9744 20554
rect 9800 20498 9810 20554
rect 7874 20430 9810 20498
rect 7874 20374 7884 20430
rect 7940 20374 8008 20430
rect 8064 20374 8132 20430
rect 8188 20374 8256 20430
rect 8312 20374 8380 20430
rect 8436 20374 8504 20430
rect 8560 20374 8628 20430
rect 8684 20374 8752 20430
rect 8808 20374 8876 20430
rect 8932 20374 9000 20430
rect 9056 20374 9124 20430
rect 9180 20374 9248 20430
rect 9304 20374 9372 20430
rect 9428 20374 9496 20430
rect 9552 20374 9620 20430
rect 9676 20374 9744 20430
rect 9800 20374 9810 20430
rect 7874 20306 9810 20374
rect 7874 20250 7884 20306
rect 7940 20250 8008 20306
rect 8064 20250 8132 20306
rect 8188 20250 8256 20306
rect 8312 20250 8380 20306
rect 8436 20250 8504 20306
rect 8560 20250 8628 20306
rect 8684 20250 8752 20306
rect 8808 20250 8876 20306
rect 8932 20250 9000 20306
rect 9056 20250 9124 20306
rect 9180 20250 9248 20306
rect 9304 20250 9372 20306
rect 9428 20250 9496 20306
rect 9552 20250 9620 20306
rect 9676 20250 9744 20306
rect 9800 20250 9810 20306
rect 7874 20182 9810 20250
rect 7874 20126 7884 20182
rect 7940 20126 8008 20182
rect 8064 20126 8132 20182
rect 8188 20126 8256 20182
rect 8312 20126 8380 20182
rect 8436 20126 8504 20182
rect 8560 20126 8628 20182
rect 8684 20126 8752 20182
rect 8808 20126 8876 20182
rect 8932 20126 9000 20182
rect 9056 20126 9124 20182
rect 9180 20126 9248 20182
rect 9304 20126 9372 20182
rect 9428 20126 9496 20182
rect 9552 20126 9620 20182
rect 9676 20126 9744 20182
rect 9800 20126 9810 20182
rect 7874 20058 9810 20126
rect 7874 20002 7884 20058
rect 7940 20002 8008 20058
rect 8064 20002 8132 20058
rect 8188 20002 8256 20058
rect 8312 20002 8380 20058
rect 8436 20002 8504 20058
rect 8560 20002 8628 20058
rect 8684 20002 8752 20058
rect 8808 20002 8876 20058
rect 8932 20002 9000 20058
rect 9056 20002 9124 20058
rect 9180 20002 9248 20058
rect 9304 20002 9372 20058
rect 9428 20002 9496 20058
rect 9552 20002 9620 20058
rect 9676 20002 9744 20058
rect 9800 20002 9810 20058
rect 7874 19934 9810 20002
rect 7874 19878 7884 19934
rect 7940 19878 8008 19934
rect 8064 19878 8132 19934
rect 8188 19878 8256 19934
rect 8312 19878 8380 19934
rect 8436 19878 8504 19934
rect 8560 19878 8628 19934
rect 8684 19878 8752 19934
rect 8808 19878 8876 19934
rect 8932 19878 9000 19934
rect 9056 19878 9124 19934
rect 9180 19878 9248 19934
rect 9304 19878 9372 19934
rect 9428 19878 9496 19934
rect 9552 19878 9620 19934
rect 9676 19878 9744 19934
rect 9800 19878 9810 19934
rect 7874 19810 9810 19878
rect 7874 19754 7884 19810
rect 7940 19754 8008 19810
rect 8064 19754 8132 19810
rect 8188 19754 8256 19810
rect 8312 19754 8380 19810
rect 8436 19754 8504 19810
rect 8560 19754 8628 19810
rect 8684 19754 8752 19810
rect 8808 19754 8876 19810
rect 8932 19754 9000 19810
rect 9056 19754 9124 19810
rect 9180 19754 9248 19810
rect 9304 19754 9372 19810
rect 9428 19754 9496 19810
rect 9552 19754 9620 19810
rect 9676 19754 9744 19810
rect 9800 19754 9810 19810
rect 7874 19686 9810 19754
rect 7874 19630 7884 19686
rect 7940 19630 8008 19686
rect 8064 19630 8132 19686
rect 8188 19630 8256 19686
rect 8312 19630 8380 19686
rect 8436 19630 8504 19686
rect 8560 19630 8628 19686
rect 8684 19630 8752 19686
rect 8808 19630 8876 19686
rect 8932 19630 9000 19686
rect 9056 19630 9124 19686
rect 9180 19630 9248 19686
rect 9304 19630 9372 19686
rect 9428 19630 9496 19686
rect 9552 19630 9620 19686
rect 9676 19630 9744 19686
rect 9800 19630 9810 19686
rect 7874 19562 9810 19630
rect 7874 19506 7884 19562
rect 7940 19506 8008 19562
rect 8064 19506 8132 19562
rect 8188 19506 8256 19562
rect 8312 19506 8380 19562
rect 8436 19506 8504 19562
rect 8560 19506 8628 19562
rect 8684 19506 8752 19562
rect 8808 19506 8876 19562
rect 8932 19506 9000 19562
rect 9056 19506 9124 19562
rect 9180 19506 9248 19562
rect 9304 19506 9372 19562
rect 9428 19506 9496 19562
rect 9552 19506 9620 19562
rect 9676 19506 9744 19562
rect 9800 19506 9810 19562
rect 7874 19438 9810 19506
rect 7874 19382 7884 19438
rect 7940 19382 8008 19438
rect 8064 19382 8132 19438
rect 8188 19382 8256 19438
rect 8312 19382 8380 19438
rect 8436 19382 8504 19438
rect 8560 19382 8628 19438
rect 8684 19382 8752 19438
rect 8808 19382 8876 19438
rect 8932 19382 9000 19438
rect 9056 19382 9124 19438
rect 9180 19382 9248 19438
rect 9304 19382 9372 19438
rect 9428 19382 9496 19438
rect 9552 19382 9620 19438
rect 9676 19382 9744 19438
rect 9800 19382 9810 19438
rect 7874 19314 9810 19382
rect 7874 19258 7884 19314
rect 7940 19258 8008 19314
rect 8064 19258 8132 19314
rect 8188 19258 8256 19314
rect 8312 19258 8380 19314
rect 8436 19258 8504 19314
rect 8560 19258 8628 19314
rect 8684 19258 8752 19314
rect 8808 19258 8876 19314
rect 8932 19258 9000 19314
rect 9056 19258 9124 19314
rect 9180 19258 9248 19314
rect 9304 19258 9372 19314
rect 9428 19258 9496 19314
rect 9552 19258 9620 19314
rect 9676 19258 9744 19314
rect 9800 19258 9810 19314
rect 7874 19190 9810 19258
rect 7874 19134 7884 19190
rect 7940 19134 8008 19190
rect 8064 19134 8132 19190
rect 8188 19134 8256 19190
rect 8312 19134 8380 19190
rect 8436 19134 8504 19190
rect 8560 19134 8628 19190
rect 8684 19134 8752 19190
rect 8808 19134 8876 19190
rect 8932 19134 9000 19190
rect 9056 19134 9124 19190
rect 9180 19134 9248 19190
rect 9304 19134 9372 19190
rect 9428 19134 9496 19190
rect 9552 19134 9620 19190
rect 9676 19134 9744 19190
rect 9800 19134 9810 19190
rect 7874 19066 9810 19134
rect 7874 19010 7884 19066
rect 7940 19010 8008 19066
rect 8064 19010 8132 19066
rect 8188 19010 8256 19066
rect 8312 19010 8380 19066
rect 8436 19010 8504 19066
rect 8560 19010 8628 19066
rect 8684 19010 8752 19066
rect 8808 19010 8876 19066
rect 8932 19010 9000 19066
rect 9056 19010 9124 19066
rect 9180 19010 9248 19066
rect 9304 19010 9372 19066
rect 9428 19010 9496 19066
rect 9552 19010 9620 19066
rect 9676 19010 9744 19066
rect 9800 19010 9810 19066
rect 7874 18942 9810 19010
rect 7874 18886 7884 18942
rect 7940 18886 8008 18942
rect 8064 18886 8132 18942
rect 8188 18886 8256 18942
rect 8312 18886 8380 18942
rect 8436 18886 8504 18942
rect 8560 18886 8628 18942
rect 8684 18886 8752 18942
rect 8808 18886 8876 18942
rect 8932 18886 9000 18942
rect 9056 18886 9124 18942
rect 9180 18886 9248 18942
rect 9304 18886 9372 18942
rect 9428 18886 9496 18942
rect 9552 18886 9620 18942
rect 9676 18886 9744 18942
rect 9800 18886 9810 18942
rect 7874 18818 9810 18886
rect 7874 18762 7884 18818
rect 7940 18762 8008 18818
rect 8064 18762 8132 18818
rect 8188 18762 8256 18818
rect 8312 18762 8380 18818
rect 8436 18762 8504 18818
rect 8560 18762 8628 18818
rect 8684 18762 8752 18818
rect 8808 18762 8876 18818
rect 8932 18762 9000 18818
rect 9056 18762 9124 18818
rect 9180 18762 9248 18818
rect 9304 18762 9372 18818
rect 9428 18762 9496 18818
rect 9552 18762 9620 18818
rect 9676 18762 9744 18818
rect 9800 18762 9810 18818
rect 7874 18694 9810 18762
rect 7874 18638 7884 18694
rect 7940 18638 8008 18694
rect 8064 18638 8132 18694
rect 8188 18638 8256 18694
rect 8312 18638 8380 18694
rect 8436 18638 8504 18694
rect 8560 18638 8628 18694
rect 8684 18638 8752 18694
rect 8808 18638 8876 18694
rect 8932 18638 9000 18694
rect 9056 18638 9124 18694
rect 9180 18638 9248 18694
rect 9304 18638 9372 18694
rect 9428 18638 9496 18694
rect 9552 18638 9620 18694
rect 9676 18638 9744 18694
rect 9800 18638 9810 18694
rect 7874 18570 9810 18638
rect 7874 18514 7884 18570
rect 7940 18514 8008 18570
rect 8064 18514 8132 18570
rect 8188 18514 8256 18570
rect 8312 18514 8380 18570
rect 8436 18514 8504 18570
rect 8560 18514 8628 18570
rect 8684 18514 8752 18570
rect 8808 18514 8876 18570
rect 8932 18514 9000 18570
rect 9056 18514 9124 18570
rect 9180 18514 9248 18570
rect 9304 18514 9372 18570
rect 9428 18514 9496 18570
rect 9552 18514 9620 18570
rect 9676 18514 9744 18570
rect 9800 18514 9810 18570
rect 7874 18446 9810 18514
rect 7874 18390 7884 18446
rect 7940 18390 8008 18446
rect 8064 18390 8132 18446
rect 8188 18390 8256 18446
rect 8312 18390 8380 18446
rect 8436 18390 8504 18446
rect 8560 18390 8628 18446
rect 8684 18390 8752 18446
rect 8808 18390 8876 18446
rect 8932 18390 9000 18446
rect 9056 18390 9124 18446
rect 9180 18390 9248 18446
rect 9304 18390 9372 18446
rect 9428 18390 9496 18446
rect 9552 18390 9620 18446
rect 9676 18390 9744 18446
rect 9800 18390 9810 18446
rect 7874 18322 9810 18390
rect 7874 18266 7884 18322
rect 7940 18266 8008 18322
rect 8064 18266 8132 18322
rect 8188 18266 8256 18322
rect 8312 18266 8380 18322
rect 8436 18266 8504 18322
rect 8560 18266 8628 18322
rect 8684 18266 8752 18322
rect 8808 18266 8876 18322
rect 8932 18266 9000 18322
rect 9056 18266 9124 18322
rect 9180 18266 9248 18322
rect 9304 18266 9372 18322
rect 9428 18266 9496 18322
rect 9552 18266 9620 18322
rect 9676 18266 9744 18322
rect 9800 18266 9810 18322
rect 7874 18198 9810 18266
rect 7874 18142 7884 18198
rect 7940 18142 8008 18198
rect 8064 18142 8132 18198
rect 8188 18142 8256 18198
rect 8312 18142 8380 18198
rect 8436 18142 8504 18198
rect 8560 18142 8628 18198
rect 8684 18142 8752 18198
rect 8808 18142 8876 18198
rect 8932 18142 9000 18198
rect 9056 18142 9124 18198
rect 9180 18142 9248 18198
rect 9304 18142 9372 18198
rect 9428 18142 9496 18198
rect 9552 18142 9620 18198
rect 9676 18142 9744 18198
rect 9800 18142 9810 18198
rect 7874 18074 9810 18142
rect 7874 18018 7884 18074
rect 7940 18018 8008 18074
rect 8064 18018 8132 18074
rect 8188 18018 8256 18074
rect 8312 18018 8380 18074
rect 8436 18018 8504 18074
rect 8560 18018 8628 18074
rect 8684 18018 8752 18074
rect 8808 18018 8876 18074
rect 8932 18018 9000 18074
rect 9056 18018 9124 18074
rect 9180 18018 9248 18074
rect 9304 18018 9372 18074
rect 9428 18018 9496 18074
rect 9552 18018 9620 18074
rect 9676 18018 9744 18074
rect 9800 18018 9810 18074
rect 7874 17950 9810 18018
rect 7874 17894 7884 17950
rect 7940 17894 8008 17950
rect 8064 17894 8132 17950
rect 8188 17894 8256 17950
rect 8312 17894 8380 17950
rect 8436 17894 8504 17950
rect 8560 17894 8628 17950
rect 8684 17894 8752 17950
rect 8808 17894 8876 17950
rect 8932 17894 9000 17950
rect 9056 17894 9124 17950
rect 9180 17894 9248 17950
rect 9304 17894 9372 17950
rect 9428 17894 9496 17950
rect 9552 17894 9620 17950
rect 9676 17894 9744 17950
rect 9800 17894 9810 17950
rect 7874 17826 9810 17894
rect 7874 17770 7884 17826
rect 7940 17770 8008 17826
rect 8064 17770 8132 17826
rect 8188 17770 8256 17826
rect 8312 17770 8380 17826
rect 8436 17770 8504 17826
rect 8560 17770 8628 17826
rect 8684 17770 8752 17826
rect 8808 17770 8876 17826
rect 8932 17770 9000 17826
rect 9056 17770 9124 17826
rect 9180 17770 9248 17826
rect 9304 17770 9372 17826
rect 9428 17770 9496 17826
rect 9552 17770 9620 17826
rect 9676 17770 9744 17826
rect 9800 17770 9810 17826
rect 7874 17702 9810 17770
rect 7874 17646 7884 17702
rect 7940 17646 8008 17702
rect 8064 17646 8132 17702
rect 8188 17646 8256 17702
rect 8312 17646 8380 17702
rect 8436 17646 8504 17702
rect 8560 17646 8628 17702
rect 8684 17646 8752 17702
rect 8808 17646 8876 17702
rect 8932 17646 9000 17702
rect 9056 17646 9124 17702
rect 9180 17646 9248 17702
rect 9304 17646 9372 17702
rect 9428 17646 9496 17702
rect 9552 17646 9620 17702
rect 9676 17646 9744 17702
rect 9800 17646 9810 17702
rect 7874 17636 9810 17646
rect 10244 20554 12180 20564
rect 10244 20498 10254 20554
rect 10310 20498 10378 20554
rect 10434 20498 10502 20554
rect 10558 20498 10626 20554
rect 10682 20498 10750 20554
rect 10806 20498 10874 20554
rect 10930 20498 10998 20554
rect 11054 20498 11122 20554
rect 11178 20498 11246 20554
rect 11302 20498 11370 20554
rect 11426 20498 11494 20554
rect 11550 20498 11618 20554
rect 11674 20498 11742 20554
rect 11798 20498 11866 20554
rect 11922 20498 11990 20554
rect 12046 20498 12114 20554
rect 12170 20498 12180 20554
rect 10244 20430 12180 20498
rect 10244 20374 10254 20430
rect 10310 20374 10378 20430
rect 10434 20374 10502 20430
rect 10558 20374 10626 20430
rect 10682 20374 10750 20430
rect 10806 20374 10874 20430
rect 10930 20374 10998 20430
rect 11054 20374 11122 20430
rect 11178 20374 11246 20430
rect 11302 20374 11370 20430
rect 11426 20374 11494 20430
rect 11550 20374 11618 20430
rect 11674 20374 11742 20430
rect 11798 20374 11866 20430
rect 11922 20374 11990 20430
rect 12046 20374 12114 20430
rect 12170 20374 12180 20430
rect 10244 20306 12180 20374
rect 10244 20250 10254 20306
rect 10310 20250 10378 20306
rect 10434 20250 10502 20306
rect 10558 20250 10626 20306
rect 10682 20250 10750 20306
rect 10806 20250 10874 20306
rect 10930 20250 10998 20306
rect 11054 20250 11122 20306
rect 11178 20250 11246 20306
rect 11302 20250 11370 20306
rect 11426 20250 11494 20306
rect 11550 20250 11618 20306
rect 11674 20250 11742 20306
rect 11798 20250 11866 20306
rect 11922 20250 11990 20306
rect 12046 20250 12114 20306
rect 12170 20250 12180 20306
rect 10244 20182 12180 20250
rect 10244 20126 10254 20182
rect 10310 20126 10378 20182
rect 10434 20126 10502 20182
rect 10558 20126 10626 20182
rect 10682 20126 10750 20182
rect 10806 20126 10874 20182
rect 10930 20126 10998 20182
rect 11054 20126 11122 20182
rect 11178 20126 11246 20182
rect 11302 20126 11370 20182
rect 11426 20126 11494 20182
rect 11550 20126 11618 20182
rect 11674 20126 11742 20182
rect 11798 20126 11866 20182
rect 11922 20126 11990 20182
rect 12046 20126 12114 20182
rect 12170 20126 12180 20182
rect 10244 20058 12180 20126
rect 10244 20002 10254 20058
rect 10310 20002 10378 20058
rect 10434 20002 10502 20058
rect 10558 20002 10626 20058
rect 10682 20002 10750 20058
rect 10806 20002 10874 20058
rect 10930 20002 10998 20058
rect 11054 20002 11122 20058
rect 11178 20002 11246 20058
rect 11302 20002 11370 20058
rect 11426 20002 11494 20058
rect 11550 20002 11618 20058
rect 11674 20002 11742 20058
rect 11798 20002 11866 20058
rect 11922 20002 11990 20058
rect 12046 20002 12114 20058
rect 12170 20002 12180 20058
rect 10244 19934 12180 20002
rect 10244 19878 10254 19934
rect 10310 19878 10378 19934
rect 10434 19878 10502 19934
rect 10558 19878 10626 19934
rect 10682 19878 10750 19934
rect 10806 19878 10874 19934
rect 10930 19878 10998 19934
rect 11054 19878 11122 19934
rect 11178 19878 11246 19934
rect 11302 19878 11370 19934
rect 11426 19878 11494 19934
rect 11550 19878 11618 19934
rect 11674 19878 11742 19934
rect 11798 19878 11866 19934
rect 11922 19878 11990 19934
rect 12046 19878 12114 19934
rect 12170 19878 12180 19934
rect 10244 19810 12180 19878
rect 10244 19754 10254 19810
rect 10310 19754 10378 19810
rect 10434 19754 10502 19810
rect 10558 19754 10626 19810
rect 10682 19754 10750 19810
rect 10806 19754 10874 19810
rect 10930 19754 10998 19810
rect 11054 19754 11122 19810
rect 11178 19754 11246 19810
rect 11302 19754 11370 19810
rect 11426 19754 11494 19810
rect 11550 19754 11618 19810
rect 11674 19754 11742 19810
rect 11798 19754 11866 19810
rect 11922 19754 11990 19810
rect 12046 19754 12114 19810
rect 12170 19754 12180 19810
rect 10244 19686 12180 19754
rect 10244 19630 10254 19686
rect 10310 19630 10378 19686
rect 10434 19630 10502 19686
rect 10558 19630 10626 19686
rect 10682 19630 10750 19686
rect 10806 19630 10874 19686
rect 10930 19630 10998 19686
rect 11054 19630 11122 19686
rect 11178 19630 11246 19686
rect 11302 19630 11370 19686
rect 11426 19630 11494 19686
rect 11550 19630 11618 19686
rect 11674 19630 11742 19686
rect 11798 19630 11866 19686
rect 11922 19630 11990 19686
rect 12046 19630 12114 19686
rect 12170 19630 12180 19686
rect 10244 19562 12180 19630
rect 10244 19506 10254 19562
rect 10310 19506 10378 19562
rect 10434 19506 10502 19562
rect 10558 19506 10626 19562
rect 10682 19506 10750 19562
rect 10806 19506 10874 19562
rect 10930 19506 10998 19562
rect 11054 19506 11122 19562
rect 11178 19506 11246 19562
rect 11302 19506 11370 19562
rect 11426 19506 11494 19562
rect 11550 19506 11618 19562
rect 11674 19506 11742 19562
rect 11798 19506 11866 19562
rect 11922 19506 11990 19562
rect 12046 19506 12114 19562
rect 12170 19506 12180 19562
rect 10244 19438 12180 19506
rect 10244 19382 10254 19438
rect 10310 19382 10378 19438
rect 10434 19382 10502 19438
rect 10558 19382 10626 19438
rect 10682 19382 10750 19438
rect 10806 19382 10874 19438
rect 10930 19382 10998 19438
rect 11054 19382 11122 19438
rect 11178 19382 11246 19438
rect 11302 19382 11370 19438
rect 11426 19382 11494 19438
rect 11550 19382 11618 19438
rect 11674 19382 11742 19438
rect 11798 19382 11866 19438
rect 11922 19382 11990 19438
rect 12046 19382 12114 19438
rect 12170 19382 12180 19438
rect 10244 19314 12180 19382
rect 10244 19258 10254 19314
rect 10310 19258 10378 19314
rect 10434 19258 10502 19314
rect 10558 19258 10626 19314
rect 10682 19258 10750 19314
rect 10806 19258 10874 19314
rect 10930 19258 10998 19314
rect 11054 19258 11122 19314
rect 11178 19258 11246 19314
rect 11302 19258 11370 19314
rect 11426 19258 11494 19314
rect 11550 19258 11618 19314
rect 11674 19258 11742 19314
rect 11798 19258 11866 19314
rect 11922 19258 11990 19314
rect 12046 19258 12114 19314
rect 12170 19258 12180 19314
rect 10244 19190 12180 19258
rect 10244 19134 10254 19190
rect 10310 19134 10378 19190
rect 10434 19134 10502 19190
rect 10558 19134 10626 19190
rect 10682 19134 10750 19190
rect 10806 19134 10874 19190
rect 10930 19134 10998 19190
rect 11054 19134 11122 19190
rect 11178 19134 11246 19190
rect 11302 19134 11370 19190
rect 11426 19134 11494 19190
rect 11550 19134 11618 19190
rect 11674 19134 11742 19190
rect 11798 19134 11866 19190
rect 11922 19134 11990 19190
rect 12046 19134 12114 19190
rect 12170 19134 12180 19190
rect 10244 19066 12180 19134
rect 10244 19010 10254 19066
rect 10310 19010 10378 19066
rect 10434 19010 10502 19066
rect 10558 19010 10626 19066
rect 10682 19010 10750 19066
rect 10806 19010 10874 19066
rect 10930 19010 10998 19066
rect 11054 19010 11122 19066
rect 11178 19010 11246 19066
rect 11302 19010 11370 19066
rect 11426 19010 11494 19066
rect 11550 19010 11618 19066
rect 11674 19010 11742 19066
rect 11798 19010 11866 19066
rect 11922 19010 11990 19066
rect 12046 19010 12114 19066
rect 12170 19010 12180 19066
rect 10244 18942 12180 19010
rect 10244 18886 10254 18942
rect 10310 18886 10378 18942
rect 10434 18886 10502 18942
rect 10558 18886 10626 18942
rect 10682 18886 10750 18942
rect 10806 18886 10874 18942
rect 10930 18886 10998 18942
rect 11054 18886 11122 18942
rect 11178 18886 11246 18942
rect 11302 18886 11370 18942
rect 11426 18886 11494 18942
rect 11550 18886 11618 18942
rect 11674 18886 11742 18942
rect 11798 18886 11866 18942
rect 11922 18886 11990 18942
rect 12046 18886 12114 18942
rect 12170 18886 12180 18942
rect 10244 18818 12180 18886
rect 10244 18762 10254 18818
rect 10310 18762 10378 18818
rect 10434 18762 10502 18818
rect 10558 18762 10626 18818
rect 10682 18762 10750 18818
rect 10806 18762 10874 18818
rect 10930 18762 10998 18818
rect 11054 18762 11122 18818
rect 11178 18762 11246 18818
rect 11302 18762 11370 18818
rect 11426 18762 11494 18818
rect 11550 18762 11618 18818
rect 11674 18762 11742 18818
rect 11798 18762 11866 18818
rect 11922 18762 11990 18818
rect 12046 18762 12114 18818
rect 12170 18762 12180 18818
rect 10244 18694 12180 18762
rect 10244 18638 10254 18694
rect 10310 18638 10378 18694
rect 10434 18638 10502 18694
rect 10558 18638 10626 18694
rect 10682 18638 10750 18694
rect 10806 18638 10874 18694
rect 10930 18638 10998 18694
rect 11054 18638 11122 18694
rect 11178 18638 11246 18694
rect 11302 18638 11370 18694
rect 11426 18638 11494 18694
rect 11550 18638 11618 18694
rect 11674 18638 11742 18694
rect 11798 18638 11866 18694
rect 11922 18638 11990 18694
rect 12046 18638 12114 18694
rect 12170 18638 12180 18694
rect 10244 18570 12180 18638
rect 10244 18514 10254 18570
rect 10310 18514 10378 18570
rect 10434 18514 10502 18570
rect 10558 18514 10626 18570
rect 10682 18514 10750 18570
rect 10806 18514 10874 18570
rect 10930 18514 10998 18570
rect 11054 18514 11122 18570
rect 11178 18514 11246 18570
rect 11302 18514 11370 18570
rect 11426 18514 11494 18570
rect 11550 18514 11618 18570
rect 11674 18514 11742 18570
rect 11798 18514 11866 18570
rect 11922 18514 11990 18570
rect 12046 18514 12114 18570
rect 12170 18514 12180 18570
rect 10244 18446 12180 18514
rect 10244 18390 10254 18446
rect 10310 18390 10378 18446
rect 10434 18390 10502 18446
rect 10558 18390 10626 18446
rect 10682 18390 10750 18446
rect 10806 18390 10874 18446
rect 10930 18390 10998 18446
rect 11054 18390 11122 18446
rect 11178 18390 11246 18446
rect 11302 18390 11370 18446
rect 11426 18390 11494 18446
rect 11550 18390 11618 18446
rect 11674 18390 11742 18446
rect 11798 18390 11866 18446
rect 11922 18390 11990 18446
rect 12046 18390 12114 18446
rect 12170 18390 12180 18446
rect 10244 18322 12180 18390
rect 10244 18266 10254 18322
rect 10310 18266 10378 18322
rect 10434 18266 10502 18322
rect 10558 18266 10626 18322
rect 10682 18266 10750 18322
rect 10806 18266 10874 18322
rect 10930 18266 10998 18322
rect 11054 18266 11122 18322
rect 11178 18266 11246 18322
rect 11302 18266 11370 18322
rect 11426 18266 11494 18322
rect 11550 18266 11618 18322
rect 11674 18266 11742 18322
rect 11798 18266 11866 18322
rect 11922 18266 11990 18322
rect 12046 18266 12114 18322
rect 12170 18266 12180 18322
rect 10244 18198 12180 18266
rect 10244 18142 10254 18198
rect 10310 18142 10378 18198
rect 10434 18142 10502 18198
rect 10558 18142 10626 18198
rect 10682 18142 10750 18198
rect 10806 18142 10874 18198
rect 10930 18142 10998 18198
rect 11054 18142 11122 18198
rect 11178 18142 11246 18198
rect 11302 18142 11370 18198
rect 11426 18142 11494 18198
rect 11550 18142 11618 18198
rect 11674 18142 11742 18198
rect 11798 18142 11866 18198
rect 11922 18142 11990 18198
rect 12046 18142 12114 18198
rect 12170 18142 12180 18198
rect 10244 18074 12180 18142
rect 10244 18018 10254 18074
rect 10310 18018 10378 18074
rect 10434 18018 10502 18074
rect 10558 18018 10626 18074
rect 10682 18018 10750 18074
rect 10806 18018 10874 18074
rect 10930 18018 10998 18074
rect 11054 18018 11122 18074
rect 11178 18018 11246 18074
rect 11302 18018 11370 18074
rect 11426 18018 11494 18074
rect 11550 18018 11618 18074
rect 11674 18018 11742 18074
rect 11798 18018 11866 18074
rect 11922 18018 11990 18074
rect 12046 18018 12114 18074
rect 12170 18018 12180 18074
rect 10244 17950 12180 18018
rect 10244 17894 10254 17950
rect 10310 17894 10378 17950
rect 10434 17894 10502 17950
rect 10558 17894 10626 17950
rect 10682 17894 10750 17950
rect 10806 17894 10874 17950
rect 10930 17894 10998 17950
rect 11054 17894 11122 17950
rect 11178 17894 11246 17950
rect 11302 17894 11370 17950
rect 11426 17894 11494 17950
rect 11550 17894 11618 17950
rect 11674 17894 11742 17950
rect 11798 17894 11866 17950
rect 11922 17894 11990 17950
rect 12046 17894 12114 17950
rect 12170 17894 12180 17950
rect 10244 17826 12180 17894
rect 10244 17770 10254 17826
rect 10310 17770 10378 17826
rect 10434 17770 10502 17826
rect 10558 17770 10626 17826
rect 10682 17770 10750 17826
rect 10806 17770 10874 17826
rect 10930 17770 10998 17826
rect 11054 17770 11122 17826
rect 11178 17770 11246 17826
rect 11302 17770 11370 17826
rect 11426 17770 11494 17826
rect 11550 17770 11618 17826
rect 11674 17770 11742 17826
rect 11798 17770 11866 17826
rect 11922 17770 11990 17826
rect 12046 17770 12114 17826
rect 12170 17770 12180 17826
rect 10244 17702 12180 17770
rect 10244 17646 10254 17702
rect 10310 17646 10378 17702
rect 10434 17646 10502 17702
rect 10558 17646 10626 17702
rect 10682 17646 10750 17702
rect 10806 17646 10874 17702
rect 10930 17646 10998 17702
rect 11054 17646 11122 17702
rect 11178 17646 11246 17702
rect 11302 17646 11370 17702
rect 11426 17646 11494 17702
rect 11550 17646 11618 17702
rect 11674 17646 11742 17702
rect 11798 17646 11866 17702
rect 11922 17646 11990 17702
rect 12046 17646 12114 17702
rect 12170 17646 12180 17702
rect 10244 17636 12180 17646
rect 12861 20554 14673 20564
rect 12861 20498 12871 20554
rect 12927 20498 12995 20554
rect 13051 20498 13119 20554
rect 13175 20498 13243 20554
rect 13299 20498 13367 20554
rect 13423 20498 13491 20554
rect 13547 20498 13615 20554
rect 13671 20498 13739 20554
rect 13795 20498 13863 20554
rect 13919 20498 13987 20554
rect 14043 20498 14111 20554
rect 14167 20498 14235 20554
rect 14291 20498 14359 20554
rect 14415 20498 14483 20554
rect 14539 20498 14607 20554
rect 14663 20498 14673 20554
rect 12861 20430 14673 20498
rect 12861 20374 12871 20430
rect 12927 20374 12995 20430
rect 13051 20374 13119 20430
rect 13175 20374 13243 20430
rect 13299 20374 13367 20430
rect 13423 20374 13491 20430
rect 13547 20374 13615 20430
rect 13671 20374 13739 20430
rect 13795 20374 13863 20430
rect 13919 20374 13987 20430
rect 14043 20374 14111 20430
rect 14167 20374 14235 20430
rect 14291 20374 14359 20430
rect 14415 20374 14483 20430
rect 14539 20374 14607 20430
rect 14663 20374 14673 20430
rect 12861 20306 14673 20374
rect 12861 20250 12871 20306
rect 12927 20250 12995 20306
rect 13051 20250 13119 20306
rect 13175 20250 13243 20306
rect 13299 20250 13367 20306
rect 13423 20250 13491 20306
rect 13547 20250 13615 20306
rect 13671 20250 13739 20306
rect 13795 20250 13863 20306
rect 13919 20250 13987 20306
rect 14043 20250 14111 20306
rect 14167 20250 14235 20306
rect 14291 20250 14359 20306
rect 14415 20250 14483 20306
rect 14539 20250 14607 20306
rect 14663 20250 14673 20306
rect 12861 20182 14673 20250
rect 12861 20126 12871 20182
rect 12927 20126 12995 20182
rect 13051 20126 13119 20182
rect 13175 20126 13243 20182
rect 13299 20126 13367 20182
rect 13423 20126 13491 20182
rect 13547 20126 13615 20182
rect 13671 20126 13739 20182
rect 13795 20126 13863 20182
rect 13919 20126 13987 20182
rect 14043 20126 14111 20182
rect 14167 20126 14235 20182
rect 14291 20126 14359 20182
rect 14415 20126 14483 20182
rect 14539 20126 14607 20182
rect 14663 20126 14673 20182
rect 12861 20058 14673 20126
rect 12861 20002 12871 20058
rect 12927 20002 12995 20058
rect 13051 20002 13119 20058
rect 13175 20002 13243 20058
rect 13299 20002 13367 20058
rect 13423 20002 13491 20058
rect 13547 20002 13615 20058
rect 13671 20002 13739 20058
rect 13795 20002 13863 20058
rect 13919 20002 13987 20058
rect 14043 20002 14111 20058
rect 14167 20002 14235 20058
rect 14291 20002 14359 20058
rect 14415 20002 14483 20058
rect 14539 20002 14607 20058
rect 14663 20002 14673 20058
rect 12861 19934 14673 20002
rect 12861 19878 12871 19934
rect 12927 19878 12995 19934
rect 13051 19878 13119 19934
rect 13175 19878 13243 19934
rect 13299 19878 13367 19934
rect 13423 19878 13491 19934
rect 13547 19878 13615 19934
rect 13671 19878 13739 19934
rect 13795 19878 13863 19934
rect 13919 19878 13987 19934
rect 14043 19878 14111 19934
rect 14167 19878 14235 19934
rect 14291 19878 14359 19934
rect 14415 19878 14483 19934
rect 14539 19878 14607 19934
rect 14663 19878 14673 19934
rect 12861 19810 14673 19878
rect 12861 19754 12871 19810
rect 12927 19754 12995 19810
rect 13051 19754 13119 19810
rect 13175 19754 13243 19810
rect 13299 19754 13367 19810
rect 13423 19754 13491 19810
rect 13547 19754 13615 19810
rect 13671 19754 13739 19810
rect 13795 19754 13863 19810
rect 13919 19754 13987 19810
rect 14043 19754 14111 19810
rect 14167 19754 14235 19810
rect 14291 19754 14359 19810
rect 14415 19754 14483 19810
rect 14539 19754 14607 19810
rect 14663 19754 14673 19810
rect 12861 19686 14673 19754
rect 12861 19630 12871 19686
rect 12927 19630 12995 19686
rect 13051 19630 13119 19686
rect 13175 19630 13243 19686
rect 13299 19630 13367 19686
rect 13423 19630 13491 19686
rect 13547 19630 13615 19686
rect 13671 19630 13739 19686
rect 13795 19630 13863 19686
rect 13919 19630 13987 19686
rect 14043 19630 14111 19686
rect 14167 19630 14235 19686
rect 14291 19630 14359 19686
rect 14415 19630 14483 19686
rect 14539 19630 14607 19686
rect 14663 19630 14673 19686
rect 12861 19562 14673 19630
rect 12861 19506 12871 19562
rect 12927 19506 12995 19562
rect 13051 19506 13119 19562
rect 13175 19506 13243 19562
rect 13299 19506 13367 19562
rect 13423 19506 13491 19562
rect 13547 19506 13615 19562
rect 13671 19506 13739 19562
rect 13795 19506 13863 19562
rect 13919 19506 13987 19562
rect 14043 19506 14111 19562
rect 14167 19506 14235 19562
rect 14291 19506 14359 19562
rect 14415 19506 14483 19562
rect 14539 19506 14607 19562
rect 14663 19506 14673 19562
rect 12861 19438 14673 19506
rect 12861 19382 12871 19438
rect 12927 19382 12995 19438
rect 13051 19382 13119 19438
rect 13175 19382 13243 19438
rect 13299 19382 13367 19438
rect 13423 19382 13491 19438
rect 13547 19382 13615 19438
rect 13671 19382 13739 19438
rect 13795 19382 13863 19438
rect 13919 19382 13987 19438
rect 14043 19382 14111 19438
rect 14167 19382 14235 19438
rect 14291 19382 14359 19438
rect 14415 19382 14483 19438
rect 14539 19382 14607 19438
rect 14663 19382 14673 19438
rect 12861 19314 14673 19382
rect 12861 19258 12871 19314
rect 12927 19258 12995 19314
rect 13051 19258 13119 19314
rect 13175 19258 13243 19314
rect 13299 19258 13367 19314
rect 13423 19258 13491 19314
rect 13547 19258 13615 19314
rect 13671 19258 13739 19314
rect 13795 19258 13863 19314
rect 13919 19258 13987 19314
rect 14043 19258 14111 19314
rect 14167 19258 14235 19314
rect 14291 19258 14359 19314
rect 14415 19258 14483 19314
rect 14539 19258 14607 19314
rect 14663 19258 14673 19314
rect 12861 19190 14673 19258
rect 12861 19134 12871 19190
rect 12927 19134 12995 19190
rect 13051 19134 13119 19190
rect 13175 19134 13243 19190
rect 13299 19134 13367 19190
rect 13423 19134 13491 19190
rect 13547 19134 13615 19190
rect 13671 19134 13739 19190
rect 13795 19134 13863 19190
rect 13919 19134 13987 19190
rect 14043 19134 14111 19190
rect 14167 19134 14235 19190
rect 14291 19134 14359 19190
rect 14415 19134 14483 19190
rect 14539 19134 14607 19190
rect 14663 19134 14673 19190
rect 12861 19066 14673 19134
rect 12861 19010 12871 19066
rect 12927 19010 12995 19066
rect 13051 19010 13119 19066
rect 13175 19010 13243 19066
rect 13299 19010 13367 19066
rect 13423 19010 13491 19066
rect 13547 19010 13615 19066
rect 13671 19010 13739 19066
rect 13795 19010 13863 19066
rect 13919 19010 13987 19066
rect 14043 19010 14111 19066
rect 14167 19010 14235 19066
rect 14291 19010 14359 19066
rect 14415 19010 14483 19066
rect 14539 19010 14607 19066
rect 14663 19010 14673 19066
rect 12861 18942 14673 19010
rect 12861 18886 12871 18942
rect 12927 18886 12995 18942
rect 13051 18886 13119 18942
rect 13175 18886 13243 18942
rect 13299 18886 13367 18942
rect 13423 18886 13491 18942
rect 13547 18886 13615 18942
rect 13671 18886 13739 18942
rect 13795 18886 13863 18942
rect 13919 18886 13987 18942
rect 14043 18886 14111 18942
rect 14167 18886 14235 18942
rect 14291 18886 14359 18942
rect 14415 18886 14483 18942
rect 14539 18886 14607 18942
rect 14663 18886 14673 18942
rect 12861 18818 14673 18886
rect 12861 18762 12871 18818
rect 12927 18762 12995 18818
rect 13051 18762 13119 18818
rect 13175 18762 13243 18818
rect 13299 18762 13367 18818
rect 13423 18762 13491 18818
rect 13547 18762 13615 18818
rect 13671 18762 13739 18818
rect 13795 18762 13863 18818
rect 13919 18762 13987 18818
rect 14043 18762 14111 18818
rect 14167 18762 14235 18818
rect 14291 18762 14359 18818
rect 14415 18762 14483 18818
rect 14539 18762 14607 18818
rect 14663 18762 14673 18818
rect 12861 18694 14673 18762
rect 12861 18638 12871 18694
rect 12927 18638 12995 18694
rect 13051 18638 13119 18694
rect 13175 18638 13243 18694
rect 13299 18638 13367 18694
rect 13423 18638 13491 18694
rect 13547 18638 13615 18694
rect 13671 18638 13739 18694
rect 13795 18638 13863 18694
rect 13919 18638 13987 18694
rect 14043 18638 14111 18694
rect 14167 18638 14235 18694
rect 14291 18638 14359 18694
rect 14415 18638 14483 18694
rect 14539 18638 14607 18694
rect 14663 18638 14673 18694
rect 12861 18570 14673 18638
rect 12861 18514 12871 18570
rect 12927 18514 12995 18570
rect 13051 18514 13119 18570
rect 13175 18514 13243 18570
rect 13299 18514 13367 18570
rect 13423 18514 13491 18570
rect 13547 18514 13615 18570
rect 13671 18514 13739 18570
rect 13795 18514 13863 18570
rect 13919 18514 13987 18570
rect 14043 18514 14111 18570
rect 14167 18514 14235 18570
rect 14291 18514 14359 18570
rect 14415 18514 14483 18570
rect 14539 18514 14607 18570
rect 14663 18514 14673 18570
rect 12861 18446 14673 18514
rect 12861 18390 12871 18446
rect 12927 18390 12995 18446
rect 13051 18390 13119 18446
rect 13175 18390 13243 18446
rect 13299 18390 13367 18446
rect 13423 18390 13491 18446
rect 13547 18390 13615 18446
rect 13671 18390 13739 18446
rect 13795 18390 13863 18446
rect 13919 18390 13987 18446
rect 14043 18390 14111 18446
rect 14167 18390 14235 18446
rect 14291 18390 14359 18446
rect 14415 18390 14483 18446
rect 14539 18390 14607 18446
rect 14663 18390 14673 18446
rect 12861 18322 14673 18390
rect 12861 18266 12871 18322
rect 12927 18266 12995 18322
rect 13051 18266 13119 18322
rect 13175 18266 13243 18322
rect 13299 18266 13367 18322
rect 13423 18266 13491 18322
rect 13547 18266 13615 18322
rect 13671 18266 13739 18322
rect 13795 18266 13863 18322
rect 13919 18266 13987 18322
rect 14043 18266 14111 18322
rect 14167 18266 14235 18322
rect 14291 18266 14359 18322
rect 14415 18266 14483 18322
rect 14539 18266 14607 18322
rect 14663 18266 14673 18322
rect 12861 18198 14673 18266
rect 12861 18142 12871 18198
rect 12927 18142 12995 18198
rect 13051 18142 13119 18198
rect 13175 18142 13243 18198
rect 13299 18142 13367 18198
rect 13423 18142 13491 18198
rect 13547 18142 13615 18198
rect 13671 18142 13739 18198
rect 13795 18142 13863 18198
rect 13919 18142 13987 18198
rect 14043 18142 14111 18198
rect 14167 18142 14235 18198
rect 14291 18142 14359 18198
rect 14415 18142 14483 18198
rect 14539 18142 14607 18198
rect 14663 18142 14673 18198
rect 12861 18074 14673 18142
rect 12861 18018 12871 18074
rect 12927 18018 12995 18074
rect 13051 18018 13119 18074
rect 13175 18018 13243 18074
rect 13299 18018 13367 18074
rect 13423 18018 13491 18074
rect 13547 18018 13615 18074
rect 13671 18018 13739 18074
rect 13795 18018 13863 18074
rect 13919 18018 13987 18074
rect 14043 18018 14111 18074
rect 14167 18018 14235 18074
rect 14291 18018 14359 18074
rect 14415 18018 14483 18074
rect 14539 18018 14607 18074
rect 14663 18018 14673 18074
rect 12861 17950 14673 18018
rect 12861 17894 12871 17950
rect 12927 17894 12995 17950
rect 13051 17894 13119 17950
rect 13175 17894 13243 17950
rect 13299 17894 13367 17950
rect 13423 17894 13491 17950
rect 13547 17894 13615 17950
rect 13671 17894 13739 17950
rect 13795 17894 13863 17950
rect 13919 17894 13987 17950
rect 14043 17894 14111 17950
rect 14167 17894 14235 17950
rect 14291 17894 14359 17950
rect 14415 17894 14483 17950
rect 14539 17894 14607 17950
rect 14663 17894 14673 17950
rect 12861 17826 14673 17894
rect 12861 17770 12871 17826
rect 12927 17770 12995 17826
rect 13051 17770 13119 17826
rect 13175 17770 13243 17826
rect 13299 17770 13367 17826
rect 13423 17770 13491 17826
rect 13547 17770 13615 17826
rect 13671 17770 13739 17826
rect 13795 17770 13863 17826
rect 13919 17770 13987 17826
rect 14043 17770 14111 17826
rect 14167 17770 14235 17826
rect 14291 17770 14359 17826
rect 14415 17770 14483 17826
rect 14539 17770 14607 17826
rect 14663 17770 14673 17826
rect 12861 17702 14673 17770
rect 12861 17646 12871 17702
rect 12927 17646 12995 17702
rect 13051 17646 13119 17702
rect 13175 17646 13243 17702
rect 13299 17646 13367 17702
rect 13423 17646 13491 17702
rect 13547 17646 13615 17702
rect 13671 17646 13739 17702
rect 13795 17646 13863 17702
rect 13919 17646 13987 17702
rect 14043 17646 14111 17702
rect 14167 17646 14235 17702
rect 14291 17646 14359 17702
rect 14415 17646 14483 17702
rect 14539 17646 14607 17702
rect 14663 17646 14673 17702
rect 12861 17636 14673 17646
rect 305 17354 2117 17364
rect 305 17298 315 17354
rect 371 17298 439 17354
rect 495 17298 563 17354
rect 619 17298 687 17354
rect 743 17298 811 17354
rect 867 17298 935 17354
rect 991 17298 1059 17354
rect 1115 17298 1183 17354
rect 1239 17298 1307 17354
rect 1363 17298 1431 17354
rect 1487 17298 1555 17354
rect 1611 17298 1679 17354
rect 1735 17298 1803 17354
rect 1859 17298 1927 17354
rect 1983 17298 2051 17354
rect 2107 17298 2117 17354
rect 305 17230 2117 17298
rect 305 17174 315 17230
rect 371 17174 439 17230
rect 495 17174 563 17230
rect 619 17174 687 17230
rect 743 17174 811 17230
rect 867 17174 935 17230
rect 991 17174 1059 17230
rect 1115 17174 1183 17230
rect 1239 17174 1307 17230
rect 1363 17174 1431 17230
rect 1487 17174 1555 17230
rect 1611 17174 1679 17230
rect 1735 17174 1803 17230
rect 1859 17174 1927 17230
rect 1983 17174 2051 17230
rect 2107 17174 2117 17230
rect 305 17106 2117 17174
rect 305 17050 315 17106
rect 371 17050 439 17106
rect 495 17050 563 17106
rect 619 17050 687 17106
rect 743 17050 811 17106
rect 867 17050 935 17106
rect 991 17050 1059 17106
rect 1115 17050 1183 17106
rect 1239 17050 1307 17106
rect 1363 17050 1431 17106
rect 1487 17050 1555 17106
rect 1611 17050 1679 17106
rect 1735 17050 1803 17106
rect 1859 17050 1927 17106
rect 1983 17050 2051 17106
rect 2107 17050 2117 17106
rect 305 16982 2117 17050
rect 305 16926 315 16982
rect 371 16926 439 16982
rect 495 16926 563 16982
rect 619 16926 687 16982
rect 743 16926 811 16982
rect 867 16926 935 16982
rect 991 16926 1059 16982
rect 1115 16926 1183 16982
rect 1239 16926 1307 16982
rect 1363 16926 1431 16982
rect 1487 16926 1555 16982
rect 1611 16926 1679 16982
rect 1735 16926 1803 16982
rect 1859 16926 1927 16982
rect 1983 16926 2051 16982
rect 2107 16926 2117 16982
rect 305 16858 2117 16926
rect 305 16802 315 16858
rect 371 16802 439 16858
rect 495 16802 563 16858
rect 619 16802 687 16858
rect 743 16802 811 16858
rect 867 16802 935 16858
rect 991 16802 1059 16858
rect 1115 16802 1183 16858
rect 1239 16802 1307 16858
rect 1363 16802 1431 16858
rect 1487 16802 1555 16858
rect 1611 16802 1679 16858
rect 1735 16802 1803 16858
rect 1859 16802 1927 16858
rect 1983 16802 2051 16858
rect 2107 16802 2117 16858
rect 305 16734 2117 16802
rect 305 16678 315 16734
rect 371 16678 439 16734
rect 495 16678 563 16734
rect 619 16678 687 16734
rect 743 16678 811 16734
rect 867 16678 935 16734
rect 991 16678 1059 16734
rect 1115 16678 1183 16734
rect 1239 16678 1307 16734
rect 1363 16678 1431 16734
rect 1487 16678 1555 16734
rect 1611 16678 1679 16734
rect 1735 16678 1803 16734
rect 1859 16678 1927 16734
rect 1983 16678 2051 16734
rect 2107 16678 2117 16734
rect 305 16610 2117 16678
rect 305 16554 315 16610
rect 371 16554 439 16610
rect 495 16554 563 16610
rect 619 16554 687 16610
rect 743 16554 811 16610
rect 867 16554 935 16610
rect 991 16554 1059 16610
rect 1115 16554 1183 16610
rect 1239 16554 1307 16610
rect 1363 16554 1431 16610
rect 1487 16554 1555 16610
rect 1611 16554 1679 16610
rect 1735 16554 1803 16610
rect 1859 16554 1927 16610
rect 1983 16554 2051 16610
rect 2107 16554 2117 16610
rect 305 16486 2117 16554
rect 305 16430 315 16486
rect 371 16430 439 16486
rect 495 16430 563 16486
rect 619 16430 687 16486
rect 743 16430 811 16486
rect 867 16430 935 16486
rect 991 16430 1059 16486
rect 1115 16430 1183 16486
rect 1239 16430 1307 16486
rect 1363 16430 1431 16486
rect 1487 16430 1555 16486
rect 1611 16430 1679 16486
rect 1735 16430 1803 16486
rect 1859 16430 1927 16486
rect 1983 16430 2051 16486
rect 2107 16430 2117 16486
rect 305 16362 2117 16430
rect 305 16306 315 16362
rect 371 16306 439 16362
rect 495 16306 563 16362
rect 619 16306 687 16362
rect 743 16306 811 16362
rect 867 16306 935 16362
rect 991 16306 1059 16362
rect 1115 16306 1183 16362
rect 1239 16306 1307 16362
rect 1363 16306 1431 16362
rect 1487 16306 1555 16362
rect 1611 16306 1679 16362
rect 1735 16306 1803 16362
rect 1859 16306 1927 16362
rect 1983 16306 2051 16362
rect 2107 16306 2117 16362
rect 305 16238 2117 16306
rect 305 16182 315 16238
rect 371 16182 439 16238
rect 495 16182 563 16238
rect 619 16182 687 16238
rect 743 16182 811 16238
rect 867 16182 935 16238
rect 991 16182 1059 16238
rect 1115 16182 1183 16238
rect 1239 16182 1307 16238
rect 1363 16182 1431 16238
rect 1487 16182 1555 16238
rect 1611 16182 1679 16238
rect 1735 16182 1803 16238
rect 1859 16182 1927 16238
rect 1983 16182 2051 16238
rect 2107 16182 2117 16238
rect 305 16114 2117 16182
rect 305 16058 315 16114
rect 371 16058 439 16114
rect 495 16058 563 16114
rect 619 16058 687 16114
rect 743 16058 811 16114
rect 867 16058 935 16114
rect 991 16058 1059 16114
rect 1115 16058 1183 16114
rect 1239 16058 1307 16114
rect 1363 16058 1431 16114
rect 1487 16058 1555 16114
rect 1611 16058 1679 16114
rect 1735 16058 1803 16114
rect 1859 16058 1927 16114
rect 1983 16058 2051 16114
rect 2107 16058 2117 16114
rect 305 15990 2117 16058
rect 305 15934 315 15990
rect 371 15934 439 15990
rect 495 15934 563 15990
rect 619 15934 687 15990
rect 743 15934 811 15990
rect 867 15934 935 15990
rect 991 15934 1059 15990
rect 1115 15934 1183 15990
rect 1239 15934 1307 15990
rect 1363 15934 1431 15990
rect 1487 15934 1555 15990
rect 1611 15934 1679 15990
rect 1735 15934 1803 15990
rect 1859 15934 1927 15990
rect 1983 15934 2051 15990
rect 2107 15934 2117 15990
rect 305 15866 2117 15934
rect 305 15810 315 15866
rect 371 15810 439 15866
rect 495 15810 563 15866
rect 619 15810 687 15866
rect 743 15810 811 15866
rect 867 15810 935 15866
rect 991 15810 1059 15866
rect 1115 15810 1183 15866
rect 1239 15810 1307 15866
rect 1363 15810 1431 15866
rect 1487 15810 1555 15866
rect 1611 15810 1679 15866
rect 1735 15810 1803 15866
rect 1859 15810 1927 15866
rect 1983 15810 2051 15866
rect 2107 15810 2117 15866
rect 305 15742 2117 15810
rect 305 15686 315 15742
rect 371 15686 439 15742
rect 495 15686 563 15742
rect 619 15686 687 15742
rect 743 15686 811 15742
rect 867 15686 935 15742
rect 991 15686 1059 15742
rect 1115 15686 1183 15742
rect 1239 15686 1307 15742
rect 1363 15686 1431 15742
rect 1487 15686 1555 15742
rect 1611 15686 1679 15742
rect 1735 15686 1803 15742
rect 1859 15686 1927 15742
rect 1983 15686 2051 15742
rect 2107 15686 2117 15742
rect 305 15618 2117 15686
rect 305 15562 315 15618
rect 371 15562 439 15618
rect 495 15562 563 15618
rect 619 15562 687 15618
rect 743 15562 811 15618
rect 867 15562 935 15618
rect 991 15562 1059 15618
rect 1115 15562 1183 15618
rect 1239 15562 1307 15618
rect 1363 15562 1431 15618
rect 1487 15562 1555 15618
rect 1611 15562 1679 15618
rect 1735 15562 1803 15618
rect 1859 15562 1927 15618
rect 1983 15562 2051 15618
rect 2107 15562 2117 15618
rect 305 15494 2117 15562
rect 305 15438 315 15494
rect 371 15438 439 15494
rect 495 15438 563 15494
rect 619 15438 687 15494
rect 743 15438 811 15494
rect 867 15438 935 15494
rect 991 15438 1059 15494
rect 1115 15438 1183 15494
rect 1239 15438 1307 15494
rect 1363 15438 1431 15494
rect 1487 15438 1555 15494
rect 1611 15438 1679 15494
rect 1735 15438 1803 15494
rect 1859 15438 1927 15494
rect 1983 15438 2051 15494
rect 2107 15438 2117 15494
rect 305 15370 2117 15438
rect 305 15314 315 15370
rect 371 15314 439 15370
rect 495 15314 563 15370
rect 619 15314 687 15370
rect 743 15314 811 15370
rect 867 15314 935 15370
rect 991 15314 1059 15370
rect 1115 15314 1183 15370
rect 1239 15314 1307 15370
rect 1363 15314 1431 15370
rect 1487 15314 1555 15370
rect 1611 15314 1679 15370
rect 1735 15314 1803 15370
rect 1859 15314 1927 15370
rect 1983 15314 2051 15370
rect 2107 15314 2117 15370
rect 305 15246 2117 15314
rect 305 15190 315 15246
rect 371 15190 439 15246
rect 495 15190 563 15246
rect 619 15190 687 15246
rect 743 15190 811 15246
rect 867 15190 935 15246
rect 991 15190 1059 15246
rect 1115 15190 1183 15246
rect 1239 15190 1307 15246
rect 1363 15190 1431 15246
rect 1487 15190 1555 15246
rect 1611 15190 1679 15246
rect 1735 15190 1803 15246
rect 1859 15190 1927 15246
rect 1983 15190 2051 15246
rect 2107 15190 2117 15246
rect 305 15122 2117 15190
rect 305 15066 315 15122
rect 371 15066 439 15122
rect 495 15066 563 15122
rect 619 15066 687 15122
rect 743 15066 811 15122
rect 867 15066 935 15122
rect 991 15066 1059 15122
rect 1115 15066 1183 15122
rect 1239 15066 1307 15122
rect 1363 15066 1431 15122
rect 1487 15066 1555 15122
rect 1611 15066 1679 15122
rect 1735 15066 1803 15122
rect 1859 15066 1927 15122
rect 1983 15066 2051 15122
rect 2107 15066 2117 15122
rect 305 14998 2117 15066
rect 305 14942 315 14998
rect 371 14942 439 14998
rect 495 14942 563 14998
rect 619 14942 687 14998
rect 743 14942 811 14998
rect 867 14942 935 14998
rect 991 14942 1059 14998
rect 1115 14942 1183 14998
rect 1239 14942 1307 14998
rect 1363 14942 1431 14998
rect 1487 14942 1555 14998
rect 1611 14942 1679 14998
rect 1735 14942 1803 14998
rect 1859 14942 1927 14998
rect 1983 14942 2051 14998
rect 2107 14942 2117 14998
rect 305 14874 2117 14942
rect 305 14818 315 14874
rect 371 14818 439 14874
rect 495 14818 563 14874
rect 619 14818 687 14874
rect 743 14818 811 14874
rect 867 14818 935 14874
rect 991 14818 1059 14874
rect 1115 14818 1183 14874
rect 1239 14818 1307 14874
rect 1363 14818 1431 14874
rect 1487 14818 1555 14874
rect 1611 14818 1679 14874
rect 1735 14818 1803 14874
rect 1859 14818 1927 14874
rect 1983 14818 2051 14874
rect 2107 14818 2117 14874
rect 305 14750 2117 14818
rect 305 14694 315 14750
rect 371 14694 439 14750
rect 495 14694 563 14750
rect 619 14694 687 14750
rect 743 14694 811 14750
rect 867 14694 935 14750
rect 991 14694 1059 14750
rect 1115 14694 1183 14750
rect 1239 14694 1307 14750
rect 1363 14694 1431 14750
rect 1487 14694 1555 14750
rect 1611 14694 1679 14750
rect 1735 14694 1803 14750
rect 1859 14694 1927 14750
rect 1983 14694 2051 14750
rect 2107 14694 2117 14750
rect 305 14626 2117 14694
rect 305 14570 315 14626
rect 371 14570 439 14626
rect 495 14570 563 14626
rect 619 14570 687 14626
rect 743 14570 811 14626
rect 867 14570 935 14626
rect 991 14570 1059 14626
rect 1115 14570 1183 14626
rect 1239 14570 1307 14626
rect 1363 14570 1431 14626
rect 1487 14570 1555 14626
rect 1611 14570 1679 14626
rect 1735 14570 1803 14626
rect 1859 14570 1927 14626
rect 1983 14570 2051 14626
rect 2107 14570 2117 14626
rect 305 14502 2117 14570
rect 305 14446 315 14502
rect 371 14446 439 14502
rect 495 14446 563 14502
rect 619 14446 687 14502
rect 743 14446 811 14502
rect 867 14446 935 14502
rect 991 14446 1059 14502
rect 1115 14446 1183 14502
rect 1239 14446 1307 14502
rect 1363 14446 1431 14502
rect 1487 14446 1555 14502
rect 1611 14446 1679 14502
rect 1735 14446 1803 14502
rect 1859 14446 1927 14502
rect 1983 14446 2051 14502
rect 2107 14446 2117 14502
rect 305 14436 2117 14446
rect 2798 17354 4734 17364
rect 2798 17298 2808 17354
rect 2864 17298 2932 17354
rect 2988 17298 3056 17354
rect 3112 17298 3180 17354
rect 3236 17298 3304 17354
rect 3360 17298 3428 17354
rect 3484 17298 3552 17354
rect 3608 17298 3676 17354
rect 3732 17298 3800 17354
rect 3856 17298 3924 17354
rect 3980 17298 4048 17354
rect 4104 17298 4172 17354
rect 4228 17298 4296 17354
rect 4352 17298 4420 17354
rect 4476 17298 4544 17354
rect 4600 17298 4668 17354
rect 4724 17298 4734 17354
rect 2798 17230 4734 17298
rect 2798 17174 2808 17230
rect 2864 17174 2932 17230
rect 2988 17174 3056 17230
rect 3112 17174 3180 17230
rect 3236 17174 3304 17230
rect 3360 17174 3428 17230
rect 3484 17174 3552 17230
rect 3608 17174 3676 17230
rect 3732 17174 3800 17230
rect 3856 17174 3924 17230
rect 3980 17174 4048 17230
rect 4104 17174 4172 17230
rect 4228 17174 4296 17230
rect 4352 17174 4420 17230
rect 4476 17174 4544 17230
rect 4600 17174 4668 17230
rect 4724 17174 4734 17230
rect 2798 17106 4734 17174
rect 2798 17050 2808 17106
rect 2864 17050 2932 17106
rect 2988 17050 3056 17106
rect 3112 17050 3180 17106
rect 3236 17050 3304 17106
rect 3360 17050 3428 17106
rect 3484 17050 3552 17106
rect 3608 17050 3676 17106
rect 3732 17050 3800 17106
rect 3856 17050 3924 17106
rect 3980 17050 4048 17106
rect 4104 17050 4172 17106
rect 4228 17050 4296 17106
rect 4352 17050 4420 17106
rect 4476 17050 4544 17106
rect 4600 17050 4668 17106
rect 4724 17050 4734 17106
rect 2798 16982 4734 17050
rect 2798 16926 2808 16982
rect 2864 16926 2932 16982
rect 2988 16926 3056 16982
rect 3112 16926 3180 16982
rect 3236 16926 3304 16982
rect 3360 16926 3428 16982
rect 3484 16926 3552 16982
rect 3608 16926 3676 16982
rect 3732 16926 3800 16982
rect 3856 16926 3924 16982
rect 3980 16926 4048 16982
rect 4104 16926 4172 16982
rect 4228 16926 4296 16982
rect 4352 16926 4420 16982
rect 4476 16926 4544 16982
rect 4600 16926 4668 16982
rect 4724 16926 4734 16982
rect 2798 16858 4734 16926
rect 2798 16802 2808 16858
rect 2864 16802 2932 16858
rect 2988 16802 3056 16858
rect 3112 16802 3180 16858
rect 3236 16802 3304 16858
rect 3360 16802 3428 16858
rect 3484 16802 3552 16858
rect 3608 16802 3676 16858
rect 3732 16802 3800 16858
rect 3856 16802 3924 16858
rect 3980 16802 4048 16858
rect 4104 16802 4172 16858
rect 4228 16802 4296 16858
rect 4352 16802 4420 16858
rect 4476 16802 4544 16858
rect 4600 16802 4668 16858
rect 4724 16802 4734 16858
rect 2798 16734 4734 16802
rect 2798 16678 2808 16734
rect 2864 16678 2932 16734
rect 2988 16678 3056 16734
rect 3112 16678 3180 16734
rect 3236 16678 3304 16734
rect 3360 16678 3428 16734
rect 3484 16678 3552 16734
rect 3608 16678 3676 16734
rect 3732 16678 3800 16734
rect 3856 16678 3924 16734
rect 3980 16678 4048 16734
rect 4104 16678 4172 16734
rect 4228 16678 4296 16734
rect 4352 16678 4420 16734
rect 4476 16678 4544 16734
rect 4600 16678 4668 16734
rect 4724 16678 4734 16734
rect 2798 16610 4734 16678
rect 2798 16554 2808 16610
rect 2864 16554 2932 16610
rect 2988 16554 3056 16610
rect 3112 16554 3180 16610
rect 3236 16554 3304 16610
rect 3360 16554 3428 16610
rect 3484 16554 3552 16610
rect 3608 16554 3676 16610
rect 3732 16554 3800 16610
rect 3856 16554 3924 16610
rect 3980 16554 4048 16610
rect 4104 16554 4172 16610
rect 4228 16554 4296 16610
rect 4352 16554 4420 16610
rect 4476 16554 4544 16610
rect 4600 16554 4668 16610
rect 4724 16554 4734 16610
rect 2798 16486 4734 16554
rect 2798 16430 2808 16486
rect 2864 16430 2932 16486
rect 2988 16430 3056 16486
rect 3112 16430 3180 16486
rect 3236 16430 3304 16486
rect 3360 16430 3428 16486
rect 3484 16430 3552 16486
rect 3608 16430 3676 16486
rect 3732 16430 3800 16486
rect 3856 16430 3924 16486
rect 3980 16430 4048 16486
rect 4104 16430 4172 16486
rect 4228 16430 4296 16486
rect 4352 16430 4420 16486
rect 4476 16430 4544 16486
rect 4600 16430 4668 16486
rect 4724 16430 4734 16486
rect 2798 16362 4734 16430
rect 2798 16306 2808 16362
rect 2864 16306 2932 16362
rect 2988 16306 3056 16362
rect 3112 16306 3180 16362
rect 3236 16306 3304 16362
rect 3360 16306 3428 16362
rect 3484 16306 3552 16362
rect 3608 16306 3676 16362
rect 3732 16306 3800 16362
rect 3856 16306 3924 16362
rect 3980 16306 4048 16362
rect 4104 16306 4172 16362
rect 4228 16306 4296 16362
rect 4352 16306 4420 16362
rect 4476 16306 4544 16362
rect 4600 16306 4668 16362
rect 4724 16306 4734 16362
rect 2798 16238 4734 16306
rect 2798 16182 2808 16238
rect 2864 16182 2932 16238
rect 2988 16182 3056 16238
rect 3112 16182 3180 16238
rect 3236 16182 3304 16238
rect 3360 16182 3428 16238
rect 3484 16182 3552 16238
rect 3608 16182 3676 16238
rect 3732 16182 3800 16238
rect 3856 16182 3924 16238
rect 3980 16182 4048 16238
rect 4104 16182 4172 16238
rect 4228 16182 4296 16238
rect 4352 16182 4420 16238
rect 4476 16182 4544 16238
rect 4600 16182 4668 16238
rect 4724 16182 4734 16238
rect 2798 16114 4734 16182
rect 2798 16058 2808 16114
rect 2864 16058 2932 16114
rect 2988 16058 3056 16114
rect 3112 16058 3180 16114
rect 3236 16058 3304 16114
rect 3360 16058 3428 16114
rect 3484 16058 3552 16114
rect 3608 16058 3676 16114
rect 3732 16058 3800 16114
rect 3856 16058 3924 16114
rect 3980 16058 4048 16114
rect 4104 16058 4172 16114
rect 4228 16058 4296 16114
rect 4352 16058 4420 16114
rect 4476 16058 4544 16114
rect 4600 16058 4668 16114
rect 4724 16058 4734 16114
rect 2798 15990 4734 16058
rect 2798 15934 2808 15990
rect 2864 15934 2932 15990
rect 2988 15934 3056 15990
rect 3112 15934 3180 15990
rect 3236 15934 3304 15990
rect 3360 15934 3428 15990
rect 3484 15934 3552 15990
rect 3608 15934 3676 15990
rect 3732 15934 3800 15990
rect 3856 15934 3924 15990
rect 3980 15934 4048 15990
rect 4104 15934 4172 15990
rect 4228 15934 4296 15990
rect 4352 15934 4420 15990
rect 4476 15934 4544 15990
rect 4600 15934 4668 15990
rect 4724 15934 4734 15990
rect 2798 15866 4734 15934
rect 2798 15810 2808 15866
rect 2864 15810 2932 15866
rect 2988 15810 3056 15866
rect 3112 15810 3180 15866
rect 3236 15810 3304 15866
rect 3360 15810 3428 15866
rect 3484 15810 3552 15866
rect 3608 15810 3676 15866
rect 3732 15810 3800 15866
rect 3856 15810 3924 15866
rect 3980 15810 4048 15866
rect 4104 15810 4172 15866
rect 4228 15810 4296 15866
rect 4352 15810 4420 15866
rect 4476 15810 4544 15866
rect 4600 15810 4668 15866
rect 4724 15810 4734 15866
rect 2798 15742 4734 15810
rect 2798 15686 2808 15742
rect 2864 15686 2932 15742
rect 2988 15686 3056 15742
rect 3112 15686 3180 15742
rect 3236 15686 3304 15742
rect 3360 15686 3428 15742
rect 3484 15686 3552 15742
rect 3608 15686 3676 15742
rect 3732 15686 3800 15742
rect 3856 15686 3924 15742
rect 3980 15686 4048 15742
rect 4104 15686 4172 15742
rect 4228 15686 4296 15742
rect 4352 15686 4420 15742
rect 4476 15686 4544 15742
rect 4600 15686 4668 15742
rect 4724 15686 4734 15742
rect 2798 15618 4734 15686
rect 2798 15562 2808 15618
rect 2864 15562 2932 15618
rect 2988 15562 3056 15618
rect 3112 15562 3180 15618
rect 3236 15562 3304 15618
rect 3360 15562 3428 15618
rect 3484 15562 3552 15618
rect 3608 15562 3676 15618
rect 3732 15562 3800 15618
rect 3856 15562 3924 15618
rect 3980 15562 4048 15618
rect 4104 15562 4172 15618
rect 4228 15562 4296 15618
rect 4352 15562 4420 15618
rect 4476 15562 4544 15618
rect 4600 15562 4668 15618
rect 4724 15562 4734 15618
rect 2798 15494 4734 15562
rect 2798 15438 2808 15494
rect 2864 15438 2932 15494
rect 2988 15438 3056 15494
rect 3112 15438 3180 15494
rect 3236 15438 3304 15494
rect 3360 15438 3428 15494
rect 3484 15438 3552 15494
rect 3608 15438 3676 15494
rect 3732 15438 3800 15494
rect 3856 15438 3924 15494
rect 3980 15438 4048 15494
rect 4104 15438 4172 15494
rect 4228 15438 4296 15494
rect 4352 15438 4420 15494
rect 4476 15438 4544 15494
rect 4600 15438 4668 15494
rect 4724 15438 4734 15494
rect 2798 15370 4734 15438
rect 2798 15314 2808 15370
rect 2864 15314 2932 15370
rect 2988 15314 3056 15370
rect 3112 15314 3180 15370
rect 3236 15314 3304 15370
rect 3360 15314 3428 15370
rect 3484 15314 3552 15370
rect 3608 15314 3676 15370
rect 3732 15314 3800 15370
rect 3856 15314 3924 15370
rect 3980 15314 4048 15370
rect 4104 15314 4172 15370
rect 4228 15314 4296 15370
rect 4352 15314 4420 15370
rect 4476 15314 4544 15370
rect 4600 15314 4668 15370
rect 4724 15314 4734 15370
rect 2798 15246 4734 15314
rect 2798 15190 2808 15246
rect 2864 15190 2932 15246
rect 2988 15190 3056 15246
rect 3112 15190 3180 15246
rect 3236 15190 3304 15246
rect 3360 15190 3428 15246
rect 3484 15190 3552 15246
rect 3608 15190 3676 15246
rect 3732 15190 3800 15246
rect 3856 15190 3924 15246
rect 3980 15190 4048 15246
rect 4104 15190 4172 15246
rect 4228 15190 4296 15246
rect 4352 15190 4420 15246
rect 4476 15190 4544 15246
rect 4600 15190 4668 15246
rect 4724 15190 4734 15246
rect 2798 15122 4734 15190
rect 2798 15066 2808 15122
rect 2864 15066 2932 15122
rect 2988 15066 3056 15122
rect 3112 15066 3180 15122
rect 3236 15066 3304 15122
rect 3360 15066 3428 15122
rect 3484 15066 3552 15122
rect 3608 15066 3676 15122
rect 3732 15066 3800 15122
rect 3856 15066 3924 15122
rect 3980 15066 4048 15122
rect 4104 15066 4172 15122
rect 4228 15066 4296 15122
rect 4352 15066 4420 15122
rect 4476 15066 4544 15122
rect 4600 15066 4668 15122
rect 4724 15066 4734 15122
rect 2798 14998 4734 15066
rect 2798 14942 2808 14998
rect 2864 14942 2932 14998
rect 2988 14942 3056 14998
rect 3112 14942 3180 14998
rect 3236 14942 3304 14998
rect 3360 14942 3428 14998
rect 3484 14942 3552 14998
rect 3608 14942 3676 14998
rect 3732 14942 3800 14998
rect 3856 14942 3924 14998
rect 3980 14942 4048 14998
rect 4104 14942 4172 14998
rect 4228 14942 4296 14998
rect 4352 14942 4420 14998
rect 4476 14942 4544 14998
rect 4600 14942 4668 14998
rect 4724 14942 4734 14998
rect 2798 14874 4734 14942
rect 2798 14818 2808 14874
rect 2864 14818 2932 14874
rect 2988 14818 3056 14874
rect 3112 14818 3180 14874
rect 3236 14818 3304 14874
rect 3360 14818 3428 14874
rect 3484 14818 3552 14874
rect 3608 14818 3676 14874
rect 3732 14818 3800 14874
rect 3856 14818 3924 14874
rect 3980 14818 4048 14874
rect 4104 14818 4172 14874
rect 4228 14818 4296 14874
rect 4352 14818 4420 14874
rect 4476 14818 4544 14874
rect 4600 14818 4668 14874
rect 4724 14818 4734 14874
rect 2798 14750 4734 14818
rect 2798 14694 2808 14750
rect 2864 14694 2932 14750
rect 2988 14694 3056 14750
rect 3112 14694 3180 14750
rect 3236 14694 3304 14750
rect 3360 14694 3428 14750
rect 3484 14694 3552 14750
rect 3608 14694 3676 14750
rect 3732 14694 3800 14750
rect 3856 14694 3924 14750
rect 3980 14694 4048 14750
rect 4104 14694 4172 14750
rect 4228 14694 4296 14750
rect 4352 14694 4420 14750
rect 4476 14694 4544 14750
rect 4600 14694 4668 14750
rect 4724 14694 4734 14750
rect 2798 14626 4734 14694
rect 2798 14570 2808 14626
rect 2864 14570 2932 14626
rect 2988 14570 3056 14626
rect 3112 14570 3180 14626
rect 3236 14570 3304 14626
rect 3360 14570 3428 14626
rect 3484 14570 3552 14626
rect 3608 14570 3676 14626
rect 3732 14570 3800 14626
rect 3856 14570 3924 14626
rect 3980 14570 4048 14626
rect 4104 14570 4172 14626
rect 4228 14570 4296 14626
rect 4352 14570 4420 14626
rect 4476 14570 4544 14626
rect 4600 14570 4668 14626
rect 4724 14570 4734 14626
rect 2798 14502 4734 14570
rect 2798 14446 2808 14502
rect 2864 14446 2932 14502
rect 2988 14446 3056 14502
rect 3112 14446 3180 14502
rect 3236 14446 3304 14502
rect 3360 14446 3428 14502
rect 3484 14446 3552 14502
rect 3608 14446 3676 14502
rect 3732 14446 3800 14502
rect 3856 14446 3924 14502
rect 3980 14446 4048 14502
rect 4104 14446 4172 14502
rect 4228 14446 4296 14502
rect 4352 14446 4420 14502
rect 4476 14446 4544 14502
rect 4600 14446 4668 14502
rect 4724 14446 4734 14502
rect 2798 14436 4734 14446
rect 5168 17354 7104 17364
rect 5168 17298 5178 17354
rect 5234 17298 5302 17354
rect 5358 17298 5426 17354
rect 5482 17298 5550 17354
rect 5606 17298 5674 17354
rect 5730 17298 5798 17354
rect 5854 17298 5922 17354
rect 5978 17298 6046 17354
rect 6102 17298 6170 17354
rect 6226 17298 6294 17354
rect 6350 17298 6418 17354
rect 6474 17298 6542 17354
rect 6598 17298 6666 17354
rect 6722 17298 6790 17354
rect 6846 17298 6914 17354
rect 6970 17298 7038 17354
rect 7094 17298 7104 17354
rect 5168 17230 7104 17298
rect 5168 17174 5178 17230
rect 5234 17174 5302 17230
rect 5358 17174 5426 17230
rect 5482 17174 5550 17230
rect 5606 17174 5674 17230
rect 5730 17174 5798 17230
rect 5854 17174 5922 17230
rect 5978 17174 6046 17230
rect 6102 17174 6170 17230
rect 6226 17174 6294 17230
rect 6350 17174 6418 17230
rect 6474 17174 6542 17230
rect 6598 17174 6666 17230
rect 6722 17174 6790 17230
rect 6846 17174 6914 17230
rect 6970 17174 7038 17230
rect 7094 17174 7104 17230
rect 5168 17106 7104 17174
rect 5168 17050 5178 17106
rect 5234 17050 5302 17106
rect 5358 17050 5426 17106
rect 5482 17050 5550 17106
rect 5606 17050 5674 17106
rect 5730 17050 5798 17106
rect 5854 17050 5922 17106
rect 5978 17050 6046 17106
rect 6102 17050 6170 17106
rect 6226 17050 6294 17106
rect 6350 17050 6418 17106
rect 6474 17050 6542 17106
rect 6598 17050 6666 17106
rect 6722 17050 6790 17106
rect 6846 17050 6914 17106
rect 6970 17050 7038 17106
rect 7094 17050 7104 17106
rect 5168 16982 7104 17050
rect 5168 16926 5178 16982
rect 5234 16926 5302 16982
rect 5358 16926 5426 16982
rect 5482 16926 5550 16982
rect 5606 16926 5674 16982
rect 5730 16926 5798 16982
rect 5854 16926 5922 16982
rect 5978 16926 6046 16982
rect 6102 16926 6170 16982
rect 6226 16926 6294 16982
rect 6350 16926 6418 16982
rect 6474 16926 6542 16982
rect 6598 16926 6666 16982
rect 6722 16926 6790 16982
rect 6846 16926 6914 16982
rect 6970 16926 7038 16982
rect 7094 16926 7104 16982
rect 5168 16858 7104 16926
rect 5168 16802 5178 16858
rect 5234 16802 5302 16858
rect 5358 16802 5426 16858
rect 5482 16802 5550 16858
rect 5606 16802 5674 16858
rect 5730 16802 5798 16858
rect 5854 16802 5922 16858
rect 5978 16802 6046 16858
rect 6102 16802 6170 16858
rect 6226 16802 6294 16858
rect 6350 16802 6418 16858
rect 6474 16802 6542 16858
rect 6598 16802 6666 16858
rect 6722 16802 6790 16858
rect 6846 16802 6914 16858
rect 6970 16802 7038 16858
rect 7094 16802 7104 16858
rect 5168 16734 7104 16802
rect 5168 16678 5178 16734
rect 5234 16678 5302 16734
rect 5358 16678 5426 16734
rect 5482 16678 5550 16734
rect 5606 16678 5674 16734
rect 5730 16678 5798 16734
rect 5854 16678 5922 16734
rect 5978 16678 6046 16734
rect 6102 16678 6170 16734
rect 6226 16678 6294 16734
rect 6350 16678 6418 16734
rect 6474 16678 6542 16734
rect 6598 16678 6666 16734
rect 6722 16678 6790 16734
rect 6846 16678 6914 16734
rect 6970 16678 7038 16734
rect 7094 16678 7104 16734
rect 5168 16610 7104 16678
rect 5168 16554 5178 16610
rect 5234 16554 5302 16610
rect 5358 16554 5426 16610
rect 5482 16554 5550 16610
rect 5606 16554 5674 16610
rect 5730 16554 5798 16610
rect 5854 16554 5922 16610
rect 5978 16554 6046 16610
rect 6102 16554 6170 16610
rect 6226 16554 6294 16610
rect 6350 16554 6418 16610
rect 6474 16554 6542 16610
rect 6598 16554 6666 16610
rect 6722 16554 6790 16610
rect 6846 16554 6914 16610
rect 6970 16554 7038 16610
rect 7094 16554 7104 16610
rect 5168 16486 7104 16554
rect 5168 16430 5178 16486
rect 5234 16430 5302 16486
rect 5358 16430 5426 16486
rect 5482 16430 5550 16486
rect 5606 16430 5674 16486
rect 5730 16430 5798 16486
rect 5854 16430 5922 16486
rect 5978 16430 6046 16486
rect 6102 16430 6170 16486
rect 6226 16430 6294 16486
rect 6350 16430 6418 16486
rect 6474 16430 6542 16486
rect 6598 16430 6666 16486
rect 6722 16430 6790 16486
rect 6846 16430 6914 16486
rect 6970 16430 7038 16486
rect 7094 16430 7104 16486
rect 5168 16362 7104 16430
rect 5168 16306 5178 16362
rect 5234 16306 5302 16362
rect 5358 16306 5426 16362
rect 5482 16306 5550 16362
rect 5606 16306 5674 16362
rect 5730 16306 5798 16362
rect 5854 16306 5922 16362
rect 5978 16306 6046 16362
rect 6102 16306 6170 16362
rect 6226 16306 6294 16362
rect 6350 16306 6418 16362
rect 6474 16306 6542 16362
rect 6598 16306 6666 16362
rect 6722 16306 6790 16362
rect 6846 16306 6914 16362
rect 6970 16306 7038 16362
rect 7094 16306 7104 16362
rect 5168 16238 7104 16306
rect 5168 16182 5178 16238
rect 5234 16182 5302 16238
rect 5358 16182 5426 16238
rect 5482 16182 5550 16238
rect 5606 16182 5674 16238
rect 5730 16182 5798 16238
rect 5854 16182 5922 16238
rect 5978 16182 6046 16238
rect 6102 16182 6170 16238
rect 6226 16182 6294 16238
rect 6350 16182 6418 16238
rect 6474 16182 6542 16238
rect 6598 16182 6666 16238
rect 6722 16182 6790 16238
rect 6846 16182 6914 16238
rect 6970 16182 7038 16238
rect 7094 16182 7104 16238
rect 5168 16114 7104 16182
rect 5168 16058 5178 16114
rect 5234 16058 5302 16114
rect 5358 16058 5426 16114
rect 5482 16058 5550 16114
rect 5606 16058 5674 16114
rect 5730 16058 5798 16114
rect 5854 16058 5922 16114
rect 5978 16058 6046 16114
rect 6102 16058 6170 16114
rect 6226 16058 6294 16114
rect 6350 16058 6418 16114
rect 6474 16058 6542 16114
rect 6598 16058 6666 16114
rect 6722 16058 6790 16114
rect 6846 16058 6914 16114
rect 6970 16058 7038 16114
rect 7094 16058 7104 16114
rect 5168 15990 7104 16058
rect 5168 15934 5178 15990
rect 5234 15934 5302 15990
rect 5358 15934 5426 15990
rect 5482 15934 5550 15990
rect 5606 15934 5674 15990
rect 5730 15934 5798 15990
rect 5854 15934 5922 15990
rect 5978 15934 6046 15990
rect 6102 15934 6170 15990
rect 6226 15934 6294 15990
rect 6350 15934 6418 15990
rect 6474 15934 6542 15990
rect 6598 15934 6666 15990
rect 6722 15934 6790 15990
rect 6846 15934 6914 15990
rect 6970 15934 7038 15990
rect 7094 15934 7104 15990
rect 5168 15866 7104 15934
rect 5168 15810 5178 15866
rect 5234 15810 5302 15866
rect 5358 15810 5426 15866
rect 5482 15810 5550 15866
rect 5606 15810 5674 15866
rect 5730 15810 5798 15866
rect 5854 15810 5922 15866
rect 5978 15810 6046 15866
rect 6102 15810 6170 15866
rect 6226 15810 6294 15866
rect 6350 15810 6418 15866
rect 6474 15810 6542 15866
rect 6598 15810 6666 15866
rect 6722 15810 6790 15866
rect 6846 15810 6914 15866
rect 6970 15810 7038 15866
rect 7094 15810 7104 15866
rect 5168 15742 7104 15810
rect 5168 15686 5178 15742
rect 5234 15686 5302 15742
rect 5358 15686 5426 15742
rect 5482 15686 5550 15742
rect 5606 15686 5674 15742
rect 5730 15686 5798 15742
rect 5854 15686 5922 15742
rect 5978 15686 6046 15742
rect 6102 15686 6170 15742
rect 6226 15686 6294 15742
rect 6350 15686 6418 15742
rect 6474 15686 6542 15742
rect 6598 15686 6666 15742
rect 6722 15686 6790 15742
rect 6846 15686 6914 15742
rect 6970 15686 7038 15742
rect 7094 15686 7104 15742
rect 5168 15618 7104 15686
rect 5168 15562 5178 15618
rect 5234 15562 5302 15618
rect 5358 15562 5426 15618
rect 5482 15562 5550 15618
rect 5606 15562 5674 15618
rect 5730 15562 5798 15618
rect 5854 15562 5922 15618
rect 5978 15562 6046 15618
rect 6102 15562 6170 15618
rect 6226 15562 6294 15618
rect 6350 15562 6418 15618
rect 6474 15562 6542 15618
rect 6598 15562 6666 15618
rect 6722 15562 6790 15618
rect 6846 15562 6914 15618
rect 6970 15562 7038 15618
rect 7094 15562 7104 15618
rect 5168 15494 7104 15562
rect 5168 15438 5178 15494
rect 5234 15438 5302 15494
rect 5358 15438 5426 15494
rect 5482 15438 5550 15494
rect 5606 15438 5674 15494
rect 5730 15438 5798 15494
rect 5854 15438 5922 15494
rect 5978 15438 6046 15494
rect 6102 15438 6170 15494
rect 6226 15438 6294 15494
rect 6350 15438 6418 15494
rect 6474 15438 6542 15494
rect 6598 15438 6666 15494
rect 6722 15438 6790 15494
rect 6846 15438 6914 15494
rect 6970 15438 7038 15494
rect 7094 15438 7104 15494
rect 5168 15370 7104 15438
rect 5168 15314 5178 15370
rect 5234 15314 5302 15370
rect 5358 15314 5426 15370
rect 5482 15314 5550 15370
rect 5606 15314 5674 15370
rect 5730 15314 5798 15370
rect 5854 15314 5922 15370
rect 5978 15314 6046 15370
rect 6102 15314 6170 15370
rect 6226 15314 6294 15370
rect 6350 15314 6418 15370
rect 6474 15314 6542 15370
rect 6598 15314 6666 15370
rect 6722 15314 6790 15370
rect 6846 15314 6914 15370
rect 6970 15314 7038 15370
rect 7094 15314 7104 15370
rect 5168 15246 7104 15314
rect 5168 15190 5178 15246
rect 5234 15190 5302 15246
rect 5358 15190 5426 15246
rect 5482 15190 5550 15246
rect 5606 15190 5674 15246
rect 5730 15190 5798 15246
rect 5854 15190 5922 15246
rect 5978 15190 6046 15246
rect 6102 15190 6170 15246
rect 6226 15190 6294 15246
rect 6350 15190 6418 15246
rect 6474 15190 6542 15246
rect 6598 15190 6666 15246
rect 6722 15190 6790 15246
rect 6846 15190 6914 15246
rect 6970 15190 7038 15246
rect 7094 15190 7104 15246
rect 5168 15122 7104 15190
rect 5168 15066 5178 15122
rect 5234 15066 5302 15122
rect 5358 15066 5426 15122
rect 5482 15066 5550 15122
rect 5606 15066 5674 15122
rect 5730 15066 5798 15122
rect 5854 15066 5922 15122
rect 5978 15066 6046 15122
rect 6102 15066 6170 15122
rect 6226 15066 6294 15122
rect 6350 15066 6418 15122
rect 6474 15066 6542 15122
rect 6598 15066 6666 15122
rect 6722 15066 6790 15122
rect 6846 15066 6914 15122
rect 6970 15066 7038 15122
rect 7094 15066 7104 15122
rect 5168 14998 7104 15066
rect 5168 14942 5178 14998
rect 5234 14942 5302 14998
rect 5358 14942 5426 14998
rect 5482 14942 5550 14998
rect 5606 14942 5674 14998
rect 5730 14942 5798 14998
rect 5854 14942 5922 14998
rect 5978 14942 6046 14998
rect 6102 14942 6170 14998
rect 6226 14942 6294 14998
rect 6350 14942 6418 14998
rect 6474 14942 6542 14998
rect 6598 14942 6666 14998
rect 6722 14942 6790 14998
rect 6846 14942 6914 14998
rect 6970 14942 7038 14998
rect 7094 14942 7104 14998
rect 5168 14874 7104 14942
rect 5168 14818 5178 14874
rect 5234 14818 5302 14874
rect 5358 14818 5426 14874
rect 5482 14818 5550 14874
rect 5606 14818 5674 14874
rect 5730 14818 5798 14874
rect 5854 14818 5922 14874
rect 5978 14818 6046 14874
rect 6102 14818 6170 14874
rect 6226 14818 6294 14874
rect 6350 14818 6418 14874
rect 6474 14818 6542 14874
rect 6598 14818 6666 14874
rect 6722 14818 6790 14874
rect 6846 14818 6914 14874
rect 6970 14818 7038 14874
rect 7094 14818 7104 14874
rect 5168 14750 7104 14818
rect 5168 14694 5178 14750
rect 5234 14694 5302 14750
rect 5358 14694 5426 14750
rect 5482 14694 5550 14750
rect 5606 14694 5674 14750
rect 5730 14694 5798 14750
rect 5854 14694 5922 14750
rect 5978 14694 6046 14750
rect 6102 14694 6170 14750
rect 6226 14694 6294 14750
rect 6350 14694 6418 14750
rect 6474 14694 6542 14750
rect 6598 14694 6666 14750
rect 6722 14694 6790 14750
rect 6846 14694 6914 14750
rect 6970 14694 7038 14750
rect 7094 14694 7104 14750
rect 5168 14626 7104 14694
rect 5168 14570 5178 14626
rect 5234 14570 5302 14626
rect 5358 14570 5426 14626
rect 5482 14570 5550 14626
rect 5606 14570 5674 14626
rect 5730 14570 5798 14626
rect 5854 14570 5922 14626
rect 5978 14570 6046 14626
rect 6102 14570 6170 14626
rect 6226 14570 6294 14626
rect 6350 14570 6418 14626
rect 6474 14570 6542 14626
rect 6598 14570 6666 14626
rect 6722 14570 6790 14626
rect 6846 14570 6914 14626
rect 6970 14570 7038 14626
rect 7094 14570 7104 14626
rect 5168 14502 7104 14570
rect 5168 14446 5178 14502
rect 5234 14446 5302 14502
rect 5358 14446 5426 14502
rect 5482 14446 5550 14502
rect 5606 14446 5674 14502
rect 5730 14446 5798 14502
rect 5854 14446 5922 14502
rect 5978 14446 6046 14502
rect 6102 14446 6170 14502
rect 6226 14446 6294 14502
rect 6350 14446 6418 14502
rect 6474 14446 6542 14502
rect 6598 14446 6666 14502
rect 6722 14446 6790 14502
rect 6846 14446 6914 14502
rect 6970 14446 7038 14502
rect 7094 14446 7104 14502
rect 5168 14436 7104 14446
rect 7874 17354 9810 17364
rect 7874 17298 7884 17354
rect 7940 17298 8008 17354
rect 8064 17298 8132 17354
rect 8188 17298 8256 17354
rect 8312 17298 8380 17354
rect 8436 17298 8504 17354
rect 8560 17298 8628 17354
rect 8684 17298 8752 17354
rect 8808 17298 8876 17354
rect 8932 17298 9000 17354
rect 9056 17298 9124 17354
rect 9180 17298 9248 17354
rect 9304 17298 9372 17354
rect 9428 17298 9496 17354
rect 9552 17298 9620 17354
rect 9676 17298 9744 17354
rect 9800 17298 9810 17354
rect 7874 17230 9810 17298
rect 7874 17174 7884 17230
rect 7940 17174 8008 17230
rect 8064 17174 8132 17230
rect 8188 17174 8256 17230
rect 8312 17174 8380 17230
rect 8436 17174 8504 17230
rect 8560 17174 8628 17230
rect 8684 17174 8752 17230
rect 8808 17174 8876 17230
rect 8932 17174 9000 17230
rect 9056 17174 9124 17230
rect 9180 17174 9248 17230
rect 9304 17174 9372 17230
rect 9428 17174 9496 17230
rect 9552 17174 9620 17230
rect 9676 17174 9744 17230
rect 9800 17174 9810 17230
rect 7874 17106 9810 17174
rect 7874 17050 7884 17106
rect 7940 17050 8008 17106
rect 8064 17050 8132 17106
rect 8188 17050 8256 17106
rect 8312 17050 8380 17106
rect 8436 17050 8504 17106
rect 8560 17050 8628 17106
rect 8684 17050 8752 17106
rect 8808 17050 8876 17106
rect 8932 17050 9000 17106
rect 9056 17050 9124 17106
rect 9180 17050 9248 17106
rect 9304 17050 9372 17106
rect 9428 17050 9496 17106
rect 9552 17050 9620 17106
rect 9676 17050 9744 17106
rect 9800 17050 9810 17106
rect 7874 16982 9810 17050
rect 7874 16926 7884 16982
rect 7940 16926 8008 16982
rect 8064 16926 8132 16982
rect 8188 16926 8256 16982
rect 8312 16926 8380 16982
rect 8436 16926 8504 16982
rect 8560 16926 8628 16982
rect 8684 16926 8752 16982
rect 8808 16926 8876 16982
rect 8932 16926 9000 16982
rect 9056 16926 9124 16982
rect 9180 16926 9248 16982
rect 9304 16926 9372 16982
rect 9428 16926 9496 16982
rect 9552 16926 9620 16982
rect 9676 16926 9744 16982
rect 9800 16926 9810 16982
rect 7874 16858 9810 16926
rect 7874 16802 7884 16858
rect 7940 16802 8008 16858
rect 8064 16802 8132 16858
rect 8188 16802 8256 16858
rect 8312 16802 8380 16858
rect 8436 16802 8504 16858
rect 8560 16802 8628 16858
rect 8684 16802 8752 16858
rect 8808 16802 8876 16858
rect 8932 16802 9000 16858
rect 9056 16802 9124 16858
rect 9180 16802 9248 16858
rect 9304 16802 9372 16858
rect 9428 16802 9496 16858
rect 9552 16802 9620 16858
rect 9676 16802 9744 16858
rect 9800 16802 9810 16858
rect 7874 16734 9810 16802
rect 7874 16678 7884 16734
rect 7940 16678 8008 16734
rect 8064 16678 8132 16734
rect 8188 16678 8256 16734
rect 8312 16678 8380 16734
rect 8436 16678 8504 16734
rect 8560 16678 8628 16734
rect 8684 16678 8752 16734
rect 8808 16678 8876 16734
rect 8932 16678 9000 16734
rect 9056 16678 9124 16734
rect 9180 16678 9248 16734
rect 9304 16678 9372 16734
rect 9428 16678 9496 16734
rect 9552 16678 9620 16734
rect 9676 16678 9744 16734
rect 9800 16678 9810 16734
rect 7874 16610 9810 16678
rect 7874 16554 7884 16610
rect 7940 16554 8008 16610
rect 8064 16554 8132 16610
rect 8188 16554 8256 16610
rect 8312 16554 8380 16610
rect 8436 16554 8504 16610
rect 8560 16554 8628 16610
rect 8684 16554 8752 16610
rect 8808 16554 8876 16610
rect 8932 16554 9000 16610
rect 9056 16554 9124 16610
rect 9180 16554 9248 16610
rect 9304 16554 9372 16610
rect 9428 16554 9496 16610
rect 9552 16554 9620 16610
rect 9676 16554 9744 16610
rect 9800 16554 9810 16610
rect 7874 16486 9810 16554
rect 7874 16430 7884 16486
rect 7940 16430 8008 16486
rect 8064 16430 8132 16486
rect 8188 16430 8256 16486
rect 8312 16430 8380 16486
rect 8436 16430 8504 16486
rect 8560 16430 8628 16486
rect 8684 16430 8752 16486
rect 8808 16430 8876 16486
rect 8932 16430 9000 16486
rect 9056 16430 9124 16486
rect 9180 16430 9248 16486
rect 9304 16430 9372 16486
rect 9428 16430 9496 16486
rect 9552 16430 9620 16486
rect 9676 16430 9744 16486
rect 9800 16430 9810 16486
rect 7874 16362 9810 16430
rect 7874 16306 7884 16362
rect 7940 16306 8008 16362
rect 8064 16306 8132 16362
rect 8188 16306 8256 16362
rect 8312 16306 8380 16362
rect 8436 16306 8504 16362
rect 8560 16306 8628 16362
rect 8684 16306 8752 16362
rect 8808 16306 8876 16362
rect 8932 16306 9000 16362
rect 9056 16306 9124 16362
rect 9180 16306 9248 16362
rect 9304 16306 9372 16362
rect 9428 16306 9496 16362
rect 9552 16306 9620 16362
rect 9676 16306 9744 16362
rect 9800 16306 9810 16362
rect 7874 16238 9810 16306
rect 7874 16182 7884 16238
rect 7940 16182 8008 16238
rect 8064 16182 8132 16238
rect 8188 16182 8256 16238
rect 8312 16182 8380 16238
rect 8436 16182 8504 16238
rect 8560 16182 8628 16238
rect 8684 16182 8752 16238
rect 8808 16182 8876 16238
rect 8932 16182 9000 16238
rect 9056 16182 9124 16238
rect 9180 16182 9248 16238
rect 9304 16182 9372 16238
rect 9428 16182 9496 16238
rect 9552 16182 9620 16238
rect 9676 16182 9744 16238
rect 9800 16182 9810 16238
rect 7874 16114 9810 16182
rect 7874 16058 7884 16114
rect 7940 16058 8008 16114
rect 8064 16058 8132 16114
rect 8188 16058 8256 16114
rect 8312 16058 8380 16114
rect 8436 16058 8504 16114
rect 8560 16058 8628 16114
rect 8684 16058 8752 16114
rect 8808 16058 8876 16114
rect 8932 16058 9000 16114
rect 9056 16058 9124 16114
rect 9180 16058 9248 16114
rect 9304 16058 9372 16114
rect 9428 16058 9496 16114
rect 9552 16058 9620 16114
rect 9676 16058 9744 16114
rect 9800 16058 9810 16114
rect 7874 15990 9810 16058
rect 7874 15934 7884 15990
rect 7940 15934 8008 15990
rect 8064 15934 8132 15990
rect 8188 15934 8256 15990
rect 8312 15934 8380 15990
rect 8436 15934 8504 15990
rect 8560 15934 8628 15990
rect 8684 15934 8752 15990
rect 8808 15934 8876 15990
rect 8932 15934 9000 15990
rect 9056 15934 9124 15990
rect 9180 15934 9248 15990
rect 9304 15934 9372 15990
rect 9428 15934 9496 15990
rect 9552 15934 9620 15990
rect 9676 15934 9744 15990
rect 9800 15934 9810 15990
rect 7874 15866 9810 15934
rect 7874 15810 7884 15866
rect 7940 15810 8008 15866
rect 8064 15810 8132 15866
rect 8188 15810 8256 15866
rect 8312 15810 8380 15866
rect 8436 15810 8504 15866
rect 8560 15810 8628 15866
rect 8684 15810 8752 15866
rect 8808 15810 8876 15866
rect 8932 15810 9000 15866
rect 9056 15810 9124 15866
rect 9180 15810 9248 15866
rect 9304 15810 9372 15866
rect 9428 15810 9496 15866
rect 9552 15810 9620 15866
rect 9676 15810 9744 15866
rect 9800 15810 9810 15866
rect 7874 15742 9810 15810
rect 7874 15686 7884 15742
rect 7940 15686 8008 15742
rect 8064 15686 8132 15742
rect 8188 15686 8256 15742
rect 8312 15686 8380 15742
rect 8436 15686 8504 15742
rect 8560 15686 8628 15742
rect 8684 15686 8752 15742
rect 8808 15686 8876 15742
rect 8932 15686 9000 15742
rect 9056 15686 9124 15742
rect 9180 15686 9248 15742
rect 9304 15686 9372 15742
rect 9428 15686 9496 15742
rect 9552 15686 9620 15742
rect 9676 15686 9744 15742
rect 9800 15686 9810 15742
rect 7874 15618 9810 15686
rect 7874 15562 7884 15618
rect 7940 15562 8008 15618
rect 8064 15562 8132 15618
rect 8188 15562 8256 15618
rect 8312 15562 8380 15618
rect 8436 15562 8504 15618
rect 8560 15562 8628 15618
rect 8684 15562 8752 15618
rect 8808 15562 8876 15618
rect 8932 15562 9000 15618
rect 9056 15562 9124 15618
rect 9180 15562 9248 15618
rect 9304 15562 9372 15618
rect 9428 15562 9496 15618
rect 9552 15562 9620 15618
rect 9676 15562 9744 15618
rect 9800 15562 9810 15618
rect 7874 15494 9810 15562
rect 7874 15438 7884 15494
rect 7940 15438 8008 15494
rect 8064 15438 8132 15494
rect 8188 15438 8256 15494
rect 8312 15438 8380 15494
rect 8436 15438 8504 15494
rect 8560 15438 8628 15494
rect 8684 15438 8752 15494
rect 8808 15438 8876 15494
rect 8932 15438 9000 15494
rect 9056 15438 9124 15494
rect 9180 15438 9248 15494
rect 9304 15438 9372 15494
rect 9428 15438 9496 15494
rect 9552 15438 9620 15494
rect 9676 15438 9744 15494
rect 9800 15438 9810 15494
rect 7874 15370 9810 15438
rect 7874 15314 7884 15370
rect 7940 15314 8008 15370
rect 8064 15314 8132 15370
rect 8188 15314 8256 15370
rect 8312 15314 8380 15370
rect 8436 15314 8504 15370
rect 8560 15314 8628 15370
rect 8684 15314 8752 15370
rect 8808 15314 8876 15370
rect 8932 15314 9000 15370
rect 9056 15314 9124 15370
rect 9180 15314 9248 15370
rect 9304 15314 9372 15370
rect 9428 15314 9496 15370
rect 9552 15314 9620 15370
rect 9676 15314 9744 15370
rect 9800 15314 9810 15370
rect 7874 15246 9810 15314
rect 7874 15190 7884 15246
rect 7940 15190 8008 15246
rect 8064 15190 8132 15246
rect 8188 15190 8256 15246
rect 8312 15190 8380 15246
rect 8436 15190 8504 15246
rect 8560 15190 8628 15246
rect 8684 15190 8752 15246
rect 8808 15190 8876 15246
rect 8932 15190 9000 15246
rect 9056 15190 9124 15246
rect 9180 15190 9248 15246
rect 9304 15190 9372 15246
rect 9428 15190 9496 15246
rect 9552 15190 9620 15246
rect 9676 15190 9744 15246
rect 9800 15190 9810 15246
rect 7874 15122 9810 15190
rect 7874 15066 7884 15122
rect 7940 15066 8008 15122
rect 8064 15066 8132 15122
rect 8188 15066 8256 15122
rect 8312 15066 8380 15122
rect 8436 15066 8504 15122
rect 8560 15066 8628 15122
rect 8684 15066 8752 15122
rect 8808 15066 8876 15122
rect 8932 15066 9000 15122
rect 9056 15066 9124 15122
rect 9180 15066 9248 15122
rect 9304 15066 9372 15122
rect 9428 15066 9496 15122
rect 9552 15066 9620 15122
rect 9676 15066 9744 15122
rect 9800 15066 9810 15122
rect 7874 14998 9810 15066
rect 7874 14942 7884 14998
rect 7940 14942 8008 14998
rect 8064 14942 8132 14998
rect 8188 14942 8256 14998
rect 8312 14942 8380 14998
rect 8436 14942 8504 14998
rect 8560 14942 8628 14998
rect 8684 14942 8752 14998
rect 8808 14942 8876 14998
rect 8932 14942 9000 14998
rect 9056 14942 9124 14998
rect 9180 14942 9248 14998
rect 9304 14942 9372 14998
rect 9428 14942 9496 14998
rect 9552 14942 9620 14998
rect 9676 14942 9744 14998
rect 9800 14942 9810 14998
rect 7874 14874 9810 14942
rect 7874 14818 7884 14874
rect 7940 14818 8008 14874
rect 8064 14818 8132 14874
rect 8188 14818 8256 14874
rect 8312 14818 8380 14874
rect 8436 14818 8504 14874
rect 8560 14818 8628 14874
rect 8684 14818 8752 14874
rect 8808 14818 8876 14874
rect 8932 14818 9000 14874
rect 9056 14818 9124 14874
rect 9180 14818 9248 14874
rect 9304 14818 9372 14874
rect 9428 14818 9496 14874
rect 9552 14818 9620 14874
rect 9676 14818 9744 14874
rect 9800 14818 9810 14874
rect 7874 14750 9810 14818
rect 7874 14694 7884 14750
rect 7940 14694 8008 14750
rect 8064 14694 8132 14750
rect 8188 14694 8256 14750
rect 8312 14694 8380 14750
rect 8436 14694 8504 14750
rect 8560 14694 8628 14750
rect 8684 14694 8752 14750
rect 8808 14694 8876 14750
rect 8932 14694 9000 14750
rect 9056 14694 9124 14750
rect 9180 14694 9248 14750
rect 9304 14694 9372 14750
rect 9428 14694 9496 14750
rect 9552 14694 9620 14750
rect 9676 14694 9744 14750
rect 9800 14694 9810 14750
rect 7874 14626 9810 14694
rect 7874 14570 7884 14626
rect 7940 14570 8008 14626
rect 8064 14570 8132 14626
rect 8188 14570 8256 14626
rect 8312 14570 8380 14626
rect 8436 14570 8504 14626
rect 8560 14570 8628 14626
rect 8684 14570 8752 14626
rect 8808 14570 8876 14626
rect 8932 14570 9000 14626
rect 9056 14570 9124 14626
rect 9180 14570 9248 14626
rect 9304 14570 9372 14626
rect 9428 14570 9496 14626
rect 9552 14570 9620 14626
rect 9676 14570 9744 14626
rect 9800 14570 9810 14626
rect 7874 14502 9810 14570
rect 7874 14446 7884 14502
rect 7940 14446 8008 14502
rect 8064 14446 8132 14502
rect 8188 14446 8256 14502
rect 8312 14446 8380 14502
rect 8436 14446 8504 14502
rect 8560 14446 8628 14502
rect 8684 14446 8752 14502
rect 8808 14446 8876 14502
rect 8932 14446 9000 14502
rect 9056 14446 9124 14502
rect 9180 14446 9248 14502
rect 9304 14446 9372 14502
rect 9428 14446 9496 14502
rect 9552 14446 9620 14502
rect 9676 14446 9744 14502
rect 9800 14446 9810 14502
rect 7874 14436 9810 14446
rect 10244 17354 12180 17364
rect 10244 17298 10254 17354
rect 10310 17298 10378 17354
rect 10434 17298 10502 17354
rect 10558 17298 10626 17354
rect 10682 17298 10750 17354
rect 10806 17298 10874 17354
rect 10930 17298 10998 17354
rect 11054 17298 11122 17354
rect 11178 17298 11246 17354
rect 11302 17298 11370 17354
rect 11426 17298 11494 17354
rect 11550 17298 11618 17354
rect 11674 17298 11742 17354
rect 11798 17298 11866 17354
rect 11922 17298 11990 17354
rect 12046 17298 12114 17354
rect 12170 17298 12180 17354
rect 10244 17230 12180 17298
rect 10244 17174 10254 17230
rect 10310 17174 10378 17230
rect 10434 17174 10502 17230
rect 10558 17174 10626 17230
rect 10682 17174 10750 17230
rect 10806 17174 10874 17230
rect 10930 17174 10998 17230
rect 11054 17174 11122 17230
rect 11178 17174 11246 17230
rect 11302 17174 11370 17230
rect 11426 17174 11494 17230
rect 11550 17174 11618 17230
rect 11674 17174 11742 17230
rect 11798 17174 11866 17230
rect 11922 17174 11990 17230
rect 12046 17174 12114 17230
rect 12170 17174 12180 17230
rect 10244 17106 12180 17174
rect 10244 17050 10254 17106
rect 10310 17050 10378 17106
rect 10434 17050 10502 17106
rect 10558 17050 10626 17106
rect 10682 17050 10750 17106
rect 10806 17050 10874 17106
rect 10930 17050 10998 17106
rect 11054 17050 11122 17106
rect 11178 17050 11246 17106
rect 11302 17050 11370 17106
rect 11426 17050 11494 17106
rect 11550 17050 11618 17106
rect 11674 17050 11742 17106
rect 11798 17050 11866 17106
rect 11922 17050 11990 17106
rect 12046 17050 12114 17106
rect 12170 17050 12180 17106
rect 10244 16982 12180 17050
rect 10244 16926 10254 16982
rect 10310 16926 10378 16982
rect 10434 16926 10502 16982
rect 10558 16926 10626 16982
rect 10682 16926 10750 16982
rect 10806 16926 10874 16982
rect 10930 16926 10998 16982
rect 11054 16926 11122 16982
rect 11178 16926 11246 16982
rect 11302 16926 11370 16982
rect 11426 16926 11494 16982
rect 11550 16926 11618 16982
rect 11674 16926 11742 16982
rect 11798 16926 11866 16982
rect 11922 16926 11990 16982
rect 12046 16926 12114 16982
rect 12170 16926 12180 16982
rect 10244 16858 12180 16926
rect 10244 16802 10254 16858
rect 10310 16802 10378 16858
rect 10434 16802 10502 16858
rect 10558 16802 10626 16858
rect 10682 16802 10750 16858
rect 10806 16802 10874 16858
rect 10930 16802 10998 16858
rect 11054 16802 11122 16858
rect 11178 16802 11246 16858
rect 11302 16802 11370 16858
rect 11426 16802 11494 16858
rect 11550 16802 11618 16858
rect 11674 16802 11742 16858
rect 11798 16802 11866 16858
rect 11922 16802 11990 16858
rect 12046 16802 12114 16858
rect 12170 16802 12180 16858
rect 10244 16734 12180 16802
rect 10244 16678 10254 16734
rect 10310 16678 10378 16734
rect 10434 16678 10502 16734
rect 10558 16678 10626 16734
rect 10682 16678 10750 16734
rect 10806 16678 10874 16734
rect 10930 16678 10998 16734
rect 11054 16678 11122 16734
rect 11178 16678 11246 16734
rect 11302 16678 11370 16734
rect 11426 16678 11494 16734
rect 11550 16678 11618 16734
rect 11674 16678 11742 16734
rect 11798 16678 11866 16734
rect 11922 16678 11990 16734
rect 12046 16678 12114 16734
rect 12170 16678 12180 16734
rect 10244 16610 12180 16678
rect 10244 16554 10254 16610
rect 10310 16554 10378 16610
rect 10434 16554 10502 16610
rect 10558 16554 10626 16610
rect 10682 16554 10750 16610
rect 10806 16554 10874 16610
rect 10930 16554 10998 16610
rect 11054 16554 11122 16610
rect 11178 16554 11246 16610
rect 11302 16554 11370 16610
rect 11426 16554 11494 16610
rect 11550 16554 11618 16610
rect 11674 16554 11742 16610
rect 11798 16554 11866 16610
rect 11922 16554 11990 16610
rect 12046 16554 12114 16610
rect 12170 16554 12180 16610
rect 10244 16486 12180 16554
rect 10244 16430 10254 16486
rect 10310 16430 10378 16486
rect 10434 16430 10502 16486
rect 10558 16430 10626 16486
rect 10682 16430 10750 16486
rect 10806 16430 10874 16486
rect 10930 16430 10998 16486
rect 11054 16430 11122 16486
rect 11178 16430 11246 16486
rect 11302 16430 11370 16486
rect 11426 16430 11494 16486
rect 11550 16430 11618 16486
rect 11674 16430 11742 16486
rect 11798 16430 11866 16486
rect 11922 16430 11990 16486
rect 12046 16430 12114 16486
rect 12170 16430 12180 16486
rect 10244 16362 12180 16430
rect 10244 16306 10254 16362
rect 10310 16306 10378 16362
rect 10434 16306 10502 16362
rect 10558 16306 10626 16362
rect 10682 16306 10750 16362
rect 10806 16306 10874 16362
rect 10930 16306 10998 16362
rect 11054 16306 11122 16362
rect 11178 16306 11246 16362
rect 11302 16306 11370 16362
rect 11426 16306 11494 16362
rect 11550 16306 11618 16362
rect 11674 16306 11742 16362
rect 11798 16306 11866 16362
rect 11922 16306 11990 16362
rect 12046 16306 12114 16362
rect 12170 16306 12180 16362
rect 10244 16238 12180 16306
rect 10244 16182 10254 16238
rect 10310 16182 10378 16238
rect 10434 16182 10502 16238
rect 10558 16182 10626 16238
rect 10682 16182 10750 16238
rect 10806 16182 10874 16238
rect 10930 16182 10998 16238
rect 11054 16182 11122 16238
rect 11178 16182 11246 16238
rect 11302 16182 11370 16238
rect 11426 16182 11494 16238
rect 11550 16182 11618 16238
rect 11674 16182 11742 16238
rect 11798 16182 11866 16238
rect 11922 16182 11990 16238
rect 12046 16182 12114 16238
rect 12170 16182 12180 16238
rect 10244 16114 12180 16182
rect 10244 16058 10254 16114
rect 10310 16058 10378 16114
rect 10434 16058 10502 16114
rect 10558 16058 10626 16114
rect 10682 16058 10750 16114
rect 10806 16058 10874 16114
rect 10930 16058 10998 16114
rect 11054 16058 11122 16114
rect 11178 16058 11246 16114
rect 11302 16058 11370 16114
rect 11426 16058 11494 16114
rect 11550 16058 11618 16114
rect 11674 16058 11742 16114
rect 11798 16058 11866 16114
rect 11922 16058 11990 16114
rect 12046 16058 12114 16114
rect 12170 16058 12180 16114
rect 10244 15990 12180 16058
rect 10244 15934 10254 15990
rect 10310 15934 10378 15990
rect 10434 15934 10502 15990
rect 10558 15934 10626 15990
rect 10682 15934 10750 15990
rect 10806 15934 10874 15990
rect 10930 15934 10998 15990
rect 11054 15934 11122 15990
rect 11178 15934 11246 15990
rect 11302 15934 11370 15990
rect 11426 15934 11494 15990
rect 11550 15934 11618 15990
rect 11674 15934 11742 15990
rect 11798 15934 11866 15990
rect 11922 15934 11990 15990
rect 12046 15934 12114 15990
rect 12170 15934 12180 15990
rect 10244 15866 12180 15934
rect 10244 15810 10254 15866
rect 10310 15810 10378 15866
rect 10434 15810 10502 15866
rect 10558 15810 10626 15866
rect 10682 15810 10750 15866
rect 10806 15810 10874 15866
rect 10930 15810 10998 15866
rect 11054 15810 11122 15866
rect 11178 15810 11246 15866
rect 11302 15810 11370 15866
rect 11426 15810 11494 15866
rect 11550 15810 11618 15866
rect 11674 15810 11742 15866
rect 11798 15810 11866 15866
rect 11922 15810 11990 15866
rect 12046 15810 12114 15866
rect 12170 15810 12180 15866
rect 10244 15742 12180 15810
rect 10244 15686 10254 15742
rect 10310 15686 10378 15742
rect 10434 15686 10502 15742
rect 10558 15686 10626 15742
rect 10682 15686 10750 15742
rect 10806 15686 10874 15742
rect 10930 15686 10998 15742
rect 11054 15686 11122 15742
rect 11178 15686 11246 15742
rect 11302 15686 11370 15742
rect 11426 15686 11494 15742
rect 11550 15686 11618 15742
rect 11674 15686 11742 15742
rect 11798 15686 11866 15742
rect 11922 15686 11990 15742
rect 12046 15686 12114 15742
rect 12170 15686 12180 15742
rect 10244 15618 12180 15686
rect 10244 15562 10254 15618
rect 10310 15562 10378 15618
rect 10434 15562 10502 15618
rect 10558 15562 10626 15618
rect 10682 15562 10750 15618
rect 10806 15562 10874 15618
rect 10930 15562 10998 15618
rect 11054 15562 11122 15618
rect 11178 15562 11246 15618
rect 11302 15562 11370 15618
rect 11426 15562 11494 15618
rect 11550 15562 11618 15618
rect 11674 15562 11742 15618
rect 11798 15562 11866 15618
rect 11922 15562 11990 15618
rect 12046 15562 12114 15618
rect 12170 15562 12180 15618
rect 10244 15494 12180 15562
rect 10244 15438 10254 15494
rect 10310 15438 10378 15494
rect 10434 15438 10502 15494
rect 10558 15438 10626 15494
rect 10682 15438 10750 15494
rect 10806 15438 10874 15494
rect 10930 15438 10998 15494
rect 11054 15438 11122 15494
rect 11178 15438 11246 15494
rect 11302 15438 11370 15494
rect 11426 15438 11494 15494
rect 11550 15438 11618 15494
rect 11674 15438 11742 15494
rect 11798 15438 11866 15494
rect 11922 15438 11990 15494
rect 12046 15438 12114 15494
rect 12170 15438 12180 15494
rect 10244 15370 12180 15438
rect 10244 15314 10254 15370
rect 10310 15314 10378 15370
rect 10434 15314 10502 15370
rect 10558 15314 10626 15370
rect 10682 15314 10750 15370
rect 10806 15314 10874 15370
rect 10930 15314 10998 15370
rect 11054 15314 11122 15370
rect 11178 15314 11246 15370
rect 11302 15314 11370 15370
rect 11426 15314 11494 15370
rect 11550 15314 11618 15370
rect 11674 15314 11742 15370
rect 11798 15314 11866 15370
rect 11922 15314 11990 15370
rect 12046 15314 12114 15370
rect 12170 15314 12180 15370
rect 10244 15246 12180 15314
rect 10244 15190 10254 15246
rect 10310 15190 10378 15246
rect 10434 15190 10502 15246
rect 10558 15190 10626 15246
rect 10682 15190 10750 15246
rect 10806 15190 10874 15246
rect 10930 15190 10998 15246
rect 11054 15190 11122 15246
rect 11178 15190 11246 15246
rect 11302 15190 11370 15246
rect 11426 15190 11494 15246
rect 11550 15190 11618 15246
rect 11674 15190 11742 15246
rect 11798 15190 11866 15246
rect 11922 15190 11990 15246
rect 12046 15190 12114 15246
rect 12170 15190 12180 15246
rect 10244 15122 12180 15190
rect 10244 15066 10254 15122
rect 10310 15066 10378 15122
rect 10434 15066 10502 15122
rect 10558 15066 10626 15122
rect 10682 15066 10750 15122
rect 10806 15066 10874 15122
rect 10930 15066 10998 15122
rect 11054 15066 11122 15122
rect 11178 15066 11246 15122
rect 11302 15066 11370 15122
rect 11426 15066 11494 15122
rect 11550 15066 11618 15122
rect 11674 15066 11742 15122
rect 11798 15066 11866 15122
rect 11922 15066 11990 15122
rect 12046 15066 12114 15122
rect 12170 15066 12180 15122
rect 10244 14998 12180 15066
rect 10244 14942 10254 14998
rect 10310 14942 10378 14998
rect 10434 14942 10502 14998
rect 10558 14942 10626 14998
rect 10682 14942 10750 14998
rect 10806 14942 10874 14998
rect 10930 14942 10998 14998
rect 11054 14942 11122 14998
rect 11178 14942 11246 14998
rect 11302 14942 11370 14998
rect 11426 14942 11494 14998
rect 11550 14942 11618 14998
rect 11674 14942 11742 14998
rect 11798 14942 11866 14998
rect 11922 14942 11990 14998
rect 12046 14942 12114 14998
rect 12170 14942 12180 14998
rect 10244 14874 12180 14942
rect 10244 14818 10254 14874
rect 10310 14818 10378 14874
rect 10434 14818 10502 14874
rect 10558 14818 10626 14874
rect 10682 14818 10750 14874
rect 10806 14818 10874 14874
rect 10930 14818 10998 14874
rect 11054 14818 11122 14874
rect 11178 14818 11246 14874
rect 11302 14818 11370 14874
rect 11426 14818 11494 14874
rect 11550 14818 11618 14874
rect 11674 14818 11742 14874
rect 11798 14818 11866 14874
rect 11922 14818 11990 14874
rect 12046 14818 12114 14874
rect 12170 14818 12180 14874
rect 10244 14750 12180 14818
rect 10244 14694 10254 14750
rect 10310 14694 10378 14750
rect 10434 14694 10502 14750
rect 10558 14694 10626 14750
rect 10682 14694 10750 14750
rect 10806 14694 10874 14750
rect 10930 14694 10998 14750
rect 11054 14694 11122 14750
rect 11178 14694 11246 14750
rect 11302 14694 11370 14750
rect 11426 14694 11494 14750
rect 11550 14694 11618 14750
rect 11674 14694 11742 14750
rect 11798 14694 11866 14750
rect 11922 14694 11990 14750
rect 12046 14694 12114 14750
rect 12170 14694 12180 14750
rect 10244 14626 12180 14694
rect 10244 14570 10254 14626
rect 10310 14570 10378 14626
rect 10434 14570 10502 14626
rect 10558 14570 10626 14626
rect 10682 14570 10750 14626
rect 10806 14570 10874 14626
rect 10930 14570 10998 14626
rect 11054 14570 11122 14626
rect 11178 14570 11246 14626
rect 11302 14570 11370 14626
rect 11426 14570 11494 14626
rect 11550 14570 11618 14626
rect 11674 14570 11742 14626
rect 11798 14570 11866 14626
rect 11922 14570 11990 14626
rect 12046 14570 12114 14626
rect 12170 14570 12180 14626
rect 10244 14502 12180 14570
rect 10244 14446 10254 14502
rect 10310 14446 10378 14502
rect 10434 14446 10502 14502
rect 10558 14446 10626 14502
rect 10682 14446 10750 14502
rect 10806 14446 10874 14502
rect 10930 14446 10998 14502
rect 11054 14446 11122 14502
rect 11178 14446 11246 14502
rect 11302 14446 11370 14502
rect 11426 14446 11494 14502
rect 11550 14446 11618 14502
rect 11674 14446 11742 14502
rect 11798 14446 11866 14502
rect 11922 14446 11990 14502
rect 12046 14446 12114 14502
rect 12170 14446 12180 14502
rect 10244 14436 12180 14446
rect 12861 17354 14673 17364
rect 12861 17298 12871 17354
rect 12927 17298 12995 17354
rect 13051 17298 13119 17354
rect 13175 17298 13243 17354
rect 13299 17298 13367 17354
rect 13423 17298 13491 17354
rect 13547 17298 13615 17354
rect 13671 17298 13739 17354
rect 13795 17298 13863 17354
rect 13919 17298 13987 17354
rect 14043 17298 14111 17354
rect 14167 17298 14235 17354
rect 14291 17298 14359 17354
rect 14415 17298 14483 17354
rect 14539 17298 14607 17354
rect 14663 17298 14673 17354
rect 12861 17230 14673 17298
rect 12861 17174 12871 17230
rect 12927 17174 12995 17230
rect 13051 17174 13119 17230
rect 13175 17174 13243 17230
rect 13299 17174 13367 17230
rect 13423 17174 13491 17230
rect 13547 17174 13615 17230
rect 13671 17174 13739 17230
rect 13795 17174 13863 17230
rect 13919 17174 13987 17230
rect 14043 17174 14111 17230
rect 14167 17174 14235 17230
rect 14291 17174 14359 17230
rect 14415 17174 14483 17230
rect 14539 17174 14607 17230
rect 14663 17174 14673 17230
rect 12861 17106 14673 17174
rect 12861 17050 12871 17106
rect 12927 17050 12995 17106
rect 13051 17050 13119 17106
rect 13175 17050 13243 17106
rect 13299 17050 13367 17106
rect 13423 17050 13491 17106
rect 13547 17050 13615 17106
rect 13671 17050 13739 17106
rect 13795 17050 13863 17106
rect 13919 17050 13987 17106
rect 14043 17050 14111 17106
rect 14167 17050 14235 17106
rect 14291 17050 14359 17106
rect 14415 17050 14483 17106
rect 14539 17050 14607 17106
rect 14663 17050 14673 17106
rect 12861 16982 14673 17050
rect 12861 16926 12871 16982
rect 12927 16926 12995 16982
rect 13051 16926 13119 16982
rect 13175 16926 13243 16982
rect 13299 16926 13367 16982
rect 13423 16926 13491 16982
rect 13547 16926 13615 16982
rect 13671 16926 13739 16982
rect 13795 16926 13863 16982
rect 13919 16926 13987 16982
rect 14043 16926 14111 16982
rect 14167 16926 14235 16982
rect 14291 16926 14359 16982
rect 14415 16926 14483 16982
rect 14539 16926 14607 16982
rect 14663 16926 14673 16982
rect 12861 16858 14673 16926
rect 12861 16802 12871 16858
rect 12927 16802 12995 16858
rect 13051 16802 13119 16858
rect 13175 16802 13243 16858
rect 13299 16802 13367 16858
rect 13423 16802 13491 16858
rect 13547 16802 13615 16858
rect 13671 16802 13739 16858
rect 13795 16802 13863 16858
rect 13919 16802 13987 16858
rect 14043 16802 14111 16858
rect 14167 16802 14235 16858
rect 14291 16802 14359 16858
rect 14415 16802 14483 16858
rect 14539 16802 14607 16858
rect 14663 16802 14673 16858
rect 12861 16734 14673 16802
rect 12861 16678 12871 16734
rect 12927 16678 12995 16734
rect 13051 16678 13119 16734
rect 13175 16678 13243 16734
rect 13299 16678 13367 16734
rect 13423 16678 13491 16734
rect 13547 16678 13615 16734
rect 13671 16678 13739 16734
rect 13795 16678 13863 16734
rect 13919 16678 13987 16734
rect 14043 16678 14111 16734
rect 14167 16678 14235 16734
rect 14291 16678 14359 16734
rect 14415 16678 14483 16734
rect 14539 16678 14607 16734
rect 14663 16678 14673 16734
rect 12861 16610 14673 16678
rect 12861 16554 12871 16610
rect 12927 16554 12995 16610
rect 13051 16554 13119 16610
rect 13175 16554 13243 16610
rect 13299 16554 13367 16610
rect 13423 16554 13491 16610
rect 13547 16554 13615 16610
rect 13671 16554 13739 16610
rect 13795 16554 13863 16610
rect 13919 16554 13987 16610
rect 14043 16554 14111 16610
rect 14167 16554 14235 16610
rect 14291 16554 14359 16610
rect 14415 16554 14483 16610
rect 14539 16554 14607 16610
rect 14663 16554 14673 16610
rect 12861 16486 14673 16554
rect 12861 16430 12871 16486
rect 12927 16430 12995 16486
rect 13051 16430 13119 16486
rect 13175 16430 13243 16486
rect 13299 16430 13367 16486
rect 13423 16430 13491 16486
rect 13547 16430 13615 16486
rect 13671 16430 13739 16486
rect 13795 16430 13863 16486
rect 13919 16430 13987 16486
rect 14043 16430 14111 16486
rect 14167 16430 14235 16486
rect 14291 16430 14359 16486
rect 14415 16430 14483 16486
rect 14539 16430 14607 16486
rect 14663 16430 14673 16486
rect 12861 16362 14673 16430
rect 12861 16306 12871 16362
rect 12927 16306 12995 16362
rect 13051 16306 13119 16362
rect 13175 16306 13243 16362
rect 13299 16306 13367 16362
rect 13423 16306 13491 16362
rect 13547 16306 13615 16362
rect 13671 16306 13739 16362
rect 13795 16306 13863 16362
rect 13919 16306 13987 16362
rect 14043 16306 14111 16362
rect 14167 16306 14235 16362
rect 14291 16306 14359 16362
rect 14415 16306 14483 16362
rect 14539 16306 14607 16362
rect 14663 16306 14673 16362
rect 12861 16238 14673 16306
rect 12861 16182 12871 16238
rect 12927 16182 12995 16238
rect 13051 16182 13119 16238
rect 13175 16182 13243 16238
rect 13299 16182 13367 16238
rect 13423 16182 13491 16238
rect 13547 16182 13615 16238
rect 13671 16182 13739 16238
rect 13795 16182 13863 16238
rect 13919 16182 13987 16238
rect 14043 16182 14111 16238
rect 14167 16182 14235 16238
rect 14291 16182 14359 16238
rect 14415 16182 14483 16238
rect 14539 16182 14607 16238
rect 14663 16182 14673 16238
rect 12861 16114 14673 16182
rect 12861 16058 12871 16114
rect 12927 16058 12995 16114
rect 13051 16058 13119 16114
rect 13175 16058 13243 16114
rect 13299 16058 13367 16114
rect 13423 16058 13491 16114
rect 13547 16058 13615 16114
rect 13671 16058 13739 16114
rect 13795 16058 13863 16114
rect 13919 16058 13987 16114
rect 14043 16058 14111 16114
rect 14167 16058 14235 16114
rect 14291 16058 14359 16114
rect 14415 16058 14483 16114
rect 14539 16058 14607 16114
rect 14663 16058 14673 16114
rect 12861 15990 14673 16058
rect 12861 15934 12871 15990
rect 12927 15934 12995 15990
rect 13051 15934 13119 15990
rect 13175 15934 13243 15990
rect 13299 15934 13367 15990
rect 13423 15934 13491 15990
rect 13547 15934 13615 15990
rect 13671 15934 13739 15990
rect 13795 15934 13863 15990
rect 13919 15934 13987 15990
rect 14043 15934 14111 15990
rect 14167 15934 14235 15990
rect 14291 15934 14359 15990
rect 14415 15934 14483 15990
rect 14539 15934 14607 15990
rect 14663 15934 14673 15990
rect 12861 15866 14673 15934
rect 12861 15810 12871 15866
rect 12927 15810 12995 15866
rect 13051 15810 13119 15866
rect 13175 15810 13243 15866
rect 13299 15810 13367 15866
rect 13423 15810 13491 15866
rect 13547 15810 13615 15866
rect 13671 15810 13739 15866
rect 13795 15810 13863 15866
rect 13919 15810 13987 15866
rect 14043 15810 14111 15866
rect 14167 15810 14235 15866
rect 14291 15810 14359 15866
rect 14415 15810 14483 15866
rect 14539 15810 14607 15866
rect 14663 15810 14673 15866
rect 12861 15742 14673 15810
rect 12861 15686 12871 15742
rect 12927 15686 12995 15742
rect 13051 15686 13119 15742
rect 13175 15686 13243 15742
rect 13299 15686 13367 15742
rect 13423 15686 13491 15742
rect 13547 15686 13615 15742
rect 13671 15686 13739 15742
rect 13795 15686 13863 15742
rect 13919 15686 13987 15742
rect 14043 15686 14111 15742
rect 14167 15686 14235 15742
rect 14291 15686 14359 15742
rect 14415 15686 14483 15742
rect 14539 15686 14607 15742
rect 14663 15686 14673 15742
rect 12861 15618 14673 15686
rect 12861 15562 12871 15618
rect 12927 15562 12995 15618
rect 13051 15562 13119 15618
rect 13175 15562 13243 15618
rect 13299 15562 13367 15618
rect 13423 15562 13491 15618
rect 13547 15562 13615 15618
rect 13671 15562 13739 15618
rect 13795 15562 13863 15618
rect 13919 15562 13987 15618
rect 14043 15562 14111 15618
rect 14167 15562 14235 15618
rect 14291 15562 14359 15618
rect 14415 15562 14483 15618
rect 14539 15562 14607 15618
rect 14663 15562 14673 15618
rect 12861 15494 14673 15562
rect 12861 15438 12871 15494
rect 12927 15438 12995 15494
rect 13051 15438 13119 15494
rect 13175 15438 13243 15494
rect 13299 15438 13367 15494
rect 13423 15438 13491 15494
rect 13547 15438 13615 15494
rect 13671 15438 13739 15494
rect 13795 15438 13863 15494
rect 13919 15438 13987 15494
rect 14043 15438 14111 15494
rect 14167 15438 14235 15494
rect 14291 15438 14359 15494
rect 14415 15438 14483 15494
rect 14539 15438 14607 15494
rect 14663 15438 14673 15494
rect 12861 15370 14673 15438
rect 12861 15314 12871 15370
rect 12927 15314 12995 15370
rect 13051 15314 13119 15370
rect 13175 15314 13243 15370
rect 13299 15314 13367 15370
rect 13423 15314 13491 15370
rect 13547 15314 13615 15370
rect 13671 15314 13739 15370
rect 13795 15314 13863 15370
rect 13919 15314 13987 15370
rect 14043 15314 14111 15370
rect 14167 15314 14235 15370
rect 14291 15314 14359 15370
rect 14415 15314 14483 15370
rect 14539 15314 14607 15370
rect 14663 15314 14673 15370
rect 12861 15246 14673 15314
rect 12861 15190 12871 15246
rect 12927 15190 12995 15246
rect 13051 15190 13119 15246
rect 13175 15190 13243 15246
rect 13299 15190 13367 15246
rect 13423 15190 13491 15246
rect 13547 15190 13615 15246
rect 13671 15190 13739 15246
rect 13795 15190 13863 15246
rect 13919 15190 13987 15246
rect 14043 15190 14111 15246
rect 14167 15190 14235 15246
rect 14291 15190 14359 15246
rect 14415 15190 14483 15246
rect 14539 15190 14607 15246
rect 14663 15190 14673 15246
rect 12861 15122 14673 15190
rect 12861 15066 12871 15122
rect 12927 15066 12995 15122
rect 13051 15066 13119 15122
rect 13175 15066 13243 15122
rect 13299 15066 13367 15122
rect 13423 15066 13491 15122
rect 13547 15066 13615 15122
rect 13671 15066 13739 15122
rect 13795 15066 13863 15122
rect 13919 15066 13987 15122
rect 14043 15066 14111 15122
rect 14167 15066 14235 15122
rect 14291 15066 14359 15122
rect 14415 15066 14483 15122
rect 14539 15066 14607 15122
rect 14663 15066 14673 15122
rect 12861 14998 14673 15066
rect 12861 14942 12871 14998
rect 12927 14942 12995 14998
rect 13051 14942 13119 14998
rect 13175 14942 13243 14998
rect 13299 14942 13367 14998
rect 13423 14942 13491 14998
rect 13547 14942 13615 14998
rect 13671 14942 13739 14998
rect 13795 14942 13863 14998
rect 13919 14942 13987 14998
rect 14043 14942 14111 14998
rect 14167 14942 14235 14998
rect 14291 14942 14359 14998
rect 14415 14942 14483 14998
rect 14539 14942 14607 14998
rect 14663 14942 14673 14998
rect 12861 14874 14673 14942
rect 12861 14818 12871 14874
rect 12927 14818 12995 14874
rect 13051 14818 13119 14874
rect 13175 14818 13243 14874
rect 13299 14818 13367 14874
rect 13423 14818 13491 14874
rect 13547 14818 13615 14874
rect 13671 14818 13739 14874
rect 13795 14818 13863 14874
rect 13919 14818 13987 14874
rect 14043 14818 14111 14874
rect 14167 14818 14235 14874
rect 14291 14818 14359 14874
rect 14415 14818 14483 14874
rect 14539 14818 14607 14874
rect 14663 14818 14673 14874
rect 12861 14750 14673 14818
rect 12861 14694 12871 14750
rect 12927 14694 12995 14750
rect 13051 14694 13119 14750
rect 13175 14694 13243 14750
rect 13299 14694 13367 14750
rect 13423 14694 13491 14750
rect 13547 14694 13615 14750
rect 13671 14694 13739 14750
rect 13795 14694 13863 14750
rect 13919 14694 13987 14750
rect 14043 14694 14111 14750
rect 14167 14694 14235 14750
rect 14291 14694 14359 14750
rect 14415 14694 14483 14750
rect 14539 14694 14607 14750
rect 14663 14694 14673 14750
rect 12861 14626 14673 14694
rect 12861 14570 12871 14626
rect 12927 14570 12995 14626
rect 13051 14570 13119 14626
rect 13175 14570 13243 14626
rect 13299 14570 13367 14626
rect 13423 14570 13491 14626
rect 13547 14570 13615 14626
rect 13671 14570 13739 14626
rect 13795 14570 13863 14626
rect 13919 14570 13987 14626
rect 14043 14570 14111 14626
rect 14167 14570 14235 14626
rect 14291 14570 14359 14626
rect 14415 14570 14483 14626
rect 14539 14570 14607 14626
rect 14663 14570 14673 14626
rect 12861 14502 14673 14570
rect 12861 14446 12871 14502
rect 12927 14446 12995 14502
rect 13051 14446 13119 14502
rect 13175 14446 13243 14502
rect 13299 14446 13367 14502
rect 13423 14446 13491 14502
rect 13547 14446 13615 14502
rect 13671 14446 13739 14502
rect 13795 14446 13863 14502
rect 13919 14446 13987 14502
rect 14043 14446 14111 14502
rect 14167 14446 14235 14502
rect 14291 14446 14359 14502
rect 14415 14446 14483 14502
rect 14539 14446 14607 14502
rect 14663 14446 14673 14502
rect 12861 14436 14673 14446
rect 2481 14148 2681 14158
rect 2481 14092 2491 14148
rect 2547 14092 2615 14148
rect 2671 14092 2681 14148
rect 2481 14024 2681 14092
rect 2481 13968 2491 14024
rect 2547 13968 2615 14024
rect 2671 13968 2681 14024
rect 2481 13900 2681 13968
rect 2481 13844 2491 13900
rect 2547 13844 2615 13900
rect 2671 13844 2681 13900
rect 2481 13776 2681 13844
rect 2481 13720 2491 13776
rect 2547 13720 2615 13776
rect 2671 13720 2681 13776
rect 2481 13652 2681 13720
rect 2481 13596 2491 13652
rect 2547 13596 2615 13652
rect 2671 13596 2681 13652
rect 2481 13528 2681 13596
rect 2481 13472 2491 13528
rect 2547 13472 2615 13528
rect 2671 13472 2681 13528
rect 2481 13404 2681 13472
rect 2481 13348 2491 13404
rect 2547 13348 2615 13404
rect 2671 13348 2681 13404
rect 2481 13280 2681 13348
rect 2481 13224 2491 13280
rect 2547 13224 2615 13280
rect 2671 13224 2681 13280
rect 2481 13156 2681 13224
rect 2481 13100 2491 13156
rect 2547 13100 2615 13156
rect 2671 13100 2681 13156
rect 2481 13032 2681 13100
rect 2481 12976 2491 13032
rect 2547 12976 2615 13032
rect 2671 12976 2681 13032
rect 2481 12908 2681 12976
rect 2481 12852 2491 12908
rect 2547 12852 2615 12908
rect 2671 12852 2681 12908
rect 2481 12842 2681 12852
rect 4851 14148 5051 14158
rect 4851 14092 4861 14148
rect 4917 14092 4985 14148
rect 5041 14092 5051 14148
rect 4851 14024 5051 14092
rect 4851 13968 4861 14024
rect 4917 13968 4985 14024
rect 5041 13968 5051 14024
rect 4851 13900 5051 13968
rect 4851 13844 4861 13900
rect 4917 13844 4985 13900
rect 5041 13844 5051 13900
rect 4851 13776 5051 13844
rect 4851 13720 4861 13776
rect 4917 13720 4985 13776
rect 5041 13720 5051 13776
rect 4851 13652 5051 13720
rect 4851 13596 4861 13652
rect 4917 13596 4985 13652
rect 5041 13596 5051 13652
rect 4851 13528 5051 13596
rect 4851 13472 4861 13528
rect 4917 13472 4985 13528
rect 5041 13472 5051 13528
rect 4851 13404 5051 13472
rect 4851 13348 4861 13404
rect 4917 13348 4985 13404
rect 5041 13348 5051 13404
rect 4851 13280 5051 13348
rect 4851 13224 4861 13280
rect 4917 13224 4985 13280
rect 5041 13224 5051 13280
rect 4851 13156 5051 13224
rect 4851 13100 4861 13156
rect 4917 13100 4985 13156
rect 5041 13100 5051 13156
rect 4851 13032 5051 13100
rect 4851 12976 4861 13032
rect 4917 12976 4985 13032
rect 5041 12976 5051 13032
rect 4851 12908 5051 12976
rect 4851 12852 4861 12908
rect 4917 12852 4985 12908
rect 5041 12852 5051 12908
rect 4851 12842 5051 12852
rect 7265 14148 7713 14158
rect 7265 14092 7275 14148
rect 7331 14092 7399 14148
rect 7455 14092 7523 14148
rect 7579 14092 7647 14148
rect 7703 14092 7713 14148
rect 7265 14024 7713 14092
rect 7265 13968 7275 14024
rect 7331 13968 7399 14024
rect 7455 13968 7523 14024
rect 7579 13968 7647 14024
rect 7703 13968 7713 14024
rect 7265 13900 7713 13968
rect 7265 13844 7275 13900
rect 7331 13844 7399 13900
rect 7455 13844 7523 13900
rect 7579 13844 7647 13900
rect 7703 13844 7713 13900
rect 7265 13776 7713 13844
rect 7265 13720 7275 13776
rect 7331 13720 7399 13776
rect 7455 13720 7523 13776
rect 7579 13720 7647 13776
rect 7703 13720 7713 13776
rect 7265 13652 7713 13720
rect 7265 13596 7275 13652
rect 7331 13596 7399 13652
rect 7455 13596 7523 13652
rect 7579 13596 7647 13652
rect 7703 13596 7713 13652
rect 7265 13528 7713 13596
rect 7265 13472 7275 13528
rect 7331 13472 7399 13528
rect 7455 13472 7523 13528
rect 7579 13472 7647 13528
rect 7703 13472 7713 13528
rect 7265 13404 7713 13472
rect 7265 13348 7275 13404
rect 7331 13348 7399 13404
rect 7455 13348 7523 13404
rect 7579 13348 7647 13404
rect 7703 13348 7713 13404
rect 7265 13280 7713 13348
rect 7265 13224 7275 13280
rect 7331 13224 7399 13280
rect 7455 13224 7523 13280
rect 7579 13224 7647 13280
rect 7703 13224 7713 13280
rect 7265 13156 7713 13224
rect 7265 13100 7275 13156
rect 7331 13100 7399 13156
rect 7455 13100 7523 13156
rect 7579 13100 7647 13156
rect 7703 13100 7713 13156
rect 7265 13032 7713 13100
rect 7265 12976 7275 13032
rect 7331 12976 7399 13032
rect 7455 12976 7523 13032
rect 7579 12976 7647 13032
rect 7703 12976 7713 13032
rect 7265 12908 7713 12976
rect 7265 12852 7275 12908
rect 7331 12852 7399 12908
rect 7455 12852 7523 12908
rect 7579 12852 7647 12908
rect 7703 12852 7713 12908
rect 7265 12842 7713 12852
rect 9927 14148 10127 14158
rect 9927 14092 9937 14148
rect 9993 14092 10061 14148
rect 10117 14092 10127 14148
rect 9927 14024 10127 14092
rect 9927 13968 9937 14024
rect 9993 13968 10061 14024
rect 10117 13968 10127 14024
rect 9927 13900 10127 13968
rect 9927 13844 9937 13900
rect 9993 13844 10061 13900
rect 10117 13844 10127 13900
rect 9927 13776 10127 13844
rect 9927 13720 9937 13776
rect 9993 13720 10061 13776
rect 10117 13720 10127 13776
rect 9927 13652 10127 13720
rect 9927 13596 9937 13652
rect 9993 13596 10061 13652
rect 10117 13596 10127 13652
rect 9927 13528 10127 13596
rect 9927 13472 9937 13528
rect 9993 13472 10061 13528
rect 10117 13472 10127 13528
rect 9927 13404 10127 13472
rect 9927 13348 9937 13404
rect 9993 13348 10061 13404
rect 10117 13348 10127 13404
rect 9927 13280 10127 13348
rect 9927 13224 9937 13280
rect 9993 13224 10061 13280
rect 10117 13224 10127 13280
rect 9927 13156 10127 13224
rect 9927 13100 9937 13156
rect 9993 13100 10061 13156
rect 10117 13100 10127 13156
rect 9927 13032 10127 13100
rect 9927 12976 9937 13032
rect 9993 12976 10061 13032
rect 10117 12976 10127 13032
rect 9927 12908 10127 12976
rect 9927 12852 9937 12908
rect 9993 12852 10061 12908
rect 10117 12852 10127 12908
rect 9927 12842 10127 12852
rect 12297 14148 12497 14158
rect 12297 14092 12307 14148
rect 12363 14092 12431 14148
rect 12487 14092 12497 14148
rect 12297 14024 12497 14092
rect 12297 13968 12307 14024
rect 12363 13968 12431 14024
rect 12487 13968 12497 14024
rect 12297 13900 12497 13968
rect 12297 13844 12307 13900
rect 12363 13844 12431 13900
rect 12487 13844 12497 13900
rect 12297 13776 12497 13844
rect 12297 13720 12307 13776
rect 12363 13720 12431 13776
rect 12487 13720 12497 13776
rect 12297 13652 12497 13720
rect 12297 13596 12307 13652
rect 12363 13596 12431 13652
rect 12487 13596 12497 13652
rect 12297 13528 12497 13596
rect 12297 13472 12307 13528
rect 12363 13472 12431 13528
rect 12487 13472 12497 13528
rect 12297 13404 12497 13472
rect 12297 13348 12307 13404
rect 12363 13348 12431 13404
rect 12487 13348 12497 13404
rect 12297 13280 12497 13348
rect 12297 13224 12307 13280
rect 12363 13224 12431 13280
rect 12487 13224 12497 13280
rect 12297 13156 12497 13224
rect 12297 13100 12307 13156
rect 12363 13100 12431 13156
rect 12487 13100 12497 13156
rect 12297 13032 12497 13100
rect 12297 12976 12307 13032
rect 12363 12976 12431 13032
rect 12487 12976 12497 13032
rect 12297 12908 12497 12976
rect 12297 12852 12307 12908
rect 12363 12852 12431 12908
rect 12487 12852 12497 12908
rect 12297 12842 12497 12852
rect 305 12548 2117 12558
rect 305 12492 315 12548
rect 371 12492 439 12548
rect 495 12492 563 12548
rect 619 12492 687 12548
rect 743 12492 811 12548
rect 867 12492 935 12548
rect 991 12492 1059 12548
rect 1115 12492 1183 12548
rect 1239 12492 1307 12548
rect 1363 12492 1431 12548
rect 1487 12492 1555 12548
rect 1611 12492 1679 12548
rect 1735 12492 1803 12548
rect 1859 12492 1927 12548
rect 1983 12492 2051 12548
rect 2107 12492 2117 12548
rect 305 12424 2117 12492
rect 305 12368 315 12424
rect 371 12368 439 12424
rect 495 12368 563 12424
rect 619 12368 687 12424
rect 743 12368 811 12424
rect 867 12368 935 12424
rect 991 12368 1059 12424
rect 1115 12368 1183 12424
rect 1239 12368 1307 12424
rect 1363 12368 1431 12424
rect 1487 12368 1555 12424
rect 1611 12368 1679 12424
rect 1735 12368 1803 12424
rect 1859 12368 1927 12424
rect 1983 12368 2051 12424
rect 2107 12368 2117 12424
rect 305 12300 2117 12368
rect 305 12244 315 12300
rect 371 12244 439 12300
rect 495 12244 563 12300
rect 619 12244 687 12300
rect 743 12244 811 12300
rect 867 12244 935 12300
rect 991 12244 1059 12300
rect 1115 12244 1183 12300
rect 1239 12244 1307 12300
rect 1363 12244 1431 12300
rect 1487 12244 1555 12300
rect 1611 12244 1679 12300
rect 1735 12244 1803 12300
rect 1859 12244 1927 12300
rect 1983 12244 2051 12300
rect 2107 12244 2117 12300
rect 305 12176 2117 12244
rect 305 12120 315 12176
rect 371 12120 439 12176
rect 495 12120 563 12176
rect 619 12120 687 12176
rect 743 12120 811 12176
rect 867 12120 935 12176
rect 991 12120 1059 12176
rect 1115 12120 1183 12176
rect 1239 12120 1307 12176
rect 1363 12120 1431 12176
rect 1487 12120 1555 12176
rect 1611 12120 1679 12176
rect 1735 12120 1803 12176
rect 1859 12120 1927 12176
rect 1983 12120 2051 12176
rect 2107 12120 2117 12176
rect 305 12052 2117 12120
rect 305 11996 315 12052
rect 371 11996 439 12052
rect 495 11996 563 12052
rect 619 11996 687 12052
rect 743 11996 811 12052
rect 867 11996 935 12052
rect 991 11996 1059 12052
rect 1115 11996 1183 12052
rect 1239 11996 1307 12052
rect 1363 11996 1431 12052
rect 1487 11996 1555 12052
rect 1611 11996 1679 12052
rect 1735 11996 1803 12052
rect 1859 11996 1927 12052
rect 1983 11996 2051 12052
rect 2107 11996 2117 12052
rect 305 11928 2117 11996
rect 305 11872 315 11928
rect 371 11872 439 11928
rect 495 11872 563 11928
rect 619 11872 687 11928
rect 743 11872 811 11928
rect 867 11872 935 11928
rect 991 11872 1059 11928
rect 1115 11872 1183 11928
rect 1239 11872 1307 11928
rect 1363 11872 1431 11928
rect 1487 11872 1555 11928
rect 1611 11872 1679 11928
rect 1735 11872 1803 11928
rect 1859 11872 1927 11928
rect 1983 11872 2051 11928
rect 2107 11872 2117 11928
rect 305 11804 2117 11872
rect 305 11748 315 11804
rect 371 11748 439 11804
rect 495 11748 563 11804
rect 619 11748 687 11804
rect 743 11748 811 11804
rect 867 11748 935 11804
rect 991 11748 1059 11804
rect 1115 11748 1183 11804
rect 1239 11748 1307 11804
rect 1363 11748 1431 11804
rect 1487 11748 1555 11804
rect 1611 11748 1679 11804
rect 1735 11748 1803 11804
rect 1859 11748 1927 11804
rect 1983 11748 2051 11804
rect 2107 11748 2117 11804
rect 305 11680 2117 11748
rect 305 11624 315 11680
rect 371 11624 439 11680
rect 495 11624 563 11680
rect 619 11624 687 11680
rect 743 11624 811 11680
rect 867 11624 935 11680
rect 991 11624 1059 11680
rect 1115 11624 1183 11680
rect 1239 11624 1307 11680
rect 1363 11624 1431 11680
rect 1487 11624 1555 11680
rect 1611 11624 1679 11680
rect 1735 11624 1803 11680
rect 1859 11624 1927 11680
rect 1983 11624 2051 11680
rect 2107 11624 2117 11680
rect 305 11556 2117 11624
rect 305 11500 315 11556
rect 371 11500 439 11556
rect 495 11500 563 11556
rect 619 11500 687 11556
rect 743 11500 811 11556
rect 867 11500 935 11556
rect 991 11500 1059 11556
rect 1115 11500 1183 11556
rect 1239 11500 1307 11556
rect 1363 11500 1431 11556
rect 1487 11500 1555 11556
rect 1611 11500 1679 11556
rect 1735 11500 1803 11556
rect 1859 11500 1927 11556
rect 1983 11500 2051 11556
rect 2107 11500 2117 11556
rect 305 11432 2117 11500
rect 305 11376 315 11432
rect 371 11376 439 11432
rect 495 11376 563 11432
rect 619 11376 687 11432
rect 743 11376 811 11432
rect 867 11376 935 11432
rect 991 11376 1059 11432
rect 1115 11376 1183 11432
rect 1239 11376 1307 11432
rect 1363 11376 1431 11432
rect 1487 11376 1555 11432
rect 1611 11376 1679 11432
rect 1735 11376 1803 11432
rect 1859 11376 1927 11432
rect 1983 11376 2051 11432
rect 2107 11376 2117 11432
rect 305 11308 2117 11376
rect 305 11252 315 11308
rect 371 11252 439 11308
rect 495 11252 563 11308
rect 619 11252 687 11308
rect 743 11252 811 11308
rect 867 11252 935 11308
rect 991 11252 1059 11308
rect 1115 11252 1183 11308
rect 1239 11252 1307 11308
rect 1363 11252 1431 11308
rect 1487 11252 1555 11308
rect 1611 11252 1679 11308
rect 1735 11252 1803 11308
rect 1859 11252 1927 11308
rect 1983 11252 2051 11308
rect 2107 11252 2117 11308
rect 305 11242 2117 11252
rect 2798 12548 4734 12558
rect 2798 12492 2808 12548
rect 2864 12492 2932 12548
rect 2988 12492 3056 12548
rect 3112 12492 3180 12548
rect 3236 12492 3304 12548
rect 3360 12492 3428 12548
rect 3484 12492 3552 12548
rect 3608 12492 3676 12548
rect 3732 12492 3800 12548
rect 3856 12492 3924 12548
rect 3980 12492 4048 12548
rect 4104 12492 4172 12548
rect 4228 12492 4296 12548
rect 4352 12492 4420 12548
rect 4476 12492 4544 12548
rect 4600 12492 4668 12548
rect 4724 12492 4734 12548
rect 2798 12424 4734 12492
rect 2798 12368 2808 12424
rect 2864 12368 2932 12424
rect 2988 12368 3056 12424
rect 3112 12368 3180 12424
rect 3236 12368 3304 12424
rect 3360 12368 3428 12424
rect 3484 12368 3552 12424
rect 3608 12368 3676 12424
rect 3732 12368 3800 12424
rect 3856 12368 3924 12424
rect 3980 12368 4048 12424
rect 4104 12368 4172 12424
rect 4228 12368 4296 12424
rect 4352 12368 4420 12424
rect 4476 12368 4544 12424
rect 4600 12368 4668 12424
rect 4724 12368 4734 12424
rect 2798 12300 4734 12368
rect 2798 12244 2808 12300
rect 2864 12244 2932 12300
rect 2988 12244 3056 12300
rect 3112 12244 3180 12300
rect 3236 12244 3304 12300
rect 3360 12244 3428 12300
rect 3484 12244 3552 12300
rect 3608 12244 3676 12300
rect 3732 12244 3800 12300
rect 3856 12244 3924 12300
rect 3980 12244 4048 12300
rect 4104 12244 4172 12300
rect 4228 12244 4296 12300
rect 4352 12244 4420 12300
rect 4476 12244 4544 12300
rect 4600 12244 4668 12300
rect 4724 12244 4734 12300
rect 2798 12176 4734 12244
rect 2798 12120 2808 12176
rect 2864 12120 2932 12176
rect 2988 12120 3056 12176
rect 3112 12120 3180 12176
rect 3236 12120 3304 12176
rect 3360 12120 3428 12176
rect 3484 12120 3552 12176
rect 3608 12120 3676 12176
rect 3732 12120 3800 12176
rect 3856 12120 3924 12176
rect 3980 12120 4048 12176
rect 4104 12120 4172 12176
rect 4228 12120 4296 12176
rect 4352 12120 4420 12176
rect 4476 12120 4544 12176
rect 4600 12120 4668 12176
rect 4724 12120 4734 12176
rect 2798 12052 4734 12120
rect 2798 11996 2808 12052
rect 2864 11996 2932 12052
rect 2988 11996 3056 12052
rect 3112 11996 3180 12052
rect 3236 11996 3304 12052
rect 3360 11996 3428 12052
rect 3484 11996 3552 12052
rect 3608 11996 3676 12052
rect 3732 11996 3800 12052
rect 3856 11996 3924 12052
rect 3980 11996 4048 12052
rect 4104 11996 4172 12052
rect 4228 11996 4296 12052
rect 4352 11996 4420 12052
rect 4476 11996 4544 12052
rect 4600 11996 4668 12052
rect 4724 11996 4734 12052
rect 2798 11928 4734 11996
rect 2798 11872 2808 11928
rect 2864 11872 2932 11928
rect 2988 11872 3056 11928
rect 3112 11872 3180 11928
rect 3236 11872 3304 11928
rect 3360 11872 3428 11928
rect 3484 11872 3552 11928
rect 3608 11872 3676 11928
rect 3732 11872 3800 11928
rect 3856 11872 3924 11928
rect 3980 11872 4048 11928
rect 4104 11872 4172 11928
rect 4228 11872 4296 11928
rect 4352 11872 4420 11928
rect 4476 11872 4544 11928
rect 4600 11872 4668 11928
rect 4724 11872 4734 11928
rect 2798 11804 4734 11872
rect 2798 11748 2808 11804
rect 2864 11748 2932 11804
rect 2988 11748 3056 11804
rect 3112 11748 3180 11804
rect 3236 11748 3304 11804
rect 3360 11748 3428 11804
rect 3484 11748 3552 11804
rect 3608 11748 3676 11804
rect 3732 11748 3800 11804
rect 3856 11748 3924 11804
rect 3980 11748 4048 11804
rect 4104 11748 4172 11804
rect 4228 11748 4296 11804
rect 4352 11748 4420 11804
rect 4476 11748 4544 11804
rect 4600 11748 4668 11804
rect 4724 11748 4734 11804
rect 2798 11680 4734 11748
rect 2798 11624 2808 11680
rect 2864 11624 2932 11680
rect 2988 11624 3056 11680
rect 3112 11624 3180 11680
rect 3236 11624 3304 11680
rect 3360 11624 3428 11680
rect 3484 11624 3552 11680
rect 3608 11624 3676 11680
rect 3732 11624 3800 11680
rect 3856 11624 3924 11680
rect 3980 11624 4048 11680
rect 4104 11624 4172 11680
rect 4228 11624 4296 11680
rect 4352 11624 4420 11680
rect 4476 11624 4544 11680
rect 4600 11624 4668 11680
rect 4724 11624 4734 11680
rect 2798 11556 4734 11624
rect 2798 11500 2808 11556
rect 2864 11500 2932 11556
rect 2988 11500 3056 11556
rect 3112 11500 3180 11556
rect 3236 11500 3304 11556
rect 3360 11500 3428 11556
rect 3484 11500 3552 11556
rect 3608 11500 3676 11556
rect 3732 11500 3800 11556
rect 3856 11500 3924 11556
rect 3980 11500 4048 11556
rect 4104 11500 4172 11556
rect 4228 11500 4296 11556
rect 4352 11500 4420 11556
rect 4476 11500 4544 11556
rect 4600 11500 4668 11556
rect 4724 11500 4734 11556
rect 2798 11432 4734 11500
rect 2798 11376 2808 11432
rect 2864 11376 2932 11432
rect 2988 11376 3056 11432
rect 3112 11376 3180 11432
rect 3236 11376 3304 11432
rect 3360 11376 3428 11432
rect 3484 11376 3552 11432
rect 3608 11376 3676 11432
rect 3732 11376 3800 11432
rect 3856 11376 3924 11432
rect 3980 11376 4048 11432
rect 4104 11376 4172 11432
rect 4228 11376 4296 11432
rect 4352 11376 4420 11432
rect 4476 11376 4544 11432
rect 4600 11376 4668 11432
rect 4724 11376 4734 11432
rect 2798 11308 4734 11376
rect 2798 11252 2808 11308
rect 2864 11252 2932 11308
rect 2988 11252 3056 11308
rect 3112 11252 3180 11308
rect 3236 11252 3304 11308
rect 3360 11252 3428 11308
rect 3484 11252 3552 11308
rect 3608 11252 3676 11308
rect 3732 11252 3800 11308
rect 3856 11252 3924 11308
rect 3980 11252 4048 11308
rect 4104 11252 4172 11308
rect 4228 11252 4296 11308
rect 4352 11252 4420 11308
rect 4476 11252 4544 11308
rect 4600 11252 4668 11308
rect 4724 11252 4734 11308
rect 2798 11242 4734 11252
rect 5168 12548 7104 12558
rect 5168 12492 5178 12548
rect 5234 12492 5302 12548
rect 5358 12492 5426 12548
rect 5482 12492 5550 12548
rect 5606 12492 5674 12548
rect 5730 12492 5798 12548
rect 5854 12492 5922 12548
rect 5978 12492 6046 12548
rect 6102 12492 6170 12548
rect 6226 12492 6294 12548
rect 6350 12492 6418 12548
rect 6474 12492 6542 12548
rect 6598 12492 6666 12548
rect 6722 12492 6790 12548
rect 6846 12492 6914 12548
rect 6970 12492 7038 12548
rect 7094 12492 7104 12548
rect 5168 12424 7104 12492
rect 5168 12368 5178 12424
rect 5234 12368 5302 12424
rect 5358 12368 5426 12424
rect 5482 12368 5550 12424
rect 5606 12368 5674 12424
rect 5730 12368 5798 12424
rect 5854 12368 5922 12424
rect 5978 12368 6046 12424
rect 6102 12368 6170 12424
rect 6226 12368 6294 12424
rect 6350 12368 6418 12424
rect 6474 12368 6542 12424
rect 6598 12368 6666 12424
rect 6722 12368 6790 12424
rect 6846 12368 6914 12424
rect 6970 12368 7038 12424
rect 7094 12368 7104 12424
rect 5168 12300 7104 12368
rect 5168 12244 5178 12300
rect 5234 12244 5302 12300
rect 5358 12244 5426 12300
rect 5482 12244 5550 12300
rect 5606 12244 5674 12300
rect 5730 12244 5798 12300
rect 5854 12244 5922 12300
rect 5978 12244 6046 12300
rect 6102 12244 6170 12300
rect 6226 12244 6294 12300
rect 6350 12244 6418 12300
rect 6474 12244 6542 12300
rect 6598 12244 6666 12300
rect 6722 12244 6790 12300
rect 6846 12244 6914 12300
rect 6970 12244 7038 12300
rect 7094 12244 7104 12300
rect 5168 12176 7104 12244
rect 5168 12120 5178 12176
rect 5234 12120 5302 12176
rect 5358 12120 5426 12176
rect 5482 12120 5550 12176
rect 5606 12120 5674 12176
rect 5730 12120 5798 12176
rect 5854 12120 5922 12176
rect 5978 12120 6046 12176
rect 6102 12120 6170 12176
rect 6226 12120 6294 12176
rect 6350 12120 6418 12176
rect 6474 12120 6542 12176
rect 6598 12120 6666 12176
rect 6722 12120 6790 12176
rect 6846 12120 6914 12176
rect 6970 12120 7038 12176
rect 7094 12120 7104 12176
rect 5168 12052 7104 12120
rect 5168 11996 5178 12052
rect 5234 11996 5302 12052
rect 5358 11996 5426 12052
rect 5482 11996 5550 12052
rect 5606 11996 5674 12052
rect 5730 11996 5798 12052
rect 5854 11996 5922 12052
rect 5978 11996 6046 12052
rect 6102 11996 6170 12052
rect 6226 11996 6294 12052
rect 6350 11996 6418 12052
rect 6474 11996 6542 12052
rect 6598 11996 6666 12052
rect 6722 11996 6790 12052
rect 6846 11996 6914 12052
rect 6970 11996 7038 12052
rect 7094 11996 7104 12052
rect 5168 11928 7104 11996
rect 5168 11872 5178 11928
rect 5234 11872 5302 11928
rect 5358 11872 5426 11928
rect 5482 11872 5550 11928
rect 5606 11872 5674 11928
rect 5730 11872 5798 11928
rect 5854 11872 5922 11928
rect 5978 11872 6046 11928
rect 6102 11872 6170 11928
rect 6226 11872 6294 11928
rect 6350 11872 6418 11928
rect 6474 11872 6542 11928
rect 6598 11872 6666 11928
rect 6722 11872 6790 11928
rect 6846 11872 6914 11928
rect 6970 11872 7038 11928
rect 7094 11872 7104 11928
rect 5168 11804 7104 11872
rect 5168 11748 5178 11804
rect 5234 11748 5302 11804
rect 5358 11748 5426 11804
rect 5482 11748 5550 11804
rect 5606 11748 5674 11804
rect 5730 11748 5798 11804
rect 5854 11748 5922 11804
rect 5978 11748 6046 11804
rect 6102 11748 6170 11804
rect 6226 11748 6294 11804
rect 6350 11748 6418 11804
rect 6474 11748 6542 11804
rect 6598 11748 6666 11804
rect 6722 11748 6790 11804
rect 6846 11748 6914 11804
rect 6970 11748 7038 11804
rect 7094 11748 7104 11804
rect 5168 11680 7104 11748
rect 5168 11624 5178 11680
rect 5234 11624 5302 11680
rect 5358 11624 5426 11680
rect 5482 11624 5550 11680
rect 5606 11624 5674 11680
rect 5730 11624 5798 11680
rect 5854 11624 5922 11680
rect 5978 11624 6046 11680
rect 6102 11624 6170 11680
rect 6226 11624 6294 11680
rect 6350 11624 6418 11680
rect 6474 11624 6542 11680
rect 6598 11624 6666 11680
rect 6722 11624 6790 11680
rect 6846 11624 6914 11680
rect 6970 11624 7038 11680
rect 7094 11624 7104 11680
rect 5168 11556 7104 11624
rect 5168 11500 5178 11556
rect 5234 11500 5302 11556
rect 5358 11500 5426 11556
rect 5482 11500 5550 11556
rect 5606 11500 5674 11556
rect 5730 11500 5798 11556
rect 5854 11500 5922 11556
rect 5978 11500 6046 11556
rect 6102 11500 6170 11556
rect 6226 11500 6294 11556
rect 6350 11500 6418 11556
rect 6474 11500 6542 11556
rect 6598 11500 6666 11556
rect 6722 11500 6790 11556
rect 6846 11500 6914 11556
rect 6970 11500 7038 11556
rect 7094 11500 7104 11556
rect 5168 11432 7104 11500
rect 5168 11376 5178 11432
rect 5234 11376 5302 11432
rect 5358 11376 5426 11432
rect 5482 11376 5550 11432
rect 5606 11376 5674 11432
rect 5730 11376 5798 11432
rect 5854 11376 5922 11432
rect 5978 11376 6046 11432
rect 6102 11376 6170 11432
rect 6226 11376 6294 11432
rect 6350 11376 6418 11432
rect 6474 11376 6542 11432
rect 6598 11376 6666 11432
rect 6722 11376 6790 11432
rect 6846 11376 6914 11432
rect 6970 11376 7038 11432
rect 7094 11376 7104 11432
rect 5168 11308 7104 11376
rect 5168 11252 5178 11308
rect 5234 11252 5302 11308
rect 5358 11252 5426 11308
rect 5482 11252 5550 11308
rect 5606 11252 5674 11308
rect 5730 11252 5798 11308
rect 5854 11252 5922 11308
rect 5978 11252 6046 11308
rect 6102 11252 6170 11308
rect 6226 11252 6294 11308
rect 6350 11252 6418 11308
rect 6474 11252 6542 11308
rect 6598 11252 6666 11308
rect 6722 11252 6790 11308
rect 6846 11252 6914 11308
rect 6970 11252 7038 11308
rect 7094 11252 7104 11308
rect 5168 11242 7104 11252
rect 7874 12548 9810 12558
rect 7874 12492 7884 12548
rect 7940 12492 8008 12548
rect 8064 12492 8132 12548
rect 8188 12492 8256 12548
rect 8312 12492 8380 12548
rect 8436 12492 8504 12548
rect 8560 12492 8628 12548
rect 8684 12492 8752 12548
rect 8808 12492 8876 12548
rect 8932 12492 9000 12548
rect 9056 12492 9124 12548
rect 9180 12492 9248 12548
rect 9304 12492 9372 12548
rect 9428 12492 9496 12548
rect 9552 12492 9620 12548
rect 9676 12492 9744 12548
rect 9800 12492 9810 12548
rect 7874 12424 9810 12492
rect 7874 12368 7884 12424
rect 7940 12368 8008 12424
rect 8064 12368 8132 12424
rect 8188 12368 8256 12424
rect 8312 12368 8380 12424
rect 8436 12368 8504 12424
rect 8560 12368 8628 12424
rect 8684 12368 8752 12424
rect 8808 12368 8876 12424
rect 8932 12368 9000 12424
rect 9056 12368 9124 12424
rect 9180 12368 9248 12424
rect 9304 12368 9372 12424
rect 9428 12368 9496 12424
rect 9552 12368 9620 12424
rect 9676 12368 9744 12424
rect 9800 12368 9810 12424
rect 7874 12300 9810 12368
rect 7874 12244 7884 12300
rect 7940 12244 8008 12300
rect 8064 12244 8132 12300
rect 8188 12244 8256 12300
rect 8312 12244 8380 12300
rect 8436 12244 8504 12300
rect 8560 12244 8628 12300
rect 8684 12244 8752 12300
rect 8808 12244 8876 12300
rect 8932 12244 9000 12300
rect 9056 12244 9124 12300
rect 9180 12244 9248 12300
rect 9304 12244 9372 12300
rect 9428 12244 9496 12300
rect 9552 12244 9620 12300
rect 9676 12244 9744 12300
rect 9800 12244 9810 12300
rect 7874 12176 9810 12244
rect 7874 12120 7884 12176
rect 7940 12120 8008 12176
rect 8064 12120 8132 12176
rect 8188 12120 8256 12176
rect 8312 12120 8380 12176
rect 8436 12120 8504 12176
rect 8560 12120 8628 12176
rect 8684 12120 8752 12176
rect 8808 12120 8876 12176
rect 8932 12120 9000 12176
rect 9056 12120 9124 12176
rect 9180 12120 9248 12176
rect 9304 12120 9372 12176
rect 9428 12120 9496 12176
rect 9552 12120 9620 12176
rect 9676 12120 9744 12176
rect 9800 12120 9810 12176
rect 7874 12052 9810 12120
rect 7874 11996 7884 12052
rect 7940 11996 8008 12052
rect 8064 11996 8132 12052
rect 8188 11996 8256 12052
rect 8312 11996 8380 12052
rect 8436 11996 8504 12052
rect 8560 11996 8628 12052
rect 8684 11996 8752 12052
rect 8808 11996 8876 12052
rect 8932 11996 9000 12052
rect 9056 11996 9124 12052
rect 9180 11996 9248 12052
rect 9304 11996 9372 12052
rect 9428 11996 9496 12052
rect 9552 11996 9620 12052
rect 9676 11996 9744 12052
rect 9800 11996 9810 12052
rect 7874 11928 9810 11996
rect 7874 11872 7884 11928
rect 7940 11872 8008 11928
rect 8064 11872 8132 11928
rect 8188 11872 8256 11928
rect 8312 11872 8380 11928
rect 8436 11872 8504 11928
rect 8560 11872 8628 11928
rect 8684 11872 8752 11928
rect 8808 11872 8876 11928
rect 8932 11872 9000 11928
rect 9056 11872 9124 11928
rect 9180 11872 9248 11928
rect 9304 11872 9372 11928
rect 9428 11872 9496 11928
rect 9552 11872 9620 11928
rect 9676 11872 9744 11928
rect 9800 11872 9810 11928
rect 7874 11804 9810 11872
rect 7874 11748 7884 11804
rect 7940 11748 8008 11804
rect 8064 11748 8132 11804
rect 8188 11748 8256 11804
rect 8312 11748 8380 11804
rect 8436 11748 8504 11804
rect 8560 11748 8628 11804
rect 8684 11748 8752 11804
rect 8808 11748 8876 11804
rect 8932 11748 9000 11804
rect 9056 11748 9124 11804
rect 9180 11748 9248 11804
rect 9304 11748 9372 11804
rect 9428 11748 9496 11804
rect 9552 11748 9620 11804
rect 9676 11748 9744 11804
rect 9800 11748 9810 11804
rect 7874 11680 9810 11748
rect 7874 11624 7884 11680
rect 7940 11624 8008 11680
rect 8064 11624 8132 11680
rect 8188 11624 8256 11680
rect 8312 11624 8380 11680
rect 8436 11624 8504 11680
rect 8560 11624 8628 11680
rect 8684 11624 8752 11680
rect 8808 11624 8876 11680
rect 8932 11624 9000 11680
rect 9056 11624 9124 11680
rect 9180 11624 9248 11680
rect 9304 11624 9372 11680
rect 9428 11624 9496 11680
rect 9552 11624 9620 11680
rect 9676 11624 9744 11680
rect 9800 11624 9810 11680
rect 7874 11556 9810 11624
rect 7874 11500 7884 11556
rect 7940 11500 8008 11556
rect 8064 11500 8132 11556
rect 8188 11500 8256 11556
rect 8312 11500 8380 11556
rect 8436 11500 8504 11556
rect 8560 11500 8628 11556
rect 8684 11500 8752 11556
rect 8808 11500 8876 11556
rect 8932 11500 9000 11556
rect 9056 11500 9124 11556
rect 9180 11500 9248 11556
rect 9304 11500 9372 11556
rect 9428 11500 9496 11556
rect 9552 11500 9620 11556
rect 9676 11500 9744 11556
rect 9800 11500 9810 11556
rect 7874 11432 9810 11500
rect 7874 11376 7884 11432
rect 7940 11376 8008 11432
rect 8064 11376 8132 11432
rect 8188 11376 8256 11432
rect 8312 11376 8380 11432
rect 8436 11376 8504 11432
rect 8560 11376 8628 11432
rect 8684 11376 8752 11432
rect 8808 11376 8876 11432
rect 8932 11376 9000 11432
rect 9056 11376 9124 11432
rect 9180 11376 9248 11432
rect 9304 11376 9372 11432
rect 9428 11376 9496 11432
rect 9552 11376 9620 11432
rect 9676 11376 9744 11432
rect 9800 11376 9810 11432
rect 7874 11308 9810 11376
rect 7874 11252 7884 11308
rect 7940 11252 8008 11308
rect 8064 11252 8132 11308
rect 8188 11252 8256 11308
rect 8312 11252 8380 11308
rect 8436 11252 8504 11308
rect 8560 11252 8628 11308
rect 8684 11252 8752 11308
rect 8808 11252 8876 11308
rect 8932 11252 9000 11308
rect 9056 11252 9124 11308
rect 9180 11252 9248 11308
rect 9304 11252 9372 11308
rect 9428 11252 9496 11308
rect 9552 11252 9620 11308
rect 9676 11252 9744 11308
rect 9800 11252 9810 11308
rect 7874 11242 9810 11252
rect 10244 12548 12180 12558
rect 10244 12492 10254 12548
rect 10310 12492 10378 12548
rect 10434 12492 10502 12548
rect 10558 12492 10626 12548
rect 10682 12492 10750 12548
rect 10806 12492 10874 12548
rect 10930 12492 10998 12548
rect 11054 12492 11122 12548
rect 11178 12492 11246 12548
rect 11302 12492 11370 12548
rect 11426 12492 11494 12548
rect 11550 12492 11618 12548
rect 11674 12492 11742 12548
rect 11798 12492 11866 12548
rect 11922 12492 11990 12548
rect 12046 12492 12114 12548
rect 12170 12492 12180 12548
rect 10244 12424 12180 12492
rect 10244 12368 10254 12424
rect 10310 12368 10378 12424
rect 10434 12368 10502 12424
rect 10558 12368 10626 12424
rect 10682 12368 10750 12424
rect 10806 12368 10874 12424
rect 10930 12368 10998 12424
rect 11054 12368 11122 12424
rect 11178 12368 11246 12424
rect 11302 12368 11370 12424
rect 11426 12368 11494 12424
rect 11550 12368 11618 12424
rect 11674 12368 11742 12424
rect 11798 12368 11866 12424
rect 11922 12368 11990 12424
rect 12046 12368 12114 12424
rect 12170 12368 12180 12424
rect 10244 12300 12180 12368
rect 10244 12244 10254 12300
rect 10310 12244 10378 12300
rect 10434 12244 10502 12300
rect 10558 12244 10626 12300
rect 10682 12244 10750 12300
rect 10806 12244 10874 12300
rect 10930 12244 10998 12300
rect 11054 12244 11122 12300
rect 11178 12244 11246 12300
rect 11302 12244 11370 12300
rect 11426 12244 11494 12300
rect 11550 12244 11618 12300
rect 11674 12244 11742 12300
rect 11798 12244 11866 12300
rect 11922 12244 11990 12300
rect 12046 12244 12114 12300
rect 12170 12244 12180 12300
rect 10244 12176 12180 12244
rect 10244 12120 10254 12176
rect 10310 12120 10378 12176
rect 10434 12120 10502 12176
rect 10558 12120 10626 12176
rect 10682 12120 10750 12176
rect 10806 12120 10874 12176
rect 10930 12120 10998 12176
rect 11054 12120 11122 12176
rect 11178 12120 11246 12176
rect 11302 12120 11370 12176
rect 11426 12120 11494 12176
rect 11550 12120 11618 12176
rect 11674 12120 11742 12176
rect 11798 12120 11866 12176
rect 11922 12120 11990 12176
rect 12046 12120 12114 12176
rect 12170 12120 12180 12176
rect 10244 12052 12180 12120
rect 10244 11996 10254 12052
rect 10310 11996 10378 12052
rect 10434 11996 10502 12052
rect 10558 11996 10626 12052
rect 10682 11996 10750 12052
rect 10806 11996 10874 12052
rect 10930 11996 10998 12052
rect 11054 11996 11122 12052
rect 11178 11996 11246 12052
rect 11302 11996 11370 12052
rect 11426 11996 11494 12052
rect 11550 11996 11618 12052
rect 11674 11996 11742 12052
rect 11798 11996 11866 12052
rect 11922 11996 11990 12052
rect 12046 11996 12114 12052
rect 12170 11996 12180 12052
rect 10244 11928 12180 11996
rect 10244 11872 10254 11928
rect 10310 11872 10378 11928
rect 10434 11872 10502 11928
rect 10558 11872 10626 11928
rect 10682 11872 10750 11928
rect 10806 11872 10874 11928
rect 10930 11872 10998 11928
rect 11054 11872 11122 11928
rect 11178 11872 11246 11928
rect 11302 11872 11370 11928
rect 11426 11872 11494 11928
rect 11550 11872 11618 11928
rect 11674 11872 11742 11928
rect 11798 11872 11866 11928
rect 11922 11872 11990 11928
rect 12046 11872 12114 11928
rect 12170 11872 12180 11928
rect 10244 11804 12180 11872
rect 10244 11748 10254 11804
rect 10310 11748 10378 11804
rect 10434 11748 10502 11804
rect 10558 11748 10626 11804
rect 10682 11748 10750 11804
rect 10806 11748 10874 11804
rect 10930 11748 10998 11804
rect 11054 11748 11122 11804
rect 11178 11748 11246 11804
rect 11302 11748 11370 11804
rect 11426 11748 11494 11804
rect 11550 11748 11618 11804
rect 11674 11748 11742 11804
rect 11798 11748 11866 11804
rect 11922 11748 11990 11804
rect 12046 11748 12114 11804
rect 12170 11748 12180 11804
rect 10244 11680 12180 11748
rect 10244 11624 10254 11680
rect 10310 11624 10378 11680
rect 10434 11624 10502 11680
rect 10558 11624 10626 11680
rect 10682 11624 10750 11680
rect 10806 11624 10874 11680
rect 10930 11624 10998 11680
rect 11054 11624 11122 11680
rect 11178 11624 11246 11680
rect 11302 11624 11370 11680
rect 11426 11624 11494 11680
rect 11550 11624 11618 11680
rect 11674 11624 11742 11680
rect 11798 11624 11866 11680
rect 11922 11624 11990 11680
rect 12046 11624 12114 11680
rect 12170 11624 12180 11680
rect 10244 11556 12180 11624
rect 10244 11500 10254 11556
rect 10310 11500 10378 11556
rect 10434 11500 10502 11556
rect 10558 11500 10626 11556
rect 10682 11500 10750 11556
rect 10806 11500 10874 11556
rect 10930 11500 10998 11556
rect 11054 11500 11122 11556
rect 11178 11500 11246 11556
rect 11302 11500 11370 11556
rect 11426 11500 11494 11556
rect 11550 11500 11618 11556
rect 11674 11500 11742 11556
rect 11798 11500 11866 11556
rect 11922 11500 11990 11556
rect 12046 11500 12114 11556
rect 12170 11500 12180 11556
rect 10244 11432 12180 11500
rect 10244 11376 10254 11432
rect 10310 11376 10378 11432
rect 10434 11376 10502 11432
rect 10558 11376 10626 11432
rect 10682 11376 10750 11432
rect 10806 11376 10874 11432
rect 10930 11376 10998 11432
rect 11054 11376 11122 11432
rect 11178 11376 11246 11432
rect 11302 11376 11370 11432
rect 11426 11376 11494 11432
rect 11550 11376 11618 11432
rect 11674 11376 11742 11432
rect 11798 11376 11866 11432
rect 11922 11376 11990 11432
rect 12046 11376 12114 11432
rect 12170 11376 12180 11432
rect 10244 11308 12180 11376
rect 10244 11252 10254 11308
rect 10310 11252 10378 11308
rect 10434 11252 10502 11308
rect 10558 11252 10626 11308
rect 10682 11252 10750 11308
rect 10806 11252 10874 11308
rect 10930 11252 10998 11308
rect 11054 11252 11122 11308
rect 11178 11252 11246 11308
rect 11302 11252 11370 11308
rect 11426 11252 11494 11308
rect 11550 11252 11618 11308
rect 11674 11252 11742 11308
rect 11798 11252 11866 11308
rect 11922 11252 11990 11308
rect 12046 11252 12114 11308
rect 12170 11252 12180 11308
rect 10244 11242 12180 11252
rect 12861 12548 14673 12558
rect 12861 12492 12871 12548
rect 12927 12492 12995 12548
rect 13051 12492 13119 12548
rect 13175 12492 13243 12548
rect 13299 12492 13367 12548
rect 13423 12492 13491 12548
rect 13547 12492 13615 12548
rect 13671 12492 13739 12548
rect 13795 12492 13863 12548
rect 13919 12492 13987 12548
rect 14043 12492 14111 12548
rect 14167 12492 14235 12548
rect 14291 12492 14359 12548
rect 14415 12492 14483 12548
rect 14539 12492 14607 12548
rect 14663 12492 14673 12548
rect 12861 12424 14673 12492
rect 12861 12368 12871 12424
rect 12927 12368 12995 12424
rect 13051 12368 13119 12424
rect 13175 12368 13243 12424
rect 13299 12368 13367 12424
rect 13423 12368 13491 12424
rect 13547 12368 13615 12424
rect 13671 12368 13739 12424
rect 13795 12368 13863 12424
rect 13919 12368 13987 12424
rect 14043 12368 14111 12424
rect 14167 12368 14235 12424
rect 14291 12368 14359 12424
rect 14415 12368 14483 12424
rect 14539 12368 14607 12424
rect 14663 12368 14673 12424
rect 12861 12300 14673 12368
rect 12861 12244 12871 12300
rect 12927 12244 12995 12300
rect 13051 12244 13119 12300
rect 13175 12244 13243 12300
rect 13299 12244 13367 12300
rect 13423 12244 13491 12300
rect 13547 12244 13615 12300
rect 13671 12244 13739 12300
rect 13795 12244 13863 12300
rect 13919 12244 13987 12300
rect 14043 12244 14111 12300
rect 14167 12244 14235 12300
rect 14291 12244 14359 12300
rect 14415 12244 14483 12300
rect 14539 12244 14607 12300
rect 14663 12244 14673 12300
rect 12861 12176 14673 12244
rect 12861 12120 12871 12176
rect 12927 12120 12995 12176
rect 13051 12120 13119 12176
rect 13175 12120 13243 12176
rect 13299 12120 13367 12176
rect 13423 12120 13491 12176
rect 13547 12120 13615 12176
rect 13671 12120 13739 12176
rect 13795 12120 13863 12176
rect 13919 12120 13987 12176
rect 14043 12120 14111 12176
rect 14167 12120 14235 12176
rect 14291 12120 14359 12176
rect 14415 12120 14483 12176
rect 14539 12120 14607 12176
rect 14663 12120 14673 12176
rect 12861 12052 14673 12120
rect 12861 11996 12871 12052
rect 12927 11996 12995 12052
rect 13051 11996 13119 12052
rect 13175 11996 13243 12052
rect 13299 11996 13367 12052
rect 13423 11996 13491 12052
rect 13547 11996 13615 12052
rect 13671 11996 13739 12052
rect 13795 11996 13863 12052
rect 13919 11996 13987 12052
rect 14043 11996 14111 12052
rect 14167 11996 14235 12052
rect 14291 11996 14359 12052
rect 14415 11996 14483 12052
rect 14539 11996 14607 12052
rect 14663 11996 14673 12052
rect 12861 11928 14673 11996
rect 12861 11872 12871 11928
rect 12927 11872 12995 11928
rect 13051 11872 13119 11928
rect 13175 11872 13243 11928
rect 13299 11872 13367 11928
rect 13423 11872 13491 11928
rect 13547 11872 13615 11928
rect 13671 11872 13739 11928
rect 13795 11872 13863 11928
rect 13919 11872 13987 11928
rect 14043 11872 14111 11928
rect 14167 11872 14235 11928
rect 14291 11872 14359 11928
rect 14415 11872 14483 11928
rect 14539 11872 14607 11928
rect 14663 11872 14673 11928
rect 12861 11804 14673 11872
rect 12861 11748 12871 11804
rect 12927 11748 12995 11804
rect 13051 11748 13119 11804
rect 13175 11748 13243 11804
rect 13299 11748 13367 11804
rect 13423 11748 13491 11804
rect 13547 11748 13615 11804
rect 13671 11748 13739 11804
rect 13795 11748 13863 11804
rect 13919 11748 13987 11804
rect 14043 11748 14111 11804
rect 14167 11748 14235 11804
rect 14291 11748 14359 11804
rect 14415 11748 14483 11804
rect 14539 11748 14607 11804
rect 14663 11748 14673 11804
rect 12861 11680 14673 11748
rect 12861 11624 12871 11680
rect 12927 11624 12995 11680
rect 13051 11624 13119 11680
rect 13175 11624 13243 11680
rect 13299 11624 13367 11680
rect 13423 11624 13491 11680
rect 13547 11624 13615 11680
rect 13671 11624 13739 11680
rect 13795 11624 13863 11680
rect 13919 11624 13987 11680
rect 14043 11624 14111 11680
rect 14167 11624 14235 11680
rect 14291 11624 14359 11680
rect 14415 11624 14483 11680
rect 14539 11624 14607 11680
rect 14663 11624 14673 11680
rect 12861 11556 14673 11624
rect 12861 11500 12871 11556
rect 12927 11500 12995 11556
rect 13051 11500 13119 11556
rect 13175 11500 13243 11556
rect 13299 11500 13367 11556
rect 13423 11500 13491 11556
rect 13547 11500 13615 11556
rect 13671 11500 13739 11556
rect 13795 11500 13863 11556
rect 13919 11500 13987 11556
rect 14043 11500 14111 11556
rect 14167 11500 14235 11556
rect 14291 11500 14359 11556
rect 14415 11500 14483 11556
rect 14539 11500 14607 11556
rect 14663 11500 14673 11556
rect 12861 11432 14673 11500
rect 12861 11376 12871 11432
rect 12927 11376 12995 11432
rect 13051 11376 13119 11432
rect 13175 11376 13243 11432
rect 13299 11376 13367 11432
rect 13423 11376 13491 11432
rect 13547 11376 13615 11432
rect 13671 11376 13739 11432
rect 13795 11376 13863 11432
rect 13919 11376 13987 11432
rect 14043 11376 14111 11432
rect 14167 11376 14235 11432
rect 14291 11376 14359 11432
rect 14415 11376 14483 11432
rect 14539 11376 14607 11432
rect 14663 11376 14673 11432
rect 12861 11308 14673 11376
rect 12861 11252 12871 11308
rect 12927 11252 12995 11308
rect 13051 11252 13119 11308
rect 13175 11252 13243 11308
rect 13299 11252 13367 11308
rect 13423 11252 13491 11308
rect 13547 11252 13615 11308
rect 13671 11252 13739 11308
rect 13795 11252 13863 11308
rect 13919 11252 13987 11308
rect 14043 11252 14111 11308
rect 14167 11252 14235 11308
rect 14291 11252 14359 11308
rect 14415 11252 14483 11308
rect 14539 11252 14607 11308
rect 14663 11252 14673 11308
rect 12861 11242 14673 11252
rect 2481 10954 2681 10964
rect 2481 10898 2491 10954
rect 2547 10898 2615 10954
rect 2671 10898 2681 10954
rect 2481 10830 2681 10898
rect 2481 10774 2491 10830
rect 2547 10774 2615 10830
rect 2671 10774 2681 10830
rect 2481 10706 2681 10774
rect 2481 10650 2491 10706
rect 2547 10650 2615 10706
rect 2671 10650 2681 10706
rect 2481 10582 2681 10650
rect 2481 10526 2491 10582
rect 2547 10526 2615 10582
rect 2671 10526 2681 10582
rect 2481 10458 2681 10526
rect 2481 10402 2491 10458
rect 2547 10402 2615 10458
rect 2671 10402 2681 10458
rect 2481 10334 2681 10402
rect 2481 10278 2491 10334
rect 2547 10278 2615 10334
rect 2671 10278 2681 10334
rect 2481 10210 2681 10278
rect 2481 10154 2491 10210
rect 2547 10154 2615 10210
rect 2671 10154 2681 10210
rect 2481 10086 2681 10154
rect 2481 10030 2491 10086
rect 2547 10030 2615 10086
rect 2671 10030 2681 10086
rect 2481 9962 2681 10030
rect 2481 9906 2491 9962
rect 2547 9906 2615 9962
rect 2671 9906 2681 9962
rect 2481 9838 2681 9906
rect 2481 9782 2491 9838
rect 2547 9782 2615 9838
rect 2671 9782 2681 9838
rect 2481 9714 2681 9782
rect 2481 9658 2491 9714
rect 2547 9658 2615 9714
rect 2671 9658 2681 9714
rect 2481 9590 2681 9658
rect 2481 9534 2491 9590
rect 2547 9534 2615 9590
rect 2671 9534 2681 9590
rect 2481 9466 2681 9534
rect 2481 9410 2491 9466
rect 2547 9410 2615 9466
rect 2671 9410 2681 9466
rect 2481 9342 2681 9410
rect 2481 9286 2491 9342
rect 2547 9286 2615 9342
rect 2671 9286 2681 9342
rect 2481 9218 2681 9286
rect 2481 9162 2491 9218
rect 2547 9162 2615 9218
rect 2671 9162 2681 9218
rect 2481 9094 2681 9162
rect 2481 9038 2491 9094
rect 2547 9038 2615 9094
rect 2671 9038 2681 9094
rect 2481 8970 2681 9038
rect 2481 8914 2491 8970
rect 2547 8914 2615 8970
rect 2671 8914 2681 8970
rect 2481 8846 2681 8914
rect 2481 8790 2491 8846
rect 2547 8790 2615 8846
rect 2671 8790 2681 8846
rect 2481 8722 2681 8790
rect 2481 8666 2491 8722
rect 2547 8666 2615 8722
rect 2671 8666 2681 8722
rect 2481 8598 2681 8666
rect 2481 8542 2491 8598
rect 2547 8542 2615 8598
rect 2671 8542 2681 8598
rect 2481 8474 2681 8542
rect 2481 8418 2491 8474
rect 2547 8418 2615 8474
rect 2671 8418 2681 8474
rect 2481 8350 2681 8418
rect 2481 8294 2491 8350
rect 2547 8294 2615 8350
rect 2671 8294 2681 8350
rect 2481 8226 2681 8294
rect 2481 8170 2491 8226
rect 2547 8170 2615 8226
rect 2671 8170 2681 8226
rect 2481 8102 2681 8170
rect 2481 8046 2491 8102
rect 2547 8046 2615 8102
rect 2671 8046 2681 8102
rect 2481 8036 2681 8046
rect 4851 10954 5051 10964
rect 4851 10898 4861 10954
rect 4917 10898 4985 10954
rect 5041 10898 5051 10954
rect 4851 10830 5051 10898
rect 4851 10774 4861 10830
rect 4917 10774 4985 10830
rect 5041 10774 5051 10830
rect 4851 10706 5051 10774
rect 4851 10650 4861 10706
rect 4917 10650 4985 10706
rect 5041 10650 5051 10706
rect 4851 10582 5051 10650
rect 4851 10526 4861 10582
rect 4917 10526 4985 10582
rect 5041 10526 5051 10582
rect 4851 10458 5051 10526
rect 4851 10402 4861 10458
rect 4917 10402 4985 10458
rect 5041 10402 5051 10458
rect 4851 10334 5051 10402
rect 4851 10278 4861 10334
rect 4917 10278 4985 10334
rect 5041 10278 5051 10334
rect 4851 10210 5051 10278
rect 4851 10154 4861 10210
rect 4917 10154 4985 10210
rect 5041 10154 5051 10210
rect 4851 10086 5051 10154
rect 4851 10030 4861 10086
rect 4917 10030 4985 10086
rect 5041 10030 5051 10086
rect 4851 9962 5051 10030
rect 4851 9906 4861 9962
rect 4917 9906 4985 9962
rect 5041 9906 5051 9962
rect 4851 9838 5051 9906
rect 4851 9782 4861 9838
rect 4917 9782 4985 9838
rect 5041 9782 5051 9838
rect 4851 9714 5051 9782
rect 4851 9658 4861 9714
rect 4917 9658 4985 9714
rect 5041 9658 5051 9714
rect 4851 9590 5051 9658
rect 4851 9534 4861 9590
rect 4917 9534 4985 9590
rect 5041 9534 5051 9590
rect 4851 9466 5051 9534
rect 4851 9410 4861 9466
rect 4917 9410 4985 9466
rect 5041 9410 5051 9466
rect 4851 9342 5051 9410
rect 4851 9286 4861 9342
rect 4917 9286 4985 9342
rect 5041 9286 5051 9342
rect 4851 9218 5051 9286
rect 4851 9162 4861 9218
rect 4917 9162 4985 9218
rect 5041 9162 5051 9218
rect 4851 9094 5051 9162
rect 4851 9038 4861 9094
rect 4917 9038 4985 9094
rect 5041 9038 5051 9094
rect 4851 8970 5051 9038
rect 4851 8914 4861 8970
rect 4917 8914 4985 8970
rect 5041 8914 5051 8970
rect 4851 8846 5051 8914
rect 4851 8790 4861 8846
rect 4917 8790 4985 8846
rect 5041 8790 5051 8846
rect 4851 8722 5051 8790
rect 4851 8666 4861 8722
rect 4917 8666 4985 8722
rect 5041 8666 5051 8722
rect 4851 8598 5051 8666
rect 4851 8542 4861 8598
rect 4917 8542 4985 8598
rect 5041 8542 5051 8598
rect 4851 8474 5051 8542
rect 4851 8418 4861 8474
rect 4917 8418 4985 8474
rect 5041 8418 5051 8474
rect 4851 8350 5051 8418
rect 4851 8294 4861 8350
rect 4917 8294 4985 8350
rect 5041 8294 5051 8350
rect 4851 8226 5051 8294
rect 4851 8170 4861 8226
rect 4917 8170 4985 8226
rect 5041 8170 5051 8226
rect 4851 8102 5051 8170
rect 4851 8046 4861 8102
rect 4917 8046 4985 8102
rect 5041 8046 5051 8102
rect 4851 8036 5051 8046
rect 7265 10954 7713 10964
rect 7265 10898 7275 10954
rect 7331 10898 7399 10954
rect 7455 10898 7523 10954
rect 7579 10898 7647 10954
rect 7703 10898 7713 10954
rect 7265 10830 7713 10898
rect 7265 10774 7275 10830
rect 7331 10774 7399 10830
rect 7455 10774 7523 10830
rect 7579 10774 7647 10830
rect 7703 10774 7713 10830
rect 7265 10706 7713 10774
rect 7265 10650 7275 10706
rect 7331 10650 7399 10706
rect 7455 10650 7523 10706
rect 7579 10650 7647 10706
rect 7703 10650 7713 10706
rect 7265 10582 7713 10650
rect 7265 10526 7275 10582
rect 7331 10526 7399 10582
rect 7455 10526 7523 10582
rect 7579 10526 7647 10582
rect 7703 10526 7713 10582
rect 7265 10458 7713 10526
rect 7265 10402 7275 10458
rect 7331 10402 7399 10458
rect 7455 10402 7523 10458
rect 7579 10402 7647 10458
rect 7703 10402 7713 10458
rect 7265 10334 7713 10402
rect 7265 10278 7275 10334
rect 7331 10278 7399 10334
rect 7455 10278 7523 10334
rect 7579 10278 7647 10334
rect 7703 10278 7713 10334
rect 7265 10210 7713 10278
rect 7265 10154 7275 10210
rect 7331 10154 7399 10210
rect 7455 10154 7523 10210
rect 7579 10154 7647 10210
rect 7703 10154 7713 10210
rect 7265 10086 7713 10154
rect 7265 10030 7275 10086
rect 7331 10030 7399 10086
rect 7455 10030 7523 10086
rect 7579 10030 7647 10086
rect 7703 10030 7713 10086
rect 7265 9962 7713 10030
rect 7265 9906 7275 9962
rect 7331 9906 7399 9962
rect 7455 9906 7523 9962
rect 7579 9906 7647 9962
rect 7703 9906 7713 9962
rect 7265 9838 7713 9906
rect 7265 9782 7275 9838
rect 7331 9782 7399 9838
rect 7455 9782 7523 9838
rect 7579 9782 7647 9838
rect 7703 9782 7713 9838
rect 7265 9714 7713 9782
rect 7265 9658 7275 9714
rect 7331 9658 7399 9714
rect 7455 9658 7523 9714
rect 7579 9658 7647 9714
rect 7703 9658 7713 9714
rect 7265 9590 7713 9658
rect 7265 9534 7275 9590
rect 7331 9534 7399 9590
rect 7455 9534 7523 9590
rect 7579 9534 7647 9590
rect 7703 9534 7713 9590
rect 7265 9466 7713 9534
rect 7265 9410 7275 9466
rect 7331 9410 7399 9466
rect 7455 9410 7523 9466
rect 7579 9410 7647 9466
rect 7703 9410 7713 9466
rect 7265 9342 7713 9410
rect 7265 9286 7275 9342
rect 7331 9286 7399 9342
rect 7455 9286 7523 9342
rect 7579 9286 7647 9342
rect 7703 9286 7713 9342
rect 7265 9218 7713 9286
rect 7265 9162 7275 9218
rect 7331 9162 7399 9218
rect 7455 9162 7523 9218
rect 7579 9162 7647 9218
rect 7703 9162 7713 9218
rect 7265 9094 7713 9162
rect 7265 9038 7275 9094
rect 7331 9038 7399 9094
rect 7455 9038 7523 9094
rect 7579 9038 7647 9094
rect 7703 9038 7713 9094
rect 7265 8970 7713 9038
rect 7265 8914 7275 8970
rect 7331 8914 7399 8970
rect 7455 8914 7523 8970
rect 7579 8914 7647 8970
rect 7703 8914 7713 8970
rect 7265 8846 7713 8914
rect 7265 8790 7275 8846
rect 7331 8790 7399 8846
rect 7455 8790 7523 8846
rect 7579 8790 7647 8846
rect 7703 8790 7713 8846
rect 7265 8722 7713 8790
rect 7265 8666 7275 8722
rect 7331 8666 7399 8722
rect 7455 8666 7523 8722
rect 7579 8666 7647 8722
rect 7703 8666 7713 8722
rect 7265 8598 7713 8666
rect 7265 8542 7275 8598
rect 7331 8542 7399 8598
rect 7455 8542 7523 8598
rect 7579 8542 7647 8598
rect 7703 8542 7713 8598
rect 7265 8474 7713 8542
rect 7265 8418 7275 8474
rect 7331 8418 7399 8474
rect 7455 8418 7523 8474
rect 7579 8418 7647 8474
rect 7703 8418 7713 8474
rect 7265 8350 7713 8418
rect 7265 8294 7275 8350
rect 7331 8294 7399 8350
rect 7455 8294 7523 8350
rect 7579 8294 7647 8350
rect 7703 8294 7713 8350
rect 7265 8226 7713 8294
rect 7265 8170 7275 8226
rect 7331 8170 7399 8226
rect 7455 8170 7523 8226
rect 7579 8170 7647 8226
rect 7703 8170 7713 8226
rect 7265 8102 7713 8170
rect 7265 8046 7275 8102
rect 7331 8046 7399 8102
rect 7455 8046 7523 8102
rect 7579 8046 7647 8102
rect 7703 8046 7713 8102
rect 7265 8036 7713 8046
rect 9927 10954 10127 10964
rect 9927 10898 9937 10954
rect 9993 10898 10061 10954
rect 10117 10898 10127 10954
rect 9927 10830 10127 10898
rect 9927 10774 9937 10830
rect 9993 10774 10061 10830
rect 10117 10774 10127 10830
rect 9927 10706 10127 10774
rect 9927 10650 9937 10706
rect 9993 10650 10061 10706
rect 10117 10650 10127 10706
rect 9927 10582 10127 10650
rect 9927 10526 9937 10582
rect 9993 10526 10061 10582
rect 10117 10526 10127 10582
rect 9927 10458 10127 10526
rect 9927 10402 9937 10458
rect 9993 10402 10061 10458
rect 10117 10402 10127 10458
rect 9927 10334 10127 10402
rect 9927 10278 9937 10334
rect 9993 10278 10061 10334
rect 10117 10278 10127 10334
rect 9927 10210 10127 10278
rect 9927 10154 9937 10210
rect 9993 10154 10061 10210
rect 10117 10154 10127 10210
rect 9927 10086 10127 10154
rect 9927 10030 9937 10086
rect 9993 10030 10061 10086
rect 10117 10030 10127 10086
rect 9927 9962 10127 10030
rect 9927 9906 9937 9962
rect 9993 9906 10061 9962
rect 10117 9906 10127 9962
rect 9927 9838 10127 9906
rect 9927 9782 9937 9838
rect 9993 9782 10061 9838
rect 10117 9782 10127 9838
rect 9927 9714 10127 9782
rect 9927 9658 9937 9714
rect 9993 9658 10061 9714
rect 10117 9658 10127 9714
rect 9927 9590 10127 9658
rect 9927 9534 9937 9590
rect 9993 9534 10061 9590
rect 10117 9534 10127 9590
rect 9927 9466 10127 9534
rect 9927 9410 9937 9466
rect 9993 9410 10061 9466
rect 10117 9410 10127 9466
rect 9927 9342 10127 9410
rect 9927 9286 9937 9342
rect 9993 9286 10061 9342
rect 10117 9286 10127 9342
rect 9927 9218 10127 9286
rect 9927 9162 9937 9218
rect 9993 9162 10061 9218
rect 10117 9162 10127 9218
rect 9927 9094 10127 9162
rect 9927 9038 9937 9094
rect 9993 9038 10061 9094
rect 10117 9038 10127 9094
rect 9927 8970 10127 9038
rect 9927 8914 9937 8970
rect 9993 8914 10061 8970
rect 10117 8914 10127 8970
rect 9927 8846 10127 8914
rect 9927 8790 9937 8846
rect 9993 8790 10061 8846
rect 10117 8790 10127 8846
rect 9927 8722 10127 8790
rect 9927 8666 9937 8722
rect 9993 8666 10061 8722
rect 10117 8666 10127 8722
rect 9927 8598 10127 8666
rect 9927 8542 9937 8598
rect 9993 8542 10061 8598
rect 10117 8542 10127 8598
rect 9927 8474 10127 8542
rect 9927 8418 9937 8474
rect 9993 8418 10061 8474
rect 10117 8418 10127 8474
rect 9927 8350 10127 8418
rect 9927 8294 9937 8350
rect 9993 8294 10061 8350
rect 10117 8294 10127 8350
rect 9927 8226 10127 8294
rect 9927 8170 9937 8226
rect 9993 8170 10061 8226
rect 10117 8170 10127 8226
rect 9927 8102 10127 8170
rect 9927 8046 9937 8102
rect 9993 8046 10061 8102
rect 10117 8046 10127 8102
rect 9927 8036 10127 8046
rect 12297 10954 12497 10964
rect 12297 10898 12307 10954
rect 12363 10898 12431 10954
rect 12487 10898 12497 10954
rect 12297 10830 12497 10898
rect 12297 10774 12307 10830
rect 12363 10774 12431 10830
rect 12487 10774 12497 10830
rect 12297 10706 12497 10774
rect 12297 10650 12307 10706
rect 12363 10650 12431 10706
rect 12487 10650 12497 10706
rect 12297 10582 12497 10650
rect 12297 10526 12307 10582
rect 12363 10526 12431 10582
rect 12487 10526 12497 10582
rect 12297 10458 12497 10526
rect 12297 10402 12307 10458
rect 12363 10402 12431 10458
rect 12487 10402 12497 10458
rect 12297 10334 12497 10402
rect 12297 10278 12307 10334
rect 12363 10278 12431 10334
rect 12487 10278 12497 10334
rect 12297 10210 12497 10278
rect 12297 10154 12307 10210
rect 12363 10154 12431 10210
rect 12487 10154 12497 10210
rect 12297 10086 12497 10154
rect 12297 10030 12307 10086
rect 12363 10030 12431 10086
rect 12487 10030 12497 10086
rect 12297 9962 12497 10030
rect 12297 9906 12307 9962
rect 12363 9906 12431 9962
rect 12487 9906 12497 9962
rect 12297 9838 12497 9906
rect 12297 9782 12307 9838
rect 12363 9782 12431 9838
rect 12487 9782 12497 9838
rect 12297 9714 12497 9782
rect 12297 9658 12307 9714
rect 12363 9658 12431 9714
rect 12487 9658 12497 9714
rect 12297 9590 12497 9658
rect 12297 9534 12307 9590
rect 12363 9534 12431 9590
rect 12487 9534 12497 9590
rect 12297 9466 12497 9534
rect 12297 9410 12307 9466
rect 12363 9410 12431 9466
rect 12487 9410 12497 9466
rect 12297 9342 12497 9410
rect 12297 9286 12307 9342
rect 12363 9286 12431 9342
rect 12487 9286 12497 9342
rect 12297 9218 12497 9286
rect 12297 9162 12307 9218
rect 12363 9162 12431 9218
rect 12487 9162 12497 9218
rect 12297 9094 12497 9162
rect 12297 9038 12307 9094
rect 12363 9038 12431 9094
rect 12487 9038 12497 9094
rect 12297 8970 12497 9038
rect 12297 8914 12307 8970
rect 12363 8914 12431 8970
rect 12487 8914 12497 8970
rect 12297 8846 12497 8914
rect 12297 8790 12307 8846
rect 12363 8790 12431 8846
rect 12487 8790 12497 8846
rect 12297 8722 12497 8790
rect 12297 8666 12307 8722
rect 12363 8666 12431 8722
rect 12487 8666 12497 8722
rect 12297 8598 12497 8666
rect 12297 8542 12307 8598
rect 12363 8542 12431 8598
rect 12487 8542 12497 8598
rect 12297 8474 12497 8542
rect 12297 8418 12307 8474
rect 12363 8418 12431 8474
rect 12487 8418 12497 8474
rect 12297 8350 12497 8418
rect 12297 8294 12307 8350
rect 12363 8294 12431 8350
rect 12487 8294 12497 8350
rect 12297 8226 12497 8294
rect 12297 8170 12307 8226
rect 12363 8170 12431 8226
rect 12487 8170 12497 8226
rect 12297 8102 12497 8170
rect 12297 8046 12307 8102
rect 12363 8046 12431 8102
rect 12487 8046 12497 8102
rect 12297 8036 12497 8046
rect 2481 7754 2681 7764
rect 2481 7698 2491 7754
rect 2547 7698 2615 7754
rect 2671 7698 2681 7754
rect 2481 7630 2681 7698
rect 2481 7574 2491 7630
rect 2547 7574 2615 7630
rect 2671 7574 2681 7630
rect 2481 7506 2681 7574
rect 2481 7450 2491 7506
rect 2547 7450 2615 7506
rect 2671 7450 2681 7506
rect 2481 7382 2681 7450
rect 2481 7326 2491 7382
rect 2547 7326 2615 7382
rect 2671 7326 2681 7382
rect 2481 7258 2681 7326
rect 2481 7202 2491 7258
rect 2547 7202 2615 7258
rect 2671 7202 2681 7258
rect 2481 7134 2681 7202
rect 2481 7078 2491 7134
rect 2547 7078 2615 7134
rect 2671 7078 2681 7134
rect 2481 7010 2681 7078
rect 2481 6954 2491 7010
rect 2547 6954 2615 7010
rect 2671 6954 2681 7010
rect 2481 6886 2681 6954
rect 2481 6830 2491 6886
rect 2547 6830 2615 6886
rect 2671 6830 2681 6886
rect 2481 6762 2681 6830
rect 2481 6706 2491 6762
rect 2547 6706 2615 6762
rect 2671 6706 2681 6762
rect 2481 6638 2681 6706
rect 2481 6582 2491 6638
rect 2547 6582 2615 6638
rect 2671 6582 2681 6638
rect 2481 6514 2681 6582
rect 2481 6458 2491 6514
rect 2547 6458 2615 6514
rect 2671 6458 2681 6514
rect 2481 6390 2681 6458
rect 2481 6334 2491 6390
rect 2547 6334 2615 6390
rect 2671 6334 2681 6390
rect 2481 6266 2681 6334
rect 2481 6210 2491 6266
rect 2547 6210 2615 6266
rect 2671 6210 2681 6266
rect 2481 6142 2681 6210
rect 2481 6086 2491 6142
rect 2547 6086 2615 6142
rect 2671 6086 2681 6142
rect 2481 6018 2681 6086
rect 2481 5962 2491 6018
rect 2547 5962 2615 6018
rect 2671 5962 2681 6018
rect 2481 5894 2681 5962
rect 2481 5838 2491 5894
rect 2547 5838 2615 5894
rect 2671 5838 2681 5894
rect 2481 5770 2681 5838
rect 2481 5714 2491 5770
rect 2547 5714 2615 5770
rect 2671 5714 2681 5770
rect 2481 5646 2681 5714
rect 2481 5590 2491 5646
rect 2547 5590 2615 5646
rect 2671 5590 2681 5646
rect 2481 5522 2681 5590
rect 2481 5466 2491 5522
rect 2547 5466 2615 5522
rect 2671 5466 2681 5522
rect 2481 5398 2681 5466
rect 2481 5342 2491 5398
rect 2547 5342 2615 5398
rect 2671 5342 2681 5398
rect 2481 5274 2681 5342
rect 2481 5218 2491 5274
rect 2547 5218 2615 5274
rect 2671 5218 2681 5274
rect 2481 5150 2681 5218
rect 2481 5094 2491 5150
rect 2547 5094 2615 5150
rect 2671 5094 2681 5150
rect 2481 5026 2681 5094
rect 2481 4970 2491 5026
rect 2547 4970 2615 5026
rect 2671 4970 2681 5026
rect 2481 4902 2681 4970
rect 2481 4846 2491 4902
rect 2547 4846 2615 4902
rect 2671 4846 2681 4902
rect 2481 4836 2681 4846
rect 4851 7754 5051 7764
rect 4851 7698 4861 7754
rect 4917 7698 4985 7754
rect 5041 7698 5051 7754
rect 4851 7630 5051 7698
rect 4851 7574 4861 7630
rect 4917 7574 4985 7630
rect 5041 7574 5051 7630
rect 4851 7506 5051 7574
rect 4851 7450 4861 7506
rect 4917 7450 4985 7506
rect 5041 7450 5051 7506
rect 4851 7382 5051 7450
rect 4851 7326 4861 7382
rect 4917 7326 4985 7382
rect 5041 7326 5051 7382
rect 4851 7258 5051 7326
rect 4851 7202 4861 7258
rect 4917 7202 4985 7258
rect 5041 7202 5051 7258
rect 4851 7134 5051 7202
rect 4851 7078 4861 7134
rect 4917 7078 4985 7134
rect 5041 7078 5051 7134
rect 4851 7010 5051 7078
rect 4851 6954 4861 7010
rect 4917 6954 4985 7010
rect 5041 6954 5051 7010
rect 4851 6886 5051 6954
rect 4851 6830 4861 6886
rect 4917 6830 4985 6886
rect 5041 6830 5051 6886
rect 4851 6762 5051 6830
rect 4851 6706 4861 6762
rect 4917 6706 4985 6762
rect 5041 6706 5051 6762
rect 4851 6638 5051 6706
rect 4851 6582 4861 6638
rect 4917 6582 4985 6638
rect 5041 6582 5051 6638
rect 4851 6514 5051 6582
rect 4851 6458 4861 6514
rect 4917 6458 4985 6514
rect 5041 6458 5051 6514
rect 4851 6390 5051 6458
rect 4851 6334 4861 6390
rect 4917 6334 4985 6390
rect 5041 6334 5051 6390
rect 4851 6266 5051 6334
rect 4851 6210 4861 6266
rect 4917 6210 4985 6266
rect 5041 6210 5051 6266
rect 4851 6142 5051 6210
rect 4851 6086 4861 6142
rect 4917 6086 4985 6142
rect 5041 6086 5051 6142
rect 4851 6018 5051 6086
rect 4851 5962 4861 6018
rect 4917 5962 4985 6018
rect 5041 5962 5051 6018
rect 4851 5894 5051 5962
rect 4851 5838 4861 5894
rect 4917 5838 4985 5894
rect 5041 5838 5051 5894
rect 4851 5770 5051 5838
rect 4851 5714 4861 5770
rect 4917 5714 4985 5770
rect 5041 5714 5051 5770
rect 4851 5646 5051 5714
rect 4851 5590 4861 5646
rect 4917 5590 4985 5646
rect 5041 5590 5051 5646
rect 4851 5522 5051 5590
rect 4851 5466 4861 5522
rect 4917 5466 4985 5522
rect 5041 5466 5051 5522
rect 4851 5398 5051 5466
rect 4851 5342 4861 5398
rect 4917 5342 4985 5398
rect 5041 5342 5051 5398
rect 4851 5274 5051 5342
rect 4851 5218 4861 5274
rect 4917 5218 4985 5274
rect 5041 5218 5051 5274
rect 4851 5150 5051 5218
rect 4851 5094 4861 5150
rect 4917 5094 4985 5150
rect 5041 5094 5051 5150
rect 4851 5026 5051 5094
rect 4851 4970 4861 5026
rect 4917 4970 4985 5026
rect 5041 4970 5051 5026
rect 4851 4902 5051 4970
rect 4851 4846 4861 4902
rect 4917 4846 4985 4902
rect 5041 4846 5051 4902
rect 4851 4836 5051 4846
rect 7265 7754 7713 7764
rect 7265 7698 7275 7754
rect 7331 7698 7399 7754
rect 7455 7698 7523 7754
rect 7579 7698 7647 7754
rect 7703 7698 7713 7754
rect 7265 7630 7713 7698
rect 7265 7574 7275 7630
rect 7331 7574 7399 7630
rect 7455 7574 7523 7630
rect 7579 7574 7647 7630
rect 7703 7574 7713 7630
rect 7265 7506 7713 7574
rect 7265 7450 7275 7506
rect 7331 7450 7399 7506
rect 7455 7450 7523 7506
rect 7579 7450 7647 7506
rect 7703 7450 7713 7506
rect 7265 7382 7713 7450
rect 7265 7326 7275 7382
rect 7331 7326 7399 7382
rect 7455 7326 7523 7382
rect 7579 7326 7647 7382
rect 7703 7326 7713 7382
rect 7265 7258 7713 7326
rect 7265 7202 7275 7258
rect 7331 7202 7399 7258
rect 7455 7202 7523 7258
rect 7579 7202 7647 7258
rect 7703 7202 7713 7258
rect 7265 7134 7713 7202
rect 7265 7078 7275 7134
rect 7331 7078 7399 7134
rect 7455 7078 7523 7134
rect 7579 7078 7647 7134
rect 7703 7078 7713 7134
rect 7265 7010 7713 7078
rect 7265 6954 7275 7010
rect 7331 6954 7399 7010
rect 7455 6954 7523 7010
rect 7579 6954 7647 7010
rect 7703 6954 7713 7010
rect 7265 6886 7713 6954
rect 7265 6830 7275 6886
rect 7331 6830 7399 6886
rect 7455 6830 7523 6886
rect 7579 6830 7647 6886
rect 7703 6830 7713 6886
rect 7265 6762 7713 6830
rect 7265 6706 7275 6762
rect 7331 6706 7399 6762
rect 7455 6706 7523 6762
rect 7579 6706 7647 6762
rect 7703 6706 7713 6762
rect 7265 6638 7713 6706
rect 7265 6582 7275 6638
rect 7331 6582 7399 6638
rect 7455 6582 7523 6638
rect 7579 6582 7647 6638
rect 7703 6582 7713 6638
rect 7265 6514 7713 6582
rect 7265 6458 7275 6514
rect 7331 6458 7399 6514
rect 7455 6458 7523 6514
rect 7579 6458 7647 6514
rect 7703 6458 7713 6514
rect 7265 6390 7713 6458
rect 7265 6334 7275 6390
rect 7331 6334 7399 6390
rect 7455 6334 7523 6390
rect 7579 6334 7647 6390
rect 7703 6334 7713 6390
rect 7265 6266 7713 6334
rect 7265 6210 7275 6266
rect 7331 6210 7399 6266
rect 7455 6210 7523 6266
rect 7579 6210 7647 6266
rect 7703 6210 7713 6266
rect 7265 6142 7713 6210
rect 7265 6086 7275 6142
rect 7331 6086 7399 6142
rect 7455 6086 7523 6142
rect 7579 6086 7647 6142
rect 7703 6086 7713 6142
rect 7265 6018 7713 6086
rect 7265 5962 7275 6018
rect 7331 5962 7399 6018
rect 7455 5962 7523 6018
rect 7579 5962 7647 6018
rect 7703 5962 7713 6018
rect 7265 5894 7713 5962
rect 7265 5838 7275 5894
rect 7331 5838 7399 5894
rect 7455 5838 7523 5894
rect 7579 5838 7647 5894
rect 7703 5838 7713 5894
rect 7265 5770 7713 5838
rect 7265 5714 7275 5770
rect 7331 5714 7399 5770
rect 7455 5714 7523 5770
rect 7579 5714 7647 5770
rect 7703 5714 7713 5770
rect 7265 5646 7713 5714
rect 7265 5590 7275 5646
rect 7331 5590 7399 5646
rect 7455 5590 7523 5646
rect 7579 5590 7647 5646
rect 7703 5590 7713 5646
rect 7265 5522 7713 5590
rect 7265 5466 7275 5522
rect 7331 5466 7399 5522
rect 7455 5466 7523 5522
rect 7579 5466 7647 5522
rect 7703 5466 7713 5522
rect 7265 5398 7713 5466
rect 7265 5342 7275 5398
rect 7331 5342 7399 5398
rect 7455 5342 7523 5398
rect 7579 5342 7647 5398
rect 7703 5342 7713 5398
rect 7265 5274 7713 5342
rect 7265 5218 7275 5274
rect 7331 5218 7399 5274
rect 7455 5218 7523 5274
rect 7579 5218 7647 5274
rect 7703 5218 7713 5274
rect 7265 5150 7713 5218
rect 7265 5094 7275 5150
rect 7331 5094 7399 5150
rect 7455 5094 7523 5150
rect 7579 5094 7647 5150
rect 7703 5094 7713 5150
rect 7265 5026 7713 5094
rect 7265 4970 7275 5026
rect 7331 4970 7399 5026
rect 7455 4970 7523 5026
rect 7579 4970 7647 5026
rect 7703 4970 7713 5026
rect 7265 4902 7713 4970
rect 7265 4846 7275 4902
rect 7331 4846 7399 4902
rect 7455 4846 7523 4902
rect 7579 4846 7647 4902
rect 7703 4846 7713 4902
rect 7265 4836 7713 4846
rect 9927 7754 10127 7764
rect 9927 7698 9937 7754
rect 9993 7698 10061 7754
rect 10117 7698 10127 7754
rect 9927 7630 10127 7698
rect 9927 7574 9937 7630
rect 9993 7574 10061 7630
rect 10117 7574 10127 7630
rect 9927 7506 10127 7574
rect 9927 7450 9937 7506
rect 9993 7450 10061 7506
rect 10117 7450 10127 7506
rect 9927 7382 10127 7450
rect 9927 7326 9937 7382
rect 9993 7326 10061 7382
rect 10117 7326 10127 7382
rect 9927 7258 10127 7326
rect 9927 7202 9937 7258
rect 9993 7202 10061 7258
rect 10117 7202 10127 7258
rect 9927 7134 10127 7202
rect 9927 7078 9937 7134
rect 9993 7078 10061 7134
rect 10117 7078 10127 7134
rect 9927 7010 10127 7078
rect 9927 6954 9937 7010
rect 9993 6954 10061 7010
rect 10117 6954 10127 7010
rect 9927 6886 10127 6954
rect 9927 6830 9937 6886
rect 9993 6830 10061 6886
rect 10117 6830 10127 6886
rect 9927 6762 10127 6830
rect 9927 6706 9937 6762
rect 9993 6706 10061 6762
rect 10117 6706 10127 6762
rect 9927 6638 10127 6706
rect 9927 6582 9937 6638
rect 9993 6582 10061 6638
rect 10117 6582 10127 6638
rect 9927 6514 10127 6582
rect 9927 6458 9937 6514
rect 9993 6458 10061 6514
rect 10117 6458 10127 6514
rect 9927 6390 10127 6458
rect 9927 6334 9937 6390
rect 9993 6334 10061 6390
rect 10117 6334 10127 6390
rect 9927 6266 10127 6334
rect 9927 6210 9937 6266
rect 9993 6210 10061 6266
rect 10117 6210 10127 6266
rect 9927 6142 10127 6210
rect 9927 6086 9937 6142
rect 9993 6086 10061 6142
rect 10117 6086 10127 6142
rect 9927 6018 10127 6086
rect 9927 5962 9937 6018
rect 9993 5962 10061 6018
rect 10117 5962 10127 6018
rect 9927 5894 10127 5962
rect 9927 5838 9937 5894
rect 9993 5838 10061 5894
rect 10117 5838 10127 5894
rect 9927 5770 10127 5838
rect 9927 5714 9937 5770
rect 9993 5714 10061 5770
rect 10117 5714 10127 5770
rect 9927 5646 10127 5714
rect 9927 5590 9937 5646
rect 9993 5590 10061 5646
rect 10117 5590 10127 5646
rect 9927 5522 10127 5590
rect 9927 5466 9937 5522
rect 9993 5466 10061 5522
rect 10117 5466 10127 5522
rect 9927 5398 10127 5466
rect 9927 5342 9937 5398
rect 9993 5342 10061 5398
rect 10117 5342 10127 5398
rect 9927 5274 10127 5342
rect 9927 5218 9937 5274
rect 9993 5218 10061 5274
rect 10117 5218 10127 5274
rect 9927 5150 10127 5218
rect 9927 5094 9937 5150
rect 9993 5094 10061 5150
rect 10117 5094 10127 5150
rect 9927 5026 10127 5094
rect 9927 4970 9937 5026
rect 9993 4970 10061 5026
rect 10117 4970 10127 5026
rect 9927 4902 10127 4970
rect 9927 4846 9937 4902
rect 9993 4846 10061 4902
rect 10117 4846 10127 4902
rect 9927 4836 10127 4846
rect 12297 7754 12497 7764
rect 12297 7698 12307 7754
rect 12363 7698 12431 7754
rect 12487 7698 12497 7754
rect 12297 7630 12497 7698
rect 12297 7574 12307 7630
rect 12363 7574 12431 7630
rect 12487 7574 12497 7630
rect 12297 7506 12497 7574
rect 12297 7450 12307 7506
rect 12363 7450 12431 7506
rect 12487 7450 12497 7506
rect 12297 7382 12497 7450
rect 12297 7326 12307 7382
rect 12363 7326 12431 7382
rect 12487 7326 12497 7382
rect 12297 7258 12497 7326
rect 12297 7202 12307 7258
rect 12363 7202 12431 7258
rect 12487 7202 12497 7258
rect 12297 7134 12497 7202
rect 12297 7078 12307 7134
rect 12363 7078 12431 7134
rect 12487 7078 12497 7134
rect 12297 7010 12497 7078
rect 12297 6954 12307 7010
rect 12363 6954 12431 7010
rect 12487 6954 12497 7010
rect 12297 6886 12497 6954
rect 12297 6830 12307 6886
rect 12363 6830 12431 6886
rect 12487 6830 12497 6886
rect 12297 6762 12497 6830
rect 12297 6706 12307 6762
rect 12363 6706 12431 6762
rect 12487 6706 12497 6762
rect 12297 6638 12497 6706
rect 12297 6582 12307 6638
rect 12363 6582 12431 6638
rect 12487 6582 12497 6638
rect 12297 6514 12497 6582
rect 12297 6458 12307 6514
rect 12363 6458 12431 6514
rect 12487 6458 12497 6514
rect 12297 6390 12497 6458
rect 12297 6334 12307 6390
rect 12363 6334 12431 6390
rect 12487 6334 12497 6390
rect 12297 6266 12497 6334
rect 12297 6210 12307 6266
rect 12363 6210 12431 6266
rect 12487 6210 12497 6266
rect 12297 6142 12497 6210
rect 12297 6086 12307 6142
rect 12363 6086 12431 6142
rect 12487 6086 12497 6142
rect 12297 6018 12497 6086
rect 12297 5962 12307 6018
rect 12363 5962 12431 6018
rect 12487 5962 12497 6018
rect 12297 5894 12497 5962
rect 12297 5838 12307 5894
rect 12363 5838 12431 5894
rect 12487 5838 12497 5894
rect 12297 5770 12497 5838
rect 12297 5714 12307 5770
rect 12363 5714 12431 5770
rect 12487 5714 12497 5770
rect 12297 5646 12497 5714
rect 12297 5590 12307 5646
rect 12363 5590 12431 5646
rect 12487 5590 12497 5646
rect 12297 5522 12497 5590
rect 12297 5466 12307 5522
rect 12363 5466 12431 5522
rect 12487 5466 12497 5522
rect 12297 5398 12497 5466
rect 12297 5342 12307 5398
rect 12363 5342 12431 5398
rect 12487 5342 12497 5398
rect 12297 5274 12497 5342
rect 12297 5218 12307 5274
rect 12363 5218 12431 5274
rect 12487 5218 12497 5274
rect 12297 5150 12497 5218
rect 12297 5094 12307 5150
rect 12363 5094 12431 5150
rect 12487 5094 12497 5150
rect 12297 5026 12497 5094
rect 12297 4970 12307 5026
rect 12363 4970 12431 5026
rect 12487 4970 12497 5026
rect 12297 4902 12497 4970
rect 12297 4846 12307 4902
rect 12363 4846 12431 4902
rect 12487 4846 12497 4902
rect 12297 4836 12497 4846
rect 2481 4554 2681 4564
rect 2481 4498 2491 4554
rect 2547 4498 2615 4554
rect 2671 4498 2681 4554
rect 2481 4430 2681 4498
rect 2481 4374 2491 4430
rect 2547 4374 2615 4430
rect 2671 4374 2681 4430
rect 2481 4306 2681 4374
rect 2481 4250 2491 4306
rect 2547 4250 2615 4306
rect 2671 4250 2681 4306
rect 2481 4182 2681 4250
rect 2481 4126 2491 4182
rect 2547 4126 2615 4182
rect 2671 4126 2681 4182
rect 2481 4058 2681 4126
rect 2481 4002 2491 4058
rect 2547 4002 2615 4058
rect 2671 4002 2681 4058
rect 2481 3934 2681 4002
rect 2481 3878 2491 3934
rect 2547 3878 2615 3934
rect 2671 3878 2681 3934
rect 2481 3810 2681 3878
rect 2481 3754 2491 3810
rect 2547 3754 2615 3810
rect 2671 3754 2681 3810
rect 2481 3686 2681 3754
rect 2481 3630 2491 3686
rect 2547 3630 2615 3686
rect 2671 3630 2681 3686
rect 2481 3562 2681 3630
rect 2481 3506 2491 3562
rect 2547 3506 2615 3562
rect 2671 3506 2681 3562
rect 2481 3438 2681 3506
rect 2481 3382 2491 3438
rect 2547 3382 2615 3438
rect 2671 3382 2681 3438
rect 2481 3314 2681 3382
rect 2481 3258 2491 3314
rect 2547 3258 2615 3314
rect 2671 3258 2681 3314
rect 2481 3190 2681 3258
rect 2481 3134 2491 3190
rect 2547 3134 2615 3190
rect 2671 3134 2681 3190
rect 2481 3066 2681 3134
rect 2481 3010 2491 3066
rect 2547 3010 2615 3066
rect 2671 3010 2681 3066
rect 2481 2942 2681 3010
rect 2481 2886 2491 2942
rect 2547 2886 2615 2942
rect 2671 2886 2681 2942
rect 2481 2818 2681 2886
rect 2481 2762 2491 2818
rect 2547 2762 2615 2818
rect 2671 2762 2681 2818
rect 2481 2694 2681 2762
rect 2481 2638 2491 2694
rect 2547 2638 2615 2694
rect 2671 2638 2681 2694
rect 2481 2570 2681 2638
rect 2481 2514 2491 2570
rect 2547 2514 2615 2570
rect 2671 2514 2681 2570
rect 2481 2446 2681 2514
rect 2481 2390 2491 2446
rect 2547 2390 2615 2446
rect 2671 2390 2681 2446
rect 2481 2322 2681 2390
rect 2481 2266 2491 2322
rect 2547 2266 2615 2322
rect 2671 2266 2681 2322
rect 2481 2198 2681 2266
rect 2481 2142 2491 2198
rect 2547 2142 2615 2198
rect 2671 2142 2681 2198
rect 2481 2074 2681 2142
rect 2481 2018 2491 2074
rect 2547 2018 2615 2074
rect 2671 2018 2681 2074
rect 2481 1950 2681 2018
rect 2481 1894 2491 1950
rect 2547 1894 2615 1950
rect 2671 1894 2681 1950
rect 2481 1826 2681 1894
rect 2481 1770 2491 1826
rect 2547 1770 2615 1826
rect 2671 1770 2681 1826
rect 2481 1702 2681 1770
rect 2481 1646 2491 1702
rect 2547 1646 2615 1702
rect 2671 1646 2681 1702
rect 2481 1636 2681 1646
rect 4851 4554 5051 4564
rect 4851 4498 4861 4554
rect 4917 4498 4985 4554
rect 5041 4498 5051 4554
rect 4851 4430 5051 4498
rect 4851 4374 4861 4430
rect 4917 4374 4985 4430
rect 5041 4374 5051 4430
rect 4851 4306 5051 4374
rect 4851 4250 4861 4306
rect 4917 4250 4985 4306
rect 5041 4250 5051 4306
rect 4851 4182 5051 4250
rect 4851 4126 4861 4182
rect 4917 4126 4985 4182
rect 5041 4126 5051 4182
rect 4851 4058 5051 4126
rect 4851 4002 4861 4058
rect 4917 4002 4985 4058
rect 5041 4002 5051 4058
rect 4851 3934 5051 4002
rect 4851 3878 4861 3934
rect 4917 3878 4985 3934
rect 5041 3878 5051 3934
rect 4851 3810 5051 3878
rect 4851 3754 4861 3810
rect 4917 3754 4985 3810
rect 5041 3754 5051 3810
rect 4851 3686 5051 3754
rect 4851 3630 4861 3686
rect 4917 3630 4985 3686
rect 5041 3630 5051 3686
rect 4851 3562 5051 3630
rect 4851 3506 4861 3562
rect 4917 3506 4985 3562
rect 5041 3506 5051 3562
rect 4851 3438 5051 3506
rect 4851 3382 4861 3438
rect 4917 3382 4985 3438
rect 5041 3382 5051 3438
rect 4851 3314 5051 3382
rect 4851 3258 4861 3314
rect 4917 3258 4985 3314
rect 5041 3258 5051 3314
rect 4851 3190 5051 3258
rect 4851 3134 4861 3190
rect 4917 3134 4985 3190
rect 5041 3134 5051 3190
rect 4851 3066 5051 3134
rect 4851 3010 4861 3066
rect 4917 3010 4985 3066
rect 5041 3010 5051 3066
rect 4851 2942 5051 3010
rect 4851 2886 4861 2942
rect 4917 2886 4985 2942
rect 5041 2886 5051 2942
rect 4851 2818 5051 2886
rect 4851 2762 4861 2818
rect 4917 2762 4985 2818
rect 5041 2762 5051 2818
rect 4851 2694 5051 2762
rect 4851 2638 4861 2694
rect 4917 2638 4985 2694
rect 5041 2638 5051 2694
rect 4851 2570 5051 2638
rect 4851 2514 4861 2570
rect 4917 2514 4985 2570
rect 5041 2514 5051 2570
rect 4851 2446 5051 2514
rect 4851 2390 4861 2446
rect 4917 2390 4985 2446
rect 5041 2390 5051 2446
rect 4851 2322 5051 2390
rect 4851 2266 4861 2322
rect 4917 2266 4985 2322
rect 5041 2266 5051 2322
rect 4851 2198 5051 2266
rect 4851 2142 4861 2198
rect 4917 2142 4985 2198
rect 5041 2142 5051 2198
rect 4851 2074 5051 2142
rect 4851 2018 4861 2074
rect 4917 2018 4985 2074
rect 5041 2018 5051 2074
rect 4851 1950 5051 2018
rect 4851 1894 4861 1950
rect 4917 1894 4985 1950
rect 5041 1894 5051 1950
rect 4851 1826 5051 1894
rect 4851 1770 4861 1826
rect 4917 1770 4985 1826
rect 5041 1770 5051 1826
rect 4851 1702 5051 1770
rect 4851 1646 4861 1702
rect 4917 1646 4985 1702
rect 5041 1646 5051 1702
rect 4851 1636 5051 1646
rect 7265 4554 7713 4564
rect 7265 4498 7275 4554
rect 7331 4498 7399 4554
rect 7455 4498 7523 4554
rect 7579 4498 7647 4554
rect 7703 4498 7713 4554
rect 7265 4430 7713 4498
rect 7265 4374 7275 4430
rect 7331 4374 7399 4430
rect 7455 4374 7523 4430
rect 7579 4374 7647 4430
rect 7703 4374 7713 4430
rect 7265 4306 7713 4374
rect 7265 4250 7275 4306
rect 7331 4250 7399 4306
rect 7455 4250 7523 4306
rect 7579 4250 7647 4306
rect 7703 4250 7713 4306
rect 7265 4182 7713 4250
rect 7265 4126 7275 4182
rect 7331 4126 7399 4182
rect 7455 4126 7523 4182
rect 7579 4126 7647 4182
rect 7703 4126 7713 4182
rect 7265 4058 7713 4126
rect 7265 4002 7275 4058
rect 7331 4002 7399 4058
rect 7455 4002 7523 4058
rect 7579 4002 7647 4058
rect 7703 4002 7713 4058
rect 7265 3934 7713 4002
rect 7265 3878 7275 3934
rect 7331 3878 7399 3934
rect 7455 3878 7523 3934
rect 7579 3878 7647 3934
rect 7703 3878 7713 3934
rect 7265 3810 7713 3878
rect 7265 3754 7275 3810
rect 7331 3754 7399 3810
rect 7455 3754 7523 3810
rect 7579 3754 7647 3810
rect 7703 3754 7713 3810
rect 7265 3686 7713 3754
rect 7265 3630 7275 3686
rect 7331 3630 7399 3686
rect 7455 3630 7523 3686
rect 7579 3630 7647 3686
rect 7703 3630 7713 3686
rect 7265 3562 7713 3630
rect 7265 3506 7275 3562
rect 7331 3506 7399 3562
rect 7455 3506 7523 3562
rect 7579 3506 7647 3562
rect 7703 3506 7713 3562
rect 7265 3438 7713 3506
rect 7265 3382 7275 3438
rect 7331 3382 7399 3438
rect 7455 3382 7523 3438
rect 7579 3382 7647 3438
rect 7703 3382 7713 3438
rect 7265 3314 7713 3382
rect 7265 3258 7275 3314
rect 7331 3258 7399 3314
rect 7455 3258 7523 3314
rect 7579 3258 7647 3314
rect 7703 3258 7713 3314
rect 7265 3190 7713 3258
rect 7265 3134 7275 3190
rect 7331 3134 7399 3190
rect 7455 3134 7523 3190
rect 7579 3134 7647 3190
rect 7703 3134 7713 3190
rect 7265 3066 7713 3134
rect 7265 3010 7275 3066
rect 7331 3010 7399 3066
rect 7455 3010 7523 3066
rect 7579 3010 7647 3066
rect 7703 3010 7713 3066
rect 7265 2942 7713 3010
rect 7265 2886 7275 2942
rect 7331 2886 7399 2942
rect 7455 2886 7523 2942
rect 7579 2886 7647 2942
rect 7703 2886 7713 2942
rect 7265 2818 7713 2886
rect 7265 2762 7275 2818
rect 7331 2762 7399 2818
rect 7455 2762 7523 2818
rect 7579 2762 7647 2818
rect 7703 2762 7713 2818
rect 7265 2694 7713 2762
rect 7265 2638 7275 2694
rect 7331 2638 7399 2694
rect 7455 2638 7523 2694
rect 7579 2638 7647 2694
rect 7703 2638 7713 2694
rect 7265 2570 7713 2638
rect 7265 2514 7275 2570
rect 7331 2514 7399 2570
rect 7455 2514 7523 2570
rect 7579 2514 7647 2570
rect 7703 2514 7713 2570
rect 7265 2446 7713 2514
rect 7265 2390 7275 2446
rect 7331 2390 7399 2446
rect 7455 2390 7523 2446
rect 7579 2390 7647 2446
rect 7703 2390 7713 2446
rect 7265 2322 7713 2390
rect 7265 2266 7275 2322
rect 7331 2266 7399 2322
rect 7455 2266 7523 2322
rect 7579 2266 7647 2322
rect 7703 2266 7713 2322
rect 7265 2198 7713 2266
rect 7265 2142 7275 2198
rect 7331 2142 7399 2198
rect 7455 2142 7523 2198
rect 7579 2142 7647 2198
rect 7703 2142 7713 2198
rect 7265 2074 7713 2142
rect 7265 2018 7275 2074
rect 7331 2018 7399 2074
rect 7455 2018 7523 2074
rect 7579 2018 7647 2074
rect 7703 2018 7713 2074
rect 7265 1950 7713 2018
rect 7265 1894 7275 1950
rect 7331 1894 7399 1950
rect 7455 1894 7523 1950
rect 7579 1894 7647 1950
rect 7703 1894 7713 1950
rect 7265 1826 7713 1894
rect 7265 1770 7275 1826
rect 7331 1770 7399 1826
rect 7455 1770 7523 1826
rect 7579 1770 7647 1826
rect 7703 1770 7713 1826
rect 7265 1702 7713 1770
rect 7265 1646 7275 1702
rect 7331 1646 7399 1702
rect 7455 1646 7523 1702
rect 7579 1646 7647 1702
rect 7703 1646 7713 1702
rect 7265 1636 7713 1646
rect 9927 4554 10127 4564
rect 9927 4498 9937 4554
rect 9993 4498 10061 4554
rect 10117 4498 10127 4554
rect 9927 4430 10127 4498
rect 9927 4374 9937 4430
rect 9993 4374 10061 4430
rect 10117 4374 10127 4430
rect 9927 4306 10127 4374
rect 9927 4250 9937 4306
rect 9993 4250 10061 4306
rect 10117 4250 10127 4306
rect 9927 4182 10127 4250
rect 9927 4126 9937 4182
rect 9993 4126 10061 4182
rect 10117 4126 10127 4182
rect 9927 4058 10127 4126
rect 9927 4002 9937 4058
rect 9993 4002 10061 4058
rect 10117 4002 10127 4058
rect 9927 3934 10127 4002
rect 9927 3878 9937 3934
rect 9993 3878 10061 3934
rect 10117 3878 10127 3934
rect 9927 3810 10127 3878
rect 9927 3754 9937 3810
rect 9993 3754 10061 3810
rect 10117 3754 10127 3810
rect 9927 3686 10127 3754
rect 9927 3630 9937 3686
rect 9993 3630 10061 3686
rect 10117 3630 10127 3686
rect 9927 3562 10127 3630
rect 9927 3506 9937 3562
rect 9993 3506 10061 3562
rect 10117 3506 10127 3562
rect 9927 3438 10127 3506
rect 9927 3382 9937 3438
rect 9993 3382 10061 3438
rect 10117 3382 10127 3438
rect 9927 3314 10127 3382
rect 9927 3258 9937 3314
rect 9993 3258 10061 3314
rect 10117 3258 10127 3314
rect 9927 3190 10127 3258
rect 9927 3134 9937 3190
rect 9993 3134 10061 3190
rect 10117 3134 10127 3190
rect 9927 3066 10127 3134
rect 9927 3010 9937 3066
rect 9993 3010 10061 3066
rect 10117 3010 10127 3066
rect 9927 2942 10127 3010
rect 9927 2886 9937 2942
rect 9993 2886 10061 2942
rect 10117 2886 10127 2942
rect 9927 2818 10127 2886
rect 9927 2762 9937 2818
rect 9993 2762 10061 2818
rect 10117 2762 10127 2818
rect 9927 2694 10127 2762
rect 9927 2638 9937 2694
rect 9993 2638 10061 2694
rect 10117 2638 10127 2694
rect 9927 2570 10127 2638
rect 9927 2514 9937 2570
rect 9993 2514 10061 2570
rect 10117 2514 10127 2570
rect 9927 2446 10127 2514
rect 9927 2390 9937 2446
rect 9993 2390 10061 2446
rect 10117 2390 10127 2446
rect 9927 2322 10127 2390
rect 9927 2266 9937 2322
rect 9993 2266 10061 2322
rect 10117 2266 10127 2322
rect 9927 2198 10127 2266
rect 9927 2142 9937 2198
rect 9993 2142 10061 2198
rect 10117 2142 10127 2198
rect 9927 2074 10127 2142
rect 9927 2018 9937 2074
rect 9993 2018 10061 2074
rect 10117 2018 10127 2074
rect 9927 1950 10127 2018
rect 9927 1894 9937 1950
rect 9993 1894 10061 1950
rect 10117 1894 10127 1950
rect 9927 1826 10127 1894
rect 9927 1770 9937 1826
rect 9993 1770 10061 1826
rect 10117 1770 10127 1826
rect 9927 1702 10127 1770
rect 9927 1646 9937 1702
rect 9993 1646 10061 1702
rect 10117 1646 10127 1702
rect 9927 1636 10127 1646
rect 12297 4554 12497 4564
rect 12297 4498 12307 4554
rect 12363 4498 12431 4554
rect 12487 4498 12497 4554
rect 12297 4430 12497 4498
rect 12297 4374 12307 4430
rect 12363 4374 12431 4430
rect 12487 4374 12497 4430
rect 12297 4306 12497 4374
rect 12297 4250 12307 4306
rect 12363 4250 12431 4306
rect 12487 4250 12497 4306
rect 12297 4182 12497 4250
rect 12297 4126 12307 4182
rect 12363 4126 12431 4182
rect 12487 4126 12497 4182
rect 12297 4058 12497 4126
rect 12297 4002 12307 4058
rect 12363 4002 12431 4058
rect 12487 4002 12497 4058
rect 12297 3934 12497 4002
rect 12297 3878 12307 3934
rect 12363 3878 12431 3934
rect 12487 3878 12497 3934
rect 12297 3810 12497 3878
rect 12297 3754 12307 3810
rect 12363 3754 12431 3810
rect 12487 3754 12497 3810
rect 12297 3686 12497 3754
rect 12297 3630 12307 3686
rect 12363 3630 12431 3686
rect 12487 3630 12497 3686
rect 12297 3562 12497 3630
rect 12297 3506 12307 3562
rect 12363 3506 12431 3562
rect 12487 3506 12497 3562
rect 12297 3438 12497 3506
rect 12297 3382 12307 3438
rect 12363 3382 12431 3438
rect 12487 3382 12497 3438
rect 12297 3314 12497 3382
rect 12297 3258 12307 3314
rect 12363 3258 12431 3314
rect 12487 3258 12497 3314
rect 12297 3190 12497 3258
rect 12297 3134 12307 3190
rect 12363 3134 12431 3190
rect 12487 3134 12497 3190
rect 12297 3066 12497 3134
rect 12297 3010 12307 3066
rect 12363 3010 12431 3066
rect 12487 3010 12497 3066
rect 12297 2942 12497 3010
rect 12297 2886 12307 2942
rect 12363 2886 12431 2942
rect 12487 2886 12497 2942
rect 12297 2818 12497 2886
rect 12297 2762 12307 2818
rect 12363 2762 12431 2818
rect 12487 2762 12497 2818
rect 12297 2694 12497 2762
rect 12297 2638 12307 2694
rect 12363 2638 12431 2694
rect 12487 2638 12497 2694
rect 12297 2570 12497 2638
rect 12297 2514 12307 2570
rect 12363 2514 12431 2570
rect 12487 2514 12497 2570
rect 12297 2446 12497 2514
rect 12297 2390 12307 2446
rect 12363 2390 12431 2446
rect 12487 2390 12497 2446
rect 12297 2322 12497 2390
rect 12297 2266 12307 2322
rect 12363 2266 12431 2322
rect 12487 2266 12497 2322
rect 12297 2198 12497 2266
rect 12297 2142 12307 2198
rect 12363 2142 12431 2198
rect 12487 2142 12497 2198
rect 12297 2074 12497 2142
rect 12297 2018 12307 2074
rect 12363 2018 12431 2074
rect 12487 2018 12497 2074
rect 12297 1950 12497 2018
rect 12297 1894 12307 1950
rect 12363 1894 12431 1950
rect 12487 1894 12497 1950
rect 12297 1826 12497 1894
rect 12297 1770 12307 1826
rect 12363 1770 12431 1826
rect 12487 1770 12497 1826
rect 12297 1702 12497 1770
rect 12297 1646 12307 1702
rect 12363 1646 12431 1702
rect 12487 1646 12497 1702
rect 12297 1636 12497 1646
use comp018green_esd_clamp_v5p0_DVDD  comp018green_esd_clamp_v5p0_DVDD_0
timestamp 1698431365
transform 1 0 1008 0 1 1147
box -747 -51 13709 46134
use M1_NWELL_CDNS_4066195314571  M1_NWELL_CDNS_4066195314571_0
timestamp 1698431365
transform 1 0 2735 0 1 50138
box 0 0 1 1
use M1_NWELL_CDNS_4066195314571  M1_NWELL_CDNS_4066195314571_1
timestamp 1698431365
transform 1 0 12243 0 1 50138
box 0 0 1 1
use M1_NWELL_CDNS_4066195314572  M1_NWELL_CDNS_4066195314572_0
timestamp 1698431365
transform 1 0 7489 0 1 52438
box 0 0 1 1
use M1_NWELL_CDNS_4066195314572  M1_NWELL_CDNS_4066195314572_1
timestamp 1698431365
transform 1 0 7489 0 1 47838
box 0 0 1 1
use M1_PSUB_CDNS_4066195314564  M1_PSUB_CDNS_4066195314564_0
timestamp 1698431365
transform 1 0 379 0 1 55155
box 0 0 1 1
use M1_PSUB_CDNS_4066195314564  M1_PSUB_CDNS_4066195314564_1
timestamp 1698431365
transform 1 0 14599 0 1 55155
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_0
timestamp 1698431365
transform 1 0 7489 0 1 53228
box 0 0 1 1
use M1_PSUB_CDNS_4066195314565  M1_PSUB_CDNS_4066195314565_1
timestamp 1698431365
transform 1 0 7489 0 1 57082
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_0
timestamp 1698431365
transform 1 0 3293 0 1 51539
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_1
timestamp 1698431365
transform 1 0 3293 0 1 50605
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_2
timestamp 1698431365
transform 1 0 3293 0 1 49671
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_3
timestamp 1698431365
transform 1 0 3293 0 1 48737
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_4
timestamp 1698431365
transform -1 0 11685 0 1 51539
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_5
timestamp 1698431365
transform -1 0 11685 0 1 50605
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_6
timestamp 1698431365
transform -1 0 11685 0 1 48737
box 0 0 1 1
use M1_PSUB_CDNS_4066195314566  M1_PSUB_CDNS_4066195314566_7
timestamp 1698431365
transform -1 0 11685 0 1 49671
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_0
timestamp 1698431365
transform 1 0 7489 0 -1 51852
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_1
timestamp 1698431365
transform 1 0 7489 0 1 49050
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_2
timestamp 1698431365
transform 1 0 7489 0 1 49358
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_3
timestamp 1698431365
transform 1 0 7489 0 1 49984
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_4
timestamp 1698431365
transform 1 0 7489 0 1 50292
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_5
timestamp 1698431365
transform 1 0 7489 0 1 50918
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_6
timestamp 1698431365
transform 1 0 7489 0 1 51226
box 0 0 1 1
use M1_PSUB_CDNS_4066195314567  M1_PSUB_CDNS_4066195314567_7
timestamp 1698431365
transform 1 0 7489 0 1 48424
box 0 0 1 1
use M1_PSUB_CDNS_4066195314568  M1_PSUB_CDNS_4066195314568_0
timestamp 1698431365
transform 1 0 7489 0 1 51072
box 0 0 1 1
use M1_PSUB_CDNS_4066195314568  M1_PSUB_CDNS_4066195314568_1
timestamp 1698431365
transform 1 0 7489 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_4066195314568  M1_PSUB_CDNS_4066195314568_2
timestamp 1698431365
transform 1 0 7489 0 1 49204
box 0 0 1 1
use M1_PSUB_CDNS_4066195314569  M1_PSUB_CDNS_4066195314569_0
timestamp 1698431365
transform 1 0 7489 0 -1 52006
box 0 0 1 1
use M1_PSUB_CDNS_4066195314569  M1_PSUB_CDNS_4066195314569_1
timestamp 1698431365
transform 1 0 7489 0 1 48270
box 0 0 1 1
use M1_PSUB_CDNS_4066195314570  M1_PSUB_CDNS_4066195314570_0
timestamp 1698431365
transform 1 0 3139 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_4066195314570  M1_PSUB_CDNS_4066195314570_1
timestamp 1698431365
transform -1 0 11839 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_4066195314599  M1_PSUB_CDNS_4066195314599_0
timestamp 1698431365
transform 1 0 13496 0 1 34924
box 0 0 1 1
use M1_PSUB_CDNS_40661953145100  M1_PSUB_CDNS_40661953145100_0
timestamp 1698431365
transform 1 0 14487 0 1 21924
box 0 0 1 1
use M1_PSUB_CDNS_40661953145100  M1_PSUB_CDNS_40661953145100_1
timestamp 1698431365
transform 1 0 491 0 1 21924
box 0 0 1 1
use M1_PSUB_CDNS_40661953145101  M1_PSUB_CDNS_40661953145101_0
timestamp 1698431365
transform 1 0 1241 0 1 50138
box 0 0 1 1
use M1_PSUB_CDNS_40661953145101  M1_PSUB_CDNS_40661953145101_1
timestamp 1698431365
transform 1 0 13737 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_0
timestamp 1698431365
transform 1 0 2581 0 1 53350
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_1
timestamp 1698431365
transform 1 0 4951 0 1 53350
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_2
timestamp 1698431365
transform 1 0 12397 0 1 53350
box 0 0 1 1
use M2_M1_CDNS_4066195314573  M2_M1_CDNS_4066195314573_3
timestamp 1698431365
transform 1 0 10027 0 1 53350
box 0 0 1 1
use M2_M1_CDNS_4066195314574  M2_M1_CDNS_4066195314574_0
timestamp 1698431365
transform 1 0 7489 0 1 53350
box 0 0 1 1
use M2_M1_CDNS_4066195314575  M2_M1_CDNS_4066195314575_0
timestamp 1698431365
transform 1 0 6695 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314575  M2_M1_CDNS_4066195314575_1
timestamp 1698431365
transform 1 0 8283 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314576  M2_M1_CDNS_4066195314576_0
timestamp 1698431365
transform 1 0 4951 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_4066195314576  M2_M1_CDNS_4066195314576_1
timestamp 1698431365
transform 1 0 4951 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_4066195314576  M2_M1_CDNS_4066195314576_2
timestamp 1698431365
transform -1 0 10027 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_4066195314576  M2_M1_CDNS_4066195314576_3
timestamp 1698431365
transform -1 0 10027 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_0
timestamp 1698431365
transform 1 0 3766 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_1
timestamp 1698431365
transform 1 0 3766 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_2
timestamp 1698431365
transform 1 0 6136 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_3
timestamp 1698431365
transform 1 0 6136 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_4
timestamp 1698431365
transform -1 0 8842 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_5
timestamp 1698431365
transform -1 0 8842 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_6
timestamp 1698431365
transform -1 0 11212 0 1 47838
box 0 0 1 1
use M2_M1_CDNS_4066195314577  M2_M1_CDNS_4066195314577_7
timestamp 1698431365
transform -1 0 11212 0 1 52438
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_0
timestamp 1698431365
transform 1 0 4143 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_1
timestamp 1698431365
transform 1 0 4143 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_2
timestamp 1698431365
transform 1 0 4143 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_3
timestamp 1698431365
transform 1 0 4143 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_4
timestamp 1698431365
transform -1 0 10835 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_5
timestamp 1698431365
transform -1 0 10835 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_6
timestamp 1698431365
transform -1 0 10835 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_4066195314578  M2_M1_CDNS_4066195314578_7
timestamp 1698431365
transform -1 0 10835 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_0
timestamp 1698431365
transform 1 0 6136 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_1
timestamp 1698431365
transform 1 0 6136 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_2
timestamp 1698431365
transform 1 0 6136 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_3
timestamp 1698431365
transform 1 0 6136 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_4
timestamp 1698431365
transform -1 0 8842 0 1 50605
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_5
timestamp 1698431365
transform -1 0 8842 0 1 48737
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_6
timestamp 1698431365
transform -1 0 8842 0 1 49671
box 0 0 1 1
use M2_M1_CDNS_4066195314579  M2_M1_CDNS_4066195314579_7
timestamp 1698431365
transform -1 0 8842 0 1 51539
box 0 0 1 1
use M2_M1_CDNS_4066195314580  M2_M1_CDNS_4066195314580_0
timestamp 1698431365
transform 1 0 4552 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314580  M2_M1_CDNS_4066195314580_1
timestamp 1698431365
transform 1 0 10426 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314581  M2_M1_CDNS_4066195314581_0
timestamp 1698431365
transform 1 0 3293 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314581  M2_M1_CDNS_4066195314581_1
timestamp 1698431365
transform 1 0 1377 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314581  M2_M1_CDNS_4066195314581_2
timestamp 1698431365
transform -1 0 11685 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314581  M2_M1_CDNS_4066195314581_3
timestamp 1698431365
transform -1 0 13601 0 1 55155
box 0 0 1 1
use M2_M1_CDNS_4066195314582  M2_M1_CDNS_4066195314582_0
timestamp 1698431365
transform -1 0 7489 0 1 48347
box 0 0 1 1
use M2_M1_CDNS_4066195314582  M2_M1_CDNS_4066195314582_1
timestamp 1698431365
transform -1 0 7489 0 1 51929
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_0
timestamp 1698431365
transform 1 0 4951 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_1
timestamp 1698431365
transform 1 0 4951 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_2
timestamp 1698431365
transform 1 0 4951 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_3
timestamp 1698431365
transform -1 0 10027 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_4
timestamp 1698431365
transform -1 0 10027 0 1 51072
box 0 0 1 1
use M2_M1_CDNS_4066195314583  M2_M1_CDNS_4066195314583_5
timestamp 1698431365
transform -1 0 10027 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_4066195314585  M2_M1_CDNS_4066195314585_0
timestamp 1698431365
transform 1 0 7489 0 1 57082
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_0
timestamp 1698431365
transform 1 0 4951 0 1 57082
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_1
timestamp 1698431365
transform 1 0 2581 0 1 57082
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_2
timestamp 1698431365
transform 1 0 10027 0 1 57082
box 0 0 1 1
use M2_M1_CDNS_4066195314586  M2_M1_CDNS_4066195314586_3
timestamp 1698431365
transform 1 0 12397 0 1 57082
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_0
timestamp 1698431365
transform 1 0 48 0 1 37500
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_1
timestamp 1698431365
transform 1 0 48 0 1 51900
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_2
timestamp 1698431365
transform 1 0 14930 0 1 37500
box 0 0 1 1
use M2_M1_CDNS_4066195314588  M2_M1_CDNS_4066195314588_3
timestamp 1698431365
transform 1 0 14930 0 1 51900
box 0 0 1 1
use M2_M1_CDNS_4066195314591  M2_M1_CDNS_4066195314591_0
timestamp 1698431365
transform -1 0 7489 0 1 50138
box 0 0 1 1
use M2_M1_CDNS_4066195314591  M2_M1_CDNS_4066195314591_1
timestamp 1698431365
transform -1 0 7489 0 1 49204
box 0 0 1 1
use M2_M1_CDNS_4066195314591  M2_M1_CDNS_4066195314591_2
timestamp 1698431365
transform -1 0 7489 0 1 51072
box 0 0 1 1
use M3_M2_CDNS_406619531456  M3_M2_CDNS_406619531456_0
timestamp 1698431365
transform 1 0 2581 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_406619531456  M3_M2_CDNS_406619531456_1
timestamp 1698431365
transform 1 0 4951 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_406619531456  M3_M2_CDNS_406619531456_2
timestamp 1698431365
transform 1 0 12397 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_406619531456  M3_M2_CDNS_406619531456_3
timestamp 1698431365
transform 1 0 10027 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_0
timestamp 1698431365
transform 1 0 13767 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_1
timestamp 1698431365
transform 1 0 13767 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_2
timestamp 1698431365
transform 1 0 13767 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_3
timestamp 1698431365
transform 1 0 13767 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_4
timestamp 1698431365
transform 1 0 1211 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_5
timestamp 1698431365
transform 1 0 1211 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_6
timestamp 1698431365
transform 1 0 1211 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_7
timestamp 1698431365
transform 1 0 1211 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_8
timestamp 1698431365
transform 1 0 1211 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314584  M3_M2_CDNS_4066195314584_9
timestamp 1698431365
transform 1 0 13767 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_0
timestamp 1698431365
transform 1 0 48 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_1
timestamp 1698431365
transform 1 0 48 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_2
timestamp 1698431365
transform 1 0 14930 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_4066195314587  M3_M2_CDNS_4066195314587_3
timestamp 1698431365
transform 1 0 14930 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_4066195314589  M3_M2_CDNS_4066195314589_0
timestamp 1698431365
transform 1 0 2317 0 1 37513
box 0 0 1 1
use M3_M2_CDNS_4066195314589  M3_M2_CDNS_4066195314589_1
timestamp 1698431365
transform 1 0 2317 0 1 51899
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_0
timestamp 1698431365
transform 1 0 13767 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_1
timestamp 1698431365
transform 1 0 1211 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_2
timestamp 1698431365
transform 1 0 1211 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_3
timestamp 1698431365
transform 1 0 1211 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_4
timestamp 1698431365
transform 1 0 1211 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_5
timestamp 1698431365
transform 1 0 1211 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_6
timestamp 1698431365
transform 1 0 1211 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_7
timestamp 1698431365
transform 1 0 1211 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_8
timestamp 1698431365
transform 1 0 1211 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_9
timestamp 1698431365
transform 1 0 13767 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_10
timestamp 1698431365
transform 1 0 13767 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_11
timestamp 1698431365
transform 1 0 13767 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_12
timestamp 1698431365
transform 1 0 13767 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_13
timestamp 1698431365
transform 1 0 13767 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_14
timestamp 1698431365
transform 1 0 13767 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_15
timestamp 1698431365
transform 1 0 13767 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_16
timestamp 1698431365
transform 1 0 1211 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314590  M3_M2_CDNS_4066195314590_17
timestamp 1698431365
transform 1 0 13767 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_0
timestamp 1698431365
transform 1 0 11212 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_1
timestamp 1698431365
transform 1 0 8842 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_2
timestamp 1698431365
transform 1 0 6136 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_3
timestamp 1698431365
transform 1 0 3766 0 1 11900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_4
timestamp 1698431365
transform 1 0 6136 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_5
timestamp 1698431365
transform 1 0 6136 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_6
timestamp 1698431365
transform 1 0 6136 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_7
timestamp 1698431365
transform 1 0 6136 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_8
timestamp 1698431365
transform 1 0 6136 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_9
timestamp 1698431365
transform 1 0 3766 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_10
timestamp 1698431365
transform 1 0 3766 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_11
timestamp 1698431365
transform 1 0 3766 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_12
timestamp 1698431365
transform 1 0 3766 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_13
timestamp 1698431365
transform 1 0 3766 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_14
timestamp 1698431365
transform 1 0 3766 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_15
timestamp 1698431365
transform 1 0 3766 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_16
timestamp 1698431365
transform 1 0 6136 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_17
timestamp 1698431365
transform 1 0 6136 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_18
timestamp 1698431365
transform 1 0 8842 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_19
timestamp 1698431365
transform 1 0 8842 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_20
timestamp 1698431365
transform 1 0 8842 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_21
timestamp 1698431365
transform 1 0 8842 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_22
timestamp 1698431365
transform 1 0 8842 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_23
timestamp 1698431365
transform 1 0 8842 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_24
timestamp 1698431365
transform 1 0 11212 0 1 50300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_25
timestamp 1698431365
transform 1 0 11212 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_26
timestamp 1698431365
transform 1 0 11212 0 1 39100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_27
timestamp 1698431365
transform 1 0 11212 0 1 40700
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_28
timestamp 1698431365
transform 1 0 11212 0 1 42300
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_29
timestamp 1698431365
transform 1 0 11212 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_30
timestamp 1698431365
transform 1 0 11212 0 1 47100
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_31
timestamp 1698431365
transform 1 0 8842 0 1 43900
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_32
timestamp 1698431365
transform 1 0 6136 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_33
timestamp 1698431365
transform 1 0 8842 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_34
timestamp 1698431365
transform 1 0 3766 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314592  M3_M2_CDNS_4066195314592_35
timestamp 1698431365
transform 1 0 11212 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_0
timestamp 1698431365
transform 1 0 11212 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_1
timestamp 1698431365
transform 1 0 11212 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_2
timestamp 1698431365
transform 1 0 8842 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_3
timestamp 1698431365
transform 1 0 8842 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_4
timestamp 1698431365
transform 1 0 11212 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_5
timestamp 1698431365
transform 1 0 8842 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_6
timestamp 1698431365
transform 1 0 8842 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_7
timestamp 1698431365
transform 1 0 11212 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_8
timestamp 1698431365
transform 1 0 3766 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_9
timestamp 1698431365
transform 1 0 3766 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_10
timestamp 1698431365
transform 1 0 3766 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_11
timestamp 1698431365
transform 1 0 3766 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_12
timestamp 1698431365
transform 1 0 6136 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_13
timestamp 1698431365
transform 1 0 6136 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_14
timestamp 1698431365
transform 1 0 6136 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_15
timestamp 1698431365
transform 1 0 6136 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_16
timestamp 1698431365
transform 1 0 6136 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_17
timestamp 1698431365
transform 1 0 3766 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_18
timestamp 1698431365
transform 1 0 8842 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314593  M3_M2_CDNS_4066195314593_19
timestamp 1698431365
transform 1 0 11212 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_0
timestamp 1698431365
transform 1 0 12397 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_1
timestamp 1698431365
transform 1 0 10027 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_2
timestamp 1698431365
transform 1 0 12397 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_3
timestamp 1698431365
transform 1 0 10027 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_4
timestamp 1698431365
transform 1 0 2581 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_5
timestamp 1698431365
transform 1 0 4951 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_6
timestamp 1698431365
transform 1 0 2581 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_7
timestamp 1698431365
transform 1 0 4951 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_8
timestamp 1698431365
transform 1 0 2581 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_9
timestamp 1698431365
transform 1 0 2581 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_10
timestamp 1698431365
transform 1 0 4951 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_11
timestamp 1698431365
transform 1 0 2581 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_12
timestamp 1698431365
transform 1 0 4951 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_13
timestamp 1698431365
transform 1 0 4951 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_14
timestamp 1698431365
transform 1 0 10027 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_15
timestamp 1698431365
transform 1 0 10027 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_16
timestamp 1698431365
transform 1 0 12397 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_17
timestamp 1698431365
transform 1 0 10027 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_18
timestamp 1698431365
transform 1 0 12397 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_4066195314594  M3_M2_CDNS_4066195314594_19
timestamp 1698431365
transform 1 0 12397 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_4066195314595  M3_M2_CDNS_4066195314595_0
timestamp 1698431365
transform 1 0 7489 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_0
timestamp 1698431365
transform 1 0 7489 0 1 53500
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_1
timestamp 1698431365
transform 1 0 7489 0 1 48700
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_2
timestamp 1698431365
transform 1 0 7489 0 1 45500
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_3
timestamp 1698431365
transform 1 0 7489 0 1 13500
box 0 0 1 1
use M3_M2_CDNS_4066195314596  M3_M2_CDNS_4066195314596_4
timestamp 1698431365
transform 1 0 7489 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_0
timestamp 1698431365
transform 1 0 12397 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_1
timestamp 1698431365
transform 1 0 10027 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_2
timestamp 1698431365
transform 1 0 10027 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_3
timestamp 1698431365
transform 1 0 12397 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_4
timestamp 1698431365
transform 1 0 10027 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_5
timestamp 1698431365
transform 1 0 12397 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_6
timestamp 1698431365
transform 1 0 4951 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_7
timestamp 1698431365
transform 1 0 2581 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_8
timestamp 1698431365
transform 1 0 4951 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_9
timestamp 1698431365
transform 1 0 2581 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_10
timestamp 1698431365
transform 1 0 4951 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_11
timestamp 1698431365
transform 1 0 2581 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_12
timestamp 1698431365
transform 1 0 4951 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_13
timestamp 1698431365
transform 1 0 2581 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_14
timestamp 1698431365
transform 1 0 10027 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_4066195314597  M3_M2_CDNS_4066195314597_15
timestamp 1698431365
transform 1 0 12397 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_0
timestamp 1698431365
transform 1 0 7489 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_1
timestamp 1698431365
transform 1 0 7489 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_2
timestamp 1698431365
transform 1 0 7489 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_4066195314598  M3_M2_CDNS_4066195314598_3
timestamp 1698431365
transform 1 0 7489 0 1 35100
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_0
timestamp 1698431365
transform 1 0 835 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_1
timestamp 1698431365
transform 1 0 11143 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_2
timestamp 1698431365
transform 1 0 7707 0 1 53655
box 0 0 1 1
use nmoscap_6p0_CDNS_406619531450  nmoscap_6p0_CDNS_406619531450_3
timestamp 1698431365
transform 1 0 4271 0 1 53655
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_0
timestamp 1698431365
transform 1 0 3489 0 1 51439
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_1
timestamp 1698431365
transform 1 0 3489 0 1 50505
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_2
timestamp 1698431365
transform 1 0 3489 0 1 49571
box 0 0 1 1
use np_6p0_CDNS_406619531451  np_6p0_CDNS_406619531451_3
timestamp 1698431365
transform 1 0 3489 0 1 48637
box 0 0 1 1
<< labels >>
rlabel metal3 s 705 6432 705 6432 4 DVSS
port 1 nsew
rlabel metal3 s 752 3261 752 3261 4 DVSS
port 1 nsew
rlabel metal3 s 774 9418 774 9418 4 DVSS
port 1 nsew
rlabel metal3 s 774 13611 774 13611 4 DVSS
port 1 nsew
rlabel metal3 s 774 11795 774 11795 4 DVDD
port 2 nsew
rlabel metal3 s 774 22234 774 22234 4 DVDD
port 2 nsew
rlabel metal3 s 774 19120 774 19120 4 DVDD
port 2 nsew
rlabel metal3 s 774 15905 774 15905 4 DVDD
port 2 nsew
rlabel metal3 s 774 27853 774 27853 4 DVSS
port 1 nsew
rlabel metal3 s 774 29488 774 29488 4 DVDD
port 2 nsew
rlabel metal3 s 774 25470 774 25470 4 DVDD
port 2 nsew
rlabel metal3 s 774 35106 774 35106 4 DVSS
port 1 nsew
rlabel metal3 s 774 31879 774 31879 4 DVDD
port 2 nsew
rlabel metal3 s 774 45369 774 45369 4 DVSS
port 1 nsew
rlabel metal3 s 774 43934 774 43934 4 DVDD
port 2 nsew
rlabel metal3 s 774 42169 774 42169 4 DVDD
port 2 nsew
rlabel metal3 s 774 40734 774 40734 4 DVDD
port 2 nsew
rlabel metal3 s 774 48569 774 48569 4 DVSS
port 1 nsew
rlabel metal3 s 774 53534 774 53534 4 DVSS
port 1 nsew
rlabel metal3 s 774 56560 774 56560 4 DVSS
port 1 nsew
rlabel metal3 s 774 54969 774 54969 4 DVDD
port 2 nsew
rlabel metal3 s 774 47134 774 47134 4 DVDD
port 2 nsew
<< properties >>
string GDS_END 4779612
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4757140
string path 344.175 29.750 344.175 0.000 
<< end >>
