magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
use pmos_5p04310590878118_256x8m81  pmos_5p04310590878118_256x8m81_0
timestamp 1698431365
transform 1 0 -31 0 1 0
box 0 0 1 1
<< properties >>
string GDS_END 310132
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 309178
<< end >>
