magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 124 74 244 206
rect 348 74 468 206
rect 572 74 692 206
rect 796 74 916 206
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 796 573 896 939
<< mvndiff >>
rect 36 190 124 206
rect 36 144 49 190
rect 95 144 124 190
rect 36 74 124 144
rect 244 193 348 206
rect 244 147 273 193
rect 319 147 348 193
rect 244 74 348 147
rect 468 185 572 206
rect 468 139 497 185
rect 543 139 572 185
rect 468 74 572 139
rect 692 193 796 206
rect 692 147 721 193
rect 767 147 796 193
rect 692 74 796 147
rect 916 190 1004 206
rect 916 144 945 190
rect 991 144 1004 190
rect 916 74 1004 144
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 573 582 939
rect 682 573 796 939
rect 896 861 984 939
rect 896 721 925 861
rect 971 721 984 861
rect 896 573 984 721
<< mvndiffc >>
rect 49 144 95 190
rect 273 147 319 193
rect 497 139 543 185
rect 721 147 767 193
rect 945 144 991 190
<< mvpdiffc >>
rect 69 721 115 861
rect 925 721 971 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 796 939 896 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 250 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 250 458 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 250 682 454
rect 796 500 896 573
rect 796 454 814 500
rect 860 454 896 500
rect 796 250 896 454
rect 124 206 244 250
rect 348 206 468 250
rect 572 206 692 250
rect 796 206 916 250
rect 124 30 244 74
rect 348 30 468 74
rect 572 30 692 74
rect 796 30 916 74
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 595 454 641 500
rect 814 454 860 500
<< metal1 >>
rect 0 918 1120 1098
rect 69 861 115 918
rect 69 710 115 721
rect 925 861 971 872
rect 925 603 971 721
rect 702 557 971 603
rect 142 500 203 542
rect 142 454 157 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 584 500 652 542
rect 584 454 595 500
rect 641 454 652 500
rect 142 443 203 454
rect 702 288 767 557
rect 814 500 866 511
rect 860 454 866 500
rect 814 354 866 454
rect 273 242 767 288
rect 49 190 95 201
rect 49 90 95 144
rect 273 193 319 242
rect 273 136 319 147
rect 497 185 543 196
rect 497 90 543 139
rect 721 193 767 242
rect 721 136 767 147
rect 945 190 991 201
rect 945 90 991 144
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 814 354 866 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 584 454 652 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 142 443 203 542 0 FreeSans 200 0 0 0 A4
port 4 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 945 196 991 201 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 925 603 971 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 702 557 971 603 1 ZN
port 5 nsew default output
rlabel metal1 s 702 288 767 557 1 ZN
port 5 nsew default output
rlabel metal1 s 273 242 767 288 1 ZN
port 5 nsew default output
rlabel metal1 s 721 136 767 242 1 ZN
port 5 nsew default output
rlabel metal1 s 273 136 319 242 1 ZN
port 5 nsew default output
rlabel metal1 s 69 710 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 49 196 95 201 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 196 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 196 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 196 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 101836
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 98524
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
