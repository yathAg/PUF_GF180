************************************************************************
* auCdl Netlist:
* 
* Library Name:  TCG_Library
* Top Cell Name: npolyf_u
* View Name:     schematic
* Netlisted on:  Nov 24 09:35:58 2021
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM

*.GLOBAL gnd!

*.PIN gnd!

************************************************************************
* Library Name: TCG_Library
* Cell Name:    npolyf_u
* View Name:    schematic
************************************************************************

.SUBCKT npolyf_u I1_0_0_0_0_0_0_R0_MINUS I1_0_0_0_0_0_0_R0_PLUS 
+ I1_0_0_0_1_0_0_R0_MINUS I1_0_0_0_1_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS 
+ I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS I1_0_0_1_1_0_0_R0_PLUS 
+ I1_0_0_2_0_0_0_R0_MINUS I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS 
+ I1_0_0_2_1_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS I1_0_1_0_0_0_0_R0_PLUS 
+ I1_0_1_0_1_0_0_R0_MINUS I1_0_1_0_1_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS 
+ I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS I1_0_1_1_1_0_0_R0_PLUS 
+ I1_0_1_2_0_0_0_R0_MINUS I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS 
+ I1_0_1_2_1_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS I1_0_2_0_0_0_0_R0_PLUS 
+ I1_0_2_0_1_0_0_R0_MINUS I1_0_2_0_1_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS 
+ I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS I1_0_2_1_1_0_0_R0_PLUS 
+ I1_0_2_2_0_0_0_R0_MINUS I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS 
+ I1_0_2_2_1_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS I1_1_0_0_0_0_0_R0_PLUS 
+ I1_1_0_0_1_0_0_R0_MINUS I1_1_0_0_1_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS 
+ I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS I1_1_0_1_1_0_0_R0_PLUS 
+ I1_1_0_2_0_0_0_R0_MINUS I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS 
+ I1_1_0_2_1_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS I1_1_1_0_0_0_0_R0_PLUS 
+ I1_1_1_0_1_0_0_R0_MINUS I1_1_1_0_1_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS 
+ I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS I1_1_1_1_1_0_0_R0_PLUS 
+ I1_1_1_2_0_0_0_R0_MINUS I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS 
+ I1_1_1_2_1_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS I1_1_2_0_0_0_0_R0_PLUS 
+ I1_1_2_0_1_0_0_R0_MINUS I1_1_2_0_1_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS 
+ I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS I1_1_2_1_1_0_0_R0_PLUS 
+ I1_1_2_2_0_0_0_R0_MINUS I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS 
+ I1_1_2_2_1_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS I1_2_0_0_0_0_0_R0_PLUS 
+ I1_2_0_0_1_0_0_R0_MINUS I1_2_0_0_1_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS 
+ I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS I1_2_0_1_1_0_0_R0_PLUS 
+ I1_2_0_2_0_0_0_R0_MINUS I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS 
+ I1_2_0_2_1_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS I1_2_1_0_0_0_0_R0_PLUS 
+ I1_2_1_0_1_0_0_R0_MINUS I1_2_1_0_1_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS 
+ I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS I1_2_1_1_1_0_0_R0_PLUS 
+ I1_2_1_2_0_0_0_R0_MINUS I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS 
+ I1_2_1_2_1_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS I1_2_2_0_0_0_0_R0_PLUS 
+ I1_2_2_0_1_0_0_R0_MINUS I1_2_2_0_1_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS 
+ I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS I1_2_2_1_1_0_0_R0_PLUS 
+ I1_2_2_2_0_0_0_R0_MINUS I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS 
+ I1_2_2_2_1_0_0_R0_PLUS I1_default_MINUS I1_default_PLUS gnd!
*.PININFO I1_0_0_0_0_0_0_R0_MINUS:I I1_0_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_0_1_0_0_R0_MINUS:I I1_0_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_0_0_0_R0_MINUS:I I1_0_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_1_1_0_0_R0_MINUS:I I1_0_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_0_0_0_R0_MINUS:I I1_0_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_0_2_1_0_0_R0_MINUS:I I1_0_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_0_0_0_R0_MINUS:I I1_0_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_0_1_0_0_R0_MINUS:I I1_0_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_0_0_0_R0_MINUS:I I1_0_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_1_1_0_0_R0_MINUS:I I1_0_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_0_0_0_R0_MINUS:I I1_0_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_1_2_1_0_0_R0_MINUS:I I1_0_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_0_0_0_R0_MINUS:I I1_0_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_0_1_0_0_R0_MINUS:I I1_0_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_0_0_0_R0_MINUS:I I1_0_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_1_1_0_0_R0_MINUS:I I1_0_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_0_0_0_R0_MINUS:I I1_0_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_0_2_2_1_0_0_R0_MINUS:I I1_0_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_0_0_0_R0_MINUS:I I1_1_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_0_1_0_0_R0_MINUS:I I1_1_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_0_0_0_R0_MINUS:I I1_1_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_1_1_0_0_R0_MINUS:I I1_1_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_0_0_0_R0_MINUS:I I1_1_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_0_2_1_0_0_R0_MINUS:I I1_1_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_0_0_0_R0_MINUS:I I1_1_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_0_1_0_0_R0_MINUS:I I1_1_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_0_0_0_R0_MINUS:I I1_1_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_1_1_0_0_R0_MINUS:I I1_1_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_0_0_0_R0_MINUS:I I1_1_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_1_2_1_0_0_R0_MINUS:I I1_1_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_0_0_0_R0_MINUS:I I1_1_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_0_1_0_0_R0_MINUS:I I1_1_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_0_0_0_R0_MINUS:I I1_1_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_1_1_0_0_R0_MINUS:I I1_1_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_0_0_0_R0_MINUS:I I1_1_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_1_2_2_1_0_0_R0_MINUS:I I1_1_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_0_0_0_R0_MINUS:I I1_2_0_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_0_1_0_0_R0_MINUS:I I1_2_0_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_0_0_0_R0_MINUS:I I1_2_0_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_1_1_0_0_R0_MINUS:I I1_2_0_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_0_0_0_R0_MINUS:I I1_2_0_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_0_2_1_0_0_R0_MINUS:I I1_2_0_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_0_0_0_R0_MINUS:I I1_2_1_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_0_1_0_0_R0_MINUS:I I1_2_1_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_0_0_0_R0_MINUS:I I1_2_1_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_1_1_0_0_R0_MINUS:I I1_2_1_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_0_0_0_R0_MINUS:I I1_2_1_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_1_2_1_0_0_R0_MINUS:I I1_2_1_2_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_0_0_0_R0_MINUS:I I1_2_2_0_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_0_1_0_0_R0_MINUS:I I1_2_2_0_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_0_0_0_R0_MINUS:I I1_2_2_1_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_1_1_0_0_R0_MINUS:I I1_2_2_1_1_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_0_0_0_R0_MINUS:I I1_2_2_2_0_0_0_R0_PLUS:I 
*.PININFO I1_2_2_2_1_0_0_R0_MINUS:I I1_2_2_2_1_0_0_R0_PLUS:I 
*.PININFO I1_default_MINUS:I I1_default_PLUS:I gnd!:I
RI1_2_2_2_1_0_0_R0 I1_2_2_2_1_0_0_R0_PLUS I1_2_2_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=50u w=50u r=311.93 par=8.0 s=1
RI1_2_2_2_0_0_0_R0 I1_2_2_2_0_0_0_R0_PLUS I1_2_2_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=50u r=311.93 par=1.0 s=8
RI1_2_2_1_1_0_0_R0 I1_2_2_1_1_0_0_R0_PLUS I1_2_2_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=50u w=50u r=311.93 par=3.0 s=1
RI1_2_2_1_0_0_0_R0 I1_2_2_1_0_0_0_R0_PLUS I1_2_2_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=50u r=311.93 par=1.0 s=3
RI1_2_2_0_1_0_0_R0 I1_2_2_0_1_0_0_R0_PLUS I1_2_2_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=50u r=311.93 par=1.0 s=1
RI1_2_2_0_0_0_0_R0 I1_2_2_0_0_0_0_R0_PLUS I1_2_2_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=50u r=311.93 par=1.0 s=1
RI1_2_1_2_1_0_0_R0 I1_2_1_2_1_0_0_R0_PLUS I1_2_1_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=7.6u w=50u r=48.7706 par=8.0 s=1
RI1_2_1_2_0_0_0_R0 I1_2_1_2_0_0_0_R0_PLUS I1_2_1_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=50u r=48.7706 par=1.0 s=8
RI1_2_1_1_1_0_0_R0 I1_2_1_1_1_0_0_R0_PLUS I1_2_1_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=7.6u w=50u r=48.7706 par=3.0 s=1
RI1_2_1_1_0_0_0_R0 I1_2_1_1_0_0_0_R0_PLUS I1_2_1_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=50u r=48.7706 par=1.0 s=3
RI1_2_1_0_1_0_0_R0 I1_2_1_0_1_0_0_R0_PLUS I1_2_1_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=50u r=48.7706 par=1.0 s=1
RI1_2_1_0_0_0_0_R0 I1_2_1_0_0_0_0_R0_PLUS I1_2_1_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=50u r=48.7706 par=1.0 s=1
RI1_2_0_2_1_0_0_R0 I1_2_0_2_1_0_0_R0_PLUS I1_2_0_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=1.6u w=50u r=11.5312 par=8.0 s=1
RI1_2_0_2_0_0_0_R0 I1_2_0_2_0_0_0_R0_PLUS I1_2_0_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=50u r=11.5312 par=1.0 s=8
RI1_2_0_1_1_0_0_R0 I1_2_0_1_1_0_0_R0_PLUS I1_2_0_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=1.6u w=50u r=11.5312 par=3.0 s=1
RI1_2_0_1_0_0_0_R0 I1_2_0_1_0_0_0_R0_PLUS I1_2_0_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=50u r=11.5312 par=1.0 s=3
RI1_2_0_0_1_0_0_R0 I1_2_0_0_1_0_0_R0_PLUS I1_2_0_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=50u r=11.5312 par=1.0 s=1
RI1_2_0_0_0_0_0_R0 I1_2_0_0_0_0_0_R0_PLUS I1_2_0_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=50u r=11.5312 par=1.0 s=1
RI1_1_2_2_1_0_0_R0 I1_1_2_2_1_0_0_R0_PLUS I1_1_2_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=50u w=3.62u r=4.3678K par=8.0 s=1
RI1_1_2_2_0_0_0_R0 I1_1_2_2_0_0_0_R0_PLUS I1_1_2_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=3.62u r=4.3678K par=1.0 s=8
RI1_1_2_1_1_0_0_R0 I1_1_2_1_1_0_0_R0_PLUS I1_1_2_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=50u w=3.62u r=4.3678K par=3.0 s=1
RI1_1_2_1_0_0_0_R0 I1_1_2_1_0_0_0_R0_PLUS I1_1_2_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=3.62u r=4.3678K par=1.0 s=3
RI1_1_2_0_1_0_0_R0 I1_1_2_0_1_0_0_R0_PLUS I1_1_2_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=3.62u r=4.3678K par=1.0 s=1
RI1_1_2_0_0_0_0_R0 I1_1_2_0_0_0_0_R0_PLUS I1_1_2_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=3.62u r=4.3678K par=1.0 s=1
RI1_1_1_2_1_0_0_R0 I1_1_1_2_1_0_0_R0_PLUS I1_1_1_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=7.6u w=3.62u r=682.912 par=8.0 s=1
RI1_1_1_2_0_0_0_R0 I1_1_1_2_0_0_0_R0_PLUS I1_1_1_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=3.62u r=682.912 par=1.0 s=8
RI1_1_1_1_1_0_0_R0 I1_1_1_1_1_0_0_R0_PLUS I1_1_1_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=7.6u w=3.62u r=682.912 par=3.0 s=1
RI1_1_1_1_0_0_0_R0 I1_1_1_1_0_0_0_R0_PLUS I1_1_1_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=3.62u r=682.912 par=1.0 s=3
RI1_1_1_0_1_0_0_R0 I1_1_1_0_1_0_0_R0_PLUS I1_1_1_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=3.62u r=682.912 par=1.0 s=1
RI1_1_1_0_0_0_0_R0 I1_1_1_0_0_0_0_R0_PLUS I1_1_1_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=3.62u r=682.912 par=1.0 s=1
RI1_1_0_2_1_0_0_R0 I1_1_0_2_1_0_0_R0_PLUS I1_1_0_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=1.6u w=3.62u r=161.465 par=8.0 s=1
RI1_1_0_2_0_0_0_R0 I1_1_0_2_0_0_0_R0_PLUS I1_1_0_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=3.62u r=161.465 par=1.0 s=8
RI1_1_0_1_1_0_0_R0 I1_1_0_1_1_0_0_R0_PLUS I1_1_0_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=1.6u w=3.62u r=161.465 par=3.0 s=1
RI1_1_0_1_0_0_0_R0 I1_1_0_1_0_0_0_R0_PLUS I1_1_0_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=3.62u r=161.465 par=1.0 s=3
RI1_1_0_0_1_0_0_R0 I1_1_0_0_1_0_0_R0_PLUS I1_1_0_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=3.62u r=161.465 par=1.0 s=1
RI1_1_0_0_0_0_0_R0 I1_1_0_0_0_0_0_R0_PLUS I1_1_0_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=3.62u r=161.465 par=1.0 s=1
RI1_0_2_2_1_0_0_R0 I1_0_2_2_1_0_0_R0_PLUS I1_0_2_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=50u w=800n r=20.8567K par=8.0 s=1
RI1_0_2_2_0_0_0_R0 I1_0_2_2_0_0_0_R0_PLUS I1_0_2_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=800n r=20.8567K par=1.0 s=8
RI1_0_2_1_1_0_0_R0 I1_0_2_1_1_0_0_R0_PLUS I1_0_2_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=50u w=800n r=20.8567K par=3.0 s=1
RI1_0_2_1_0_0_0_R0 I1_0_2_1_0_0_0_R0_PLUS I1_0_2_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=800n r=20.8567K par=1.0 s=3
RI1_0_2_0_1_0_0_R0 I1_0_2_0_1_0_0_R0_PLUS I1_0_2_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=800n r=20.8567K par=1.0 s=1
RI1_0_2_0_0_0_0_R0 I1_0_2_0_0_0_0_R0_PLUS I1_0_2_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=50u w=800n r=20.8567K par=1.0 s=1
RI1_0_1_2_1_0_0_R0 I1_0_1_2_1_0_0_R0_PLUS I1_0_1_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=7.6u w=800n r=3.26097K par=8.0 s=1
RI1_0_1_2_0_0_0_R0 I1_0_1_2_0_0_0_R0_PLUS I1_0_1_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=800n r=3.26097K par=1.0 s=8
RI1_0_1_1_1_0_0_R0 I1_0_1_1_1_0_0_R0_PLUS I1_0_1_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=7.6u w=800n r=3.26097K par=3.0 s=1
RI1_0_1_1_0_0_0_R0 I1_0_1_1_0_0_0_R0_PLUS I1_0_1_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=800n r=3.26097K par=1.0 s=3
RI1_0_1_0_1_0_0_R0 I1_0_1_0_1_0_0_R0_PLUS I1_0_1_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=800n r=3.26097K par=1.0 s=1
RI1_0_1_0_0_0_0_R0 I1_0_1_0_0_0_0_R0_PLUS I1_0_1_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=7.6u w=800n r=3.26097K par=1.0 s=1
RI1_0_0_2_1_0_0_R0 I1_0_0_2_1_0_0_R0_PLUS I1_0_0_2_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=8.0 l=1.6u w=800n r=771.014 par=8.0 s=1
RI1_0_0_2_0_0_0_R0 I1_0_0_2_0_0_0_R0_PLUS I1_0_0_2_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=800n r=771.014 par=1.0 s=8
RI1_0_0_1_1_0_0_R0 I1_0_0_1_1_0_0_R0_PLUS I1_0_0_1_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=3.0 l=1.6u w=800n r=771.014 par=3.0 s=1
RI1_0_0_1_0_0_0_R0 I1_0_0_1_0_0_0_R0_PLUS I1_0_0_1_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=800n r=771.014 par=1.0 s=3
RI1_0_0_0_1_0_0_R0 I1_0_0_0_1_0_0_R0_PLUS I1_0_0_0_1_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=800n r=771.014 par=1.0 s=1
RI1_0_0_0_0_0_0_R0 I1_0_0_0_0_0_0_R0_PLUS I1_0_0_0_0_0_0_R0_MINUS gnd! 
+ npolyf_u m=1.0 l=1.6u w=800n r=771.014 par=1.0 s=1
RI1_default I1_default_PLUS I1_default_MINUS gnd! npolyf_u m=1.0 
+ l=1.6u w=800.0n r=771.014 par=1.0 s=1
.ENDS

