magic
tech gf180mcuB
magscale 1 10
timestamp 1698431365
<< pwell >>
rect 1077 693 1553 993
rect 1077 1 1553 301
<< mvndiff >>
rect 1077 956 1165 993
rect 1077 910 1090 956
rect 1136 910 1165 956
rect 1077 776 1165 910
rect 1077 730 1090 776
rect 1136 730 1165 776
rect 1077 693 1165 730
rect 1465 956 1553 993
rect 1465 910 1494 956
rect 1540 910 1553 956
rect 1465 776 1553 910
rect 1465 730 1494 776
rect 1540 730 1553 776
rect 1465 693 1553 730
rect 1077 264 1165 301
rect 1077 218 1090 264
rect 1136 218 1165 264
rect 1077 84 1165 218
rect 1077 38 1090 84
rect 1136 38 1165 84
rect 1077 1 1165 38
rect 1465 264 1553 301
rect 1465 218 1494 264
rect 1540 218 1553 264
rect 1465 84 1553 218
rect 1465 38 1494 84
rect 1540 38 1553 84
rect 1465 1 1553 38
<< mvndiffc >>
rect 1090 910 1136 956
rect 1090 730 1136 776
rect 1494 910 1540 956
rect 1494 730 1540 776
rect 1090 218 1136 264
rect 1090 38 1136 84
rect 1494 218 1540 264
rect 1494 38 1540 84
<< mvnmoscap >>
rect 1165 693 1465 993
rect 1165 1 1465 301
<< polysilicon >>
rect 1165 1072 1465 1085
rect 1165 1026 1218 1072
rect 1264 1026 1366 1072
rect 1412 1026 1465 1072
rect 1165 993 1465 1026
rect 1165 660 1465 693
rect 1165 614 1218 660
rect 1264 614 1366 660
rect 1412 614 1465 660
rect 1165 601 1465 614
rect 1165 380 1465 393
rect 1165 334 1218 380
rect 1264 334 1366 380
rect 1412 334 1465 380
rect 1165 301 1465 334
rect 1165 -32 1465 1
rect 1165 -78 1218 -32
rect 1264 -78 1366 -32
rect 1412 -78 1465 -32
rect 1165 -91 1465 -78
<< polycontact >>
rect 1218 1026 1264 1072
rect 1366 1026 1412 1072
rect 1218 614 1264 660
rect 1366 614 1412 660
rect 1218 334 1264 380
rect 1366 334 1412 380
rect 1218 -78 1264 -32
rect 1366 -78 1412 -32
<< metal1 >>
rect 880 1143 1727 1343
rect 880 956 1147 1143
rect 880 910 1090 956
rect 1136 910 1147 956
rect 880 776 1147 910
rect 880 730 1090 776
rect 1136 730 1147 776
rect 880 264 1147 730
rect 1207 1072 1423 1083
rect 1207 1026 1218 1072
rect 1264 1071 1366 1072
rect 1264 1026 1290 1071
rect 1207 1019 1290 1026
rect 1342 1026 1366 1071
rect 1412 1026 1423 1072
rect 1342 1019 1423 1026
rect 1207 667 1423 1019
rect 1207 660 1290 667
rect 1207 614 1218 660
rect 1264 615 1290 660
rect 1342 660 1423 667
rect 1342 615 1366 660
rect 1264 614 1366 615
rect 1412 614 1423 660
rect 1207 603 1423 614
rect 1483 956 1727 1143
rect 1483 910 1494 956
rect 1540 910 1727 956
rect 1483 776 1727 910
rect 1483 730 1494 776
rect 1540 730 1727 776
rect 880 218 1090 264
rect 1136 218 1147 264
rect 880 84 1147 218
rect 880 38 1090 84
rect 1136 38 1147 84
rect 880 -149 1147 38
rect 1207 380 1423 391
rect 1207 334 1218 380
rect 1264 379 1366 380
rect 1264 334 1290 379
rect 1207 327 1290 334
rect 1342 334 1366 379
rect 1412 334 1423 380
rect 1342 327 1423 334
rect 1207 -25 1423 327
rect 1207 -32 1290 -25
rect 1207 -78 1218 -32
rect 1264 -77 1290 -32
rect 1342 -32 1423 -25
rect 1342 -77 1366 -32
rect 1264 -78 1366 -77
rect 1412 -78 1423 -32
rect 1207 -89 1423 -78
rect 1483 264 1727 730
rect 1483 218 1494 264
rect 1540 218 1727 264
rect 1483 84 1727 218
rect 1483 38 1494 84
rect 1540 38 1727 84
rect 1483 -149 1727 38
rect 880 -349 1727 -149
<< via1 >>
rect 1290 1019 1342 1071
rect 1290 615 1342 667
rect 1290 327 1342 379
rect 1290 -77 1342 -25
<< metal2 >>
rect 1278 1071 1354 1343
rect 1278 1019 1290 1071
rect 1342 1019 1354 1071
rect 1278 667 1354 1019
rect 1278 615 1290 667
rect 1342 615 1354 667
rect 1278 379 1354 615
rect 1278 327 1290 379
rect 1342 327 1354 379
rect 1278 -25 1354 327
rect 1278 -77 1290 -25
rect 1342 -77 1354 -25
rect 1278 -349 1354 -77
use M2_M1_CDNS_40661954729320  M2_M1_CDNS_40661954729320_0
timestamp 1698431365
transform 1 0 1316 0 -1 353
box 0 0 1 1
use M2_M1_CDNS_40661954729320  M2_M1_CDNS_40661954729320_1
timestamp 1698431365
transform 1 0 1316 0 1 641
box 0 0 1 1
use M2_M1_CDNS_40661954729320  M2_M1_CDNS_40661954729320_2
timestamp 1698431365
transform 1 0 1316 0 1 -51
box 0 0 1 1
use M2_M1_CDNS_40661954729320  M2_M1_CDNS_40661954729320_3
timestamp 1698431365
transform 1 0 1316 0 1 1045
box 0 0 1 1
<< properties >>
string GDS_END 4686750
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4683532
<< end >>
