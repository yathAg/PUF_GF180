magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< isosubstrate >>
rect 2267 55971 14818 57307
rect 4664 55935 7604 55971
rect 9908 55935 12848 55971
rect 10564 42616 14743 43682
rect 11970 40982 14743 42616
<< nwell >>
rect 354 55007 1644 56793
rect 873 54844 1644 55007
rect 873 53312 2754 54844
rect 11242 40947 11874 42043
<< pwell >>
rect 2760 56401 3760 56877
rect 4260 56401 5260 56877
rect 5760 56401 6760 56877
rect 7260 56401 8260 56877
rect 8760 56401 9760 56877
rect 10260 56401 11260 56877
rect 11760 56401 12760 56877
rect 13260 56401 14260 56877
rect 12482 42428 13082 43204
rect 13622 42428 14222 43204
rect 12482 41460 13082 42236
rect 13622 41460 14222 42236
<< mvndiff >>
rect 2760 56864 3760 56877
rect 2760 56818 2797 56864
rect 3723 56818 3760 56864
rect 2760 56789 3760 56818
rect 4260 56864 5260 56877
rect 4260 56818 4297 56864
rect 5223 56818 5260 56864
rect 4260 56789 5260 56818
rect 5760 56864 6760 56877
rect 5760 56818 5797 56864
rect 6723 56818 6760 56864
rect 5760 56789 6760 56818
rect 7260 56864 8260 56877
rect 7260 56818 7297 56864
rect 8223 56818 8260 56864
rect 7260 56789 8260 56818
rect 8760 56864 9760 56877
rect 8760 56818 8797 56864
rect 9723 56818 9760 56864
rect 8760 56789 9760 56818
rect 10260 56864 11260 56877
rect 10260 56818 10297 56864
rect 11223 56818 11260 56864
rect 10260 56789 11260 56818
rect 11760 56864 12760 56877
rect 11760 56818 11797 56864
rect 12723 56818 12760 56864
rect 11760 56789 12760 56818
rect 13260 56864 14260 56877
rect 13260 56818 13297 56864
rect 14223 56818 14260 56864
rect 13260 56789 14260 56818
rect 2760 56460 3760 56489
rect 2760 56414 2797 56460
rect 3723 56414 3760 56460
rect 2760 56401 3760 56414
rect 4260 56460 5260 56489
rect 4260 56414 4297 56460
rect 5223 56414 5260 56460
rect 4260 56401 5260 56414
rect 5760 56460 6760 56489
rect 5760 56414 5797 56460
rect 6723 56414 6760 56460
rect 5760 56401 6760 56414
rect 7260 56460 8260 56489
rect 7260 56414 7297 56460
rect 8223 56414 8260 56460
rect 7260 56401 8260 56414
rect 8760 56460 9760 56489
rect 8760 56414 8797 56460
rect 9723 56414 9760 56460
rect 8760 56401 9760 56414
rect 10260 56460 11260 56489
rect 10260 56414 10297 56460
rect 11223 56414 11260 56460
rect 10260 56401 11260 56414
rect 11760 56460 12760 56489
rect 11760 56414 11797 56460
rect 12723 56414 12760 56460
rect 11760 56401 12760 56414
rect 13260 56460 14260 56489
rect 13260 56414 13297 56460
rect 14223 56414 14260 56460
rect 13260 56401 14260 56414
rect 12482 43191 13082 43204
rect 12482 43145 12519 43191
rect 13045 43145 13082 43191
rect 12482 43116 13082 43145
rect 13622 43191 14222 43204
rect 13622 43145 13659 43191
rect 14185 43145 14222 43191
rect 13622 43116 14222 43145
rect 12482 42487 13082 42516
rect 12482 42441 12519 42487
rect 13045 42441 13082 42487
rect 12482 42428 13082 42441
rect 13622 42487 14222 42516
rect 13622 42441 13659 42487
rect 14185 42441 14222 42487
rect 13622 42428 14222 42441
rect 12482 42223 13082 42236
rect 12482 42177 12519 42223
rect 13045 42177 13082 42223
rect 12482 42148 13082 42177
rect 13622 42223 14222 42236
rect 13622 42177 13659 42223
rect 14185 42177 14222 42223
rect 13622 42148 14222 42177
rect 12482 41519 13082 41548
rect 12482 41473 12519 41519
rect 13045 41473 13082 41519
rect 12482 41460 13082 41473
rect 13622 41519 14222 41548
rect 13622 41473 13659 41519
rect 14185 41473 14222 41519
rect 13622 41460 14222 41473
<< mvndiffc >>
rect 2797 56818 3723 56864
rect 4297 56818 5223 56864
rect 5797 56818 6723 56864
rect 7297 56818 8223 56864
rect 8797 56818 9723 56864
rect 10297 56818 11223 56864
rect 11797 56818 12723 56864
rect 13297 56818 14223 56864
rect 2797 56414 3723 56460
rect 4297 56414 5223 56460
rect 5797 56414 6723 56460
rect 7297 56414 8223 56460
rect 8797 56414 9723 56460
rect 10297 56414 11223 56460
rect 11797 56414 12723 56460
rect 13297 56414 14223 56460
rect 12519 43145 13045 43191
rect 13659 43145 14185 43191
rect 12519 42441 13045 42487
rect 13659 42441 14185 42487
rect 12519 42177 13045 42223
rect 13659 42177 14185 42223
rect 12519 41473 13045 41519
rect 13659 41473 14185 41519
<< psubdiff >>
rect 2331 57202 14735 57224
rect 2331 57156 2353 57202
rect 14713 57156 14735 57202
rect 2331 57134 14735 57156
rect 2331 57038 2421 57134
rect 2331 56240 2353 57038
rect 2399 56240 2421 57038
rect 14645 57038 14735 57134
rect 2331 56144 2421 56240
rect 14645 56240 14667 57038
rect 14713 56240 14735 57038
rect 14645 56144 14735 56240
rect 2331 56122 14735 56144
rect 2331 56076 2353 56122
rect 14713 56076 14735 56122
rect 2331 56054 14735 56076
rect 10742 43628 11858 43650
rect 10742 43582 10764 43628
rect 10810 43582 10878 43628
rect 10924 43582 10992 43628
rect 11038 43582 11106 43628
rect 11152 43582 11220 43628
rect 11266 43582 11334 43628
rect 11380 43582 11448 43628
rect 11494 43582 11562 43628
rect 11608 43582 11676 43628
rect 11722 43582 11790 43628
rect 11836 43582 11858 43628
rect 10742 43514 11858 43582
rect 10742 43468 10764 43514
rect 10810 43468 10878 43514
rect 10924 43468 10992 43514
rect 11038 43468 11106 43514
rect 11152 43468 11220 43514
rect 11266 43468 11334 43514
rect 11380 43468 11448 43514
rect 11494 43468 11562 43514
rect 11608 43468 11676 43514
rect 11722 43468 11790 43514
rect 11836 43468 11858 43514
rect 10742 43400 11858 43468
rect 10742 43354 10764 43400
rect 10810 43354 10878 43400
rect 10924 43354 10992 43400
rect 11038 43354 11106 43400
rect 11152 43354 11220 43400
rect 11266 43354 11334 43400
rect 11380 43354 11448 43400
rect 11494 43354 11562 43400
rect 11608 43354 11676 43400
rect 11722 43354 11790 43400
rect 11836 43354 11858 43400
rect 10742 43286 11858 43354
rect 10742 43240 10764 43286
rect 10810 43240 10878 43286
rect 10924 43240 10992 43286
rect 11038 43240 11106 43286
rect 11152 43240 11220 43286
rect 11266 43240 11334 43286
rect 11380 43240 11448 43286
rect 11494 43240 11562 43286
rect 11608 43240 11676 43286
rect 11722 43240 11790 43286
rect 11836 43240 11858 43286
rect 10742 43172 11858 43240
rect 10742 43126 10764 43172
rect 10810 43126 10878 43172
rect 10924 43126 10992 43172
rect 11038 43126 11106 43172
rect 11152 43126 11220 43172
rect 11266 43126 11334 43172
rect 11380 43126 11448 43172
rect 11494 43126 11562 43172
rect 11608 43126 11676 43172
rect 11722 43126 11790 43172
rect 11836 43126 11858 43172
rect 10742 43058 11858 43126
rect 10742 43012 10764 43058
rect 10810 43012 10878 43058
rect 10924 43012 10992 43058
rect 11038 43012 11106 43058
rect 11152 43012 11220 43058
rect 11266 43012 11334 43058
rect 11380 43012 11448 43058
rect 11494 43012 11562 43058
rect 11608 43012 11676 43058
rect 11722 43012 11790 43058
rect 11836 43012 11858 43058
rect 10742 42944 11858 43012
rect 10742 42898 10764 42944
rect 10810 42898 10878 42944
rect 10924 42898 10992 42944
rect 11038 42898 11106 42944
rect 11152 42898 11220 42944
rect 11266 42898 11334 42944
rect 11380 42898 11448 42944
rect 11494 42898 11562 42944
rect 11608 42898 11676 42944
rect 11722 42898 11790 42944
rect 11836 42898 11858 42944
rect 10742 42830 11858 42898
rect 10742 42784 10764 42830
rect 10810 42784 10878 42830
rect 10924 42784 10992 42830
rect 11038 42784 11106 42830
rect 11152 42784 11220 42830
rect 11266 42784 11334 42830
rect 11380 42784 11448 42830
rect 11494 42784 11562 42830
rect 11608 42784 11676 42830
rect 11722 42784 11790 42830
rect 11836 42784 11858 42830
rect 10742 42716 11858 42784
rect 10742 42670 10764 42716
rect 10810 42670 10878 42716
rect 10924 42670 10992 42716
rect 11038 42670 11106 42716
rect 11152 42670 11220 42716
rect 11266 42670 11334 42716
rect 11380 42670 11448 42716
rect 11494 42670 11562 42716
rect 11608 42670 11676 42716
rect 11722 42670 11790 42716
rect 11836 42670 11858 42716
rect 10742 42648 11858 42670
rect 12053 43577 14660 43599
rect 12053 41087 12075 43577
rect 12121 43531 12182 43577
rect 14484 43531 14592 43577
rect 12121 43509 14592 43531
rect 12121 41155 12143 43509
rect 14570 41155 14592 43509
rect 12121 41133 14592 41155
rect 12121 41087 12182 41133
rect 14484 41087 14592 41133
rect 14638 41087 14660 43577
rect 12053 41065 14660 41087
rect 189 10991 279 11013
rect 189 1357 211 10991
rect 257 1357 279 10991
rect 189 1335 279 1357
rect 14723 10991 14813 11013
rect 14723 1357 14745 10991
rect 14791 1357 14813 10991
rect 14723 1335 14813 1357
rect 265 1206 14739 1228
rect 265 1160 287 1206
rect 333 1160 411 1206
rect 457 1160 535 1206
rect 581 1160 659 1206
rect 705 1160 783 1206
rect 829 1160 907 1206
rect 953 1160 1031 1206
rect 1077 1160 1155 1206
rect 1201 1160 1279 1206
rect 1325 1160 1403 1206
rect 1449 1160 1527 1206
rect 1573 1160 1651 1206
rect 1697 1160 1775 1206
rect 1821 1160 1899 1206
rect 1945 1160 2023 1206
rect 2069 1160 2147 1206
rect 2193 1160 2271 1206
rect 2317 1160 2395 1206
rect 2441 1160 2519 1206
rect 2565 1160 2643 1206
rect 2689 1160 2767 1206
rect 2813 1160 2891 1206
rect 2937 1160 3015 1206
rect 3061 1160 3139 1206
rect 3185 1160 3263 1206
rect 3309 1160 3387 1206
rect 3433 1160 3511 1206
rect 3557 1160 3635 1206
rect 3681 1160 3759 1206
rect 3805 1160 3883 1206
rect 3929 1160 4007 1206
rect 4053 1160 4131 1206
rect 4177 1160 4255 1206
rect 4301 1160 4379 1206
rect 4425 1160 4503 1206
rect 4549 1160 4627 1206
rect 4673 1160 4751 1206
rect 4797 1160 4875 1206
rect 4921 1160 4999 1206
rect 5045 1160 5123 1206
rect 5169 1160 5247 1206
rect 5293 1160 5371 1206
rect 5417 1160 5495 1206
rect 5541 1160 5619 1206
rect 5665 1160 5743 1206
rect 5789 1160 5867 1206
rect 5913 1160 5991 1206
rect 6037 1160 6115 1206
rect 6161 1160 6239 1206
rect 6285 1160 6363 1206
rect 6409 1160 6487 1206
rect 6533 1160 6611 1206
rect 6657 1160 6735 1206
rect 6781 1160 6859 1206
rect 6905 1160 6983 1206
rect 7029 1160 7107 1206
rect 7153 1160 7231 1206
rect 7277 1160 7355 1206
rect 7401 1160 7479 1206
rect 7525 1160 7603 1206
rect 7649 1160 7727 1206
rect 7773 1160 7851 1206
rect 7897 1160 7975 1206
rect 8021 1160 8099 1206
rect 8145 1160 8223 1206
rect 8269 1160 8347 1206
rect 8393 1160 8471 1206
rect 8517 1160 8595 1206
rect 8641 1160 8719 1206
rect 8765 1160 8843 1206
rect 8889 1160 8967 1206
rect 9013 1160 9091 1206
rect 9137 1160 9215 1206
rect 9261 1160 9339 1206
rect 9385 1160 9463 1206
rect 9509 1160 9587 1206
rect 9633 1160 9711 1206
rect 9757 1160 9835 1206
rect 9881 1160 9959 1206
rect 10005 1160 10083 1206
rect 10129 1160 10207 1206
rect 10253 1160 10331 1206
rect 10377 1160 10455 1206
rect 10501 1160 10579 1206
rect 10625 1160 10703 1206
rect 10749 1160 10827 1206
rect 10873 1160 10951 1206
rect 10997 1160 11075 1206
rect 11121 1160 11199 1206
rect 11245 1160 11323 1206
rect 11369 1160 11447 1206
rect 11493 1160 11571 1206
rect 11617 1160 11695 1206
rect 11741 1160 11819 1206
rect 11865 1160 11943 1206
rect 11989 1160 12067 1206
rect 12113 1160 12191 1206
rect 12237 1160 12315 1206
rect 12361 1160 12439 1206
rect 12485 1160 12563 1206
rect 12609 1160 12687 1206
rect 12733 1160 12811 1206
rect 12857 1160 12935 1206
rect 12981 1160 13059 1206
rect 13105 1160 13183 1206
rect 13229 1160 13307 1206
rect 13353 1160 13431 1206
rect 13477 1160 13555 1206
rect 13601 1160 13679 1206
rect 13725 1160 13803 1206
rect 13849 1160 13927 1206
rect 13973 1160 14051 1206
rect 14097 1160 14175 1206
rect 14221 1160 14299 1206
rect 14345 1160 14423 1206
rect 14469 1160 14547 1206
rect 14593 1160 14671 1206
rect 14717 1160 14739 1206
rect 265 1082 14739 1160
rect 265 1036 287 1082
rect 333 1036 411 1082
rect 457 1036 535 1082
rect 581 1036 659 1082
rect 705 1036 783 1082
rect 829 1036 907 1082
rect 953 1036 1031 1082
rect 1077 1036 1155 1082
rect 1201 1036 1279 1082
rect 1325 1036 1403 1082
rect 1449 1036 1527 1082
rect 1573 1036 1651 1082
rect 1697 1036 1775 1082
rect 1821 1036 1899 1082
rect 1945 1036 2023 1082
rect 2069 1036 2147 1082
rect 2193 1036 2271 1082
rect 2317 1036 2395 1082
rect 2441 1036 2519 1082
rect 2565 1036 2643 1082
rect 2689 1036 2767 1082
rect 2813 1036 2891 1082
rect 2937 1036 3015 1082
rect 3061 1036 3139 1082
rect 3185 1036 3263 1082
rect 3309 1036 3387 1082
rect 3433 1036 3511 1082
rect 3557 1036 3635 1082
rect 3681 1036 3759 1082
rect 3805 1036 3883 1082
rect 3929 1036 4007 1082
rect 4053 1036 4131 1082
rect 4177 1036 4255 1082
rect 4301 1036 4379 1082
rect 4425 1036 4503 1082
rect 4549 1036 4627 1082
rect 4673 1036 4751 1082
rect 4797 1036 4875 1082
rect 4921 1036 4999 1082
rect 5045 1036 5123 1082
rect 5169 1036 5247 1082
rect 5293 1036 5371 1082
rect 5417 1036 5495 1082
rect 5541 1036 5619 1082
rect 5665 1036 5743 1082
rect 5789 1036 5867 1082
rect 5913 1036 5991 1082
rect 6037 1036 6115 1082
rect 6161 1036 6239 1082
rect 6285 1036 6363 1082
rect 6409 1036 6487 1082
rect 6533 1036 6611 1082
rect 6657 1036 6735 1082
rect 6781 1036 6859 1082
rect 6905 1036 6983 1082
rect 7029 1036 7107 1082
rect 7153 1036 7231 1082
rect 7277 1036 7355 1082
rect 7401 1036 7479 1082
rect 7525 1036 7603 1082
rect 7649 1036 7727 1082
rect 7773 1036 7851 1082
rect 7897 1036 7975 1082
rect 8021 1036 8099 1082
rect 8145 1036 8223 1082
rect 8269 1036 8347 1082
rect 8393 1036 8471 1082
rect 8517 1036 8595 1082
rect 8641 1036 8719 1082
rect 8765 1036 8843 1082
rect 8889 1036 8967 1082
rect 9013 1036 9091 1082
rect 9137 1036 9215 1082
rect 9261 1036 9339 1082
rect 9385 1036 9463 1082
rect 9509 1036 9587 1082
rect 9633 1036 9711 1082
rect 9757 1036 9835 1082
rect 9881 1036 9959 1082
rect 10005 1036 10083 1082
rect 10129 1036 10207 1082
rect 10253 1036 10331 1082
rect 10377 1036 10455 1082
rect 10501 1036 10579 1082
rect 10625 1036 10703 1082
rect 10749 1036 10827 1082
rect 10873 1036 10951 1082
rect 10997 1036 11075 1082
rect 11121 1036 11199 1082
rect 11245 1036 11323 1082
rect 11369 1036 11447 1082
rect 11493 1036 11571 1082
rect 11617 1036 11695 1082
rect 11741 1036 11819 1082
rect 11865 1036 11943 1082
rect 11989 1036 12067 1082
rect 12113 1036 12191 1082
rect 12237 1036 12315 1082
rect 12361 1036 12439 1082
rect 12485 1036 12563 1082
rect 12609 1036 12687 1082
rect 12733 1036 12811 1082
rect 12857 1036 12935 1082
rect 12981 1036 13059 1082
rect 13105 1036 13183 1082
rect 13229 1036 13307 1082
rect 13353 1036 13431 1082
rect 13477 1036 13555 1082
rect 13601 1036 13679 1082
rect 13725 1036 13803 1082
rect 13849 1036 13927 1082
rect 13973 1036 14051 1082
rect 14097 1036 14175 1082
rect 14221 1036 14299 1082
rect 14345 1036 14423 1082
rect 14469 1036 14547 1082
rect 14593 1036 14671 1082
rect 14717 1036 14739 1082
rect 265 1014 14739 1036
<< nsubdiff >>
rect 437 56688 1561 56710
rect 437 56642 459 56688
rect 975 56642 1305 56688
rect 1539 56642 1561 56688
rect 437 56620 1561 56642
rect 437 56534 527 56620
rect 437 55266 459 56534
rect 505 55266 527 56534
rect 1471 56534 1561 56620
rect 1471 56300 1493 56534
rect 1539 56300 1561 56534
rect 1471 56064 1561 56300
rect 1471 55548 1493 56064
rect 1539 55548 1561 56064
rect 437 55180 527 55266
rect 1471 55312 1561 55548
rect 1471 55266 1493 55312
rect 1539 55266 1561 55312
rect 1471 55180 1561 55266
rect 437 55158 1561 55180
rect 437 55112 459 55158
rect 1539 55112 1561 55158
rect 437 55090 1561 55112
<< mvnsubdiff >>
rect 11290 41982 11826 41995
rect 11290 41936 11303 41982
rect 11349 41936 11419 41982
rect 11465 41936 11535 41982
rect 11581 41936 11651 41982
rect 11697 41936 11767 41982
rect 11813 41936 11826 41982
rect 11290 41923 11826 41936
rect 11290 41866 11362 41923
rect 11290 41820 11303 41866
rect 11349 41820 11362 41866
rect 11754 41866 11826 41923
rect 11290 41750 11362 41820
rect 11290 41704 11303 41750
rect 11349 41704 11362 41750
rect 11290 41634 11362 41704
rect 11290 41588 11303 41634
rect 11349 41588 11362 41634
rect 11754 41820 11767 41866
rect 11813 41820 11826 41866
rect 11754 41750 11826 41820
rect 11754 41704 11767 41750
rect 11813 41704 11826 41750
rect 11754 41634 11826 41704
rect 11290 41531 11362 41588
rect 11754 41588 11767 41634
rect 11813 41588 11826 41634
rect 11754 41531 11826 41588
rect 11290 41518 11826 41531
rect 11290 41472 11303 41518
rect 11349 41472 11419 41518
rect 11465 41472 11535 41518
rect 11581 41472 11651 41518
rect 11697 41472 11767 41518
rect 11813 41472 11826 41518
rect 11290 41459 11826 41472
rect 11290 41402 11362 41459
rect 11290 41356 11303 41402
rect 11349 41356 11362 41402
rect 11754 41402 11826 41459
rect 11290 41286 11362 41356
rect 11290 41240 11303 41286
rect 11349 41240 11362 41286
rect 11290 41170 11362 41240
rect 11290 41124 11303 41170
rect 11349 41124 11362 41170
rect 11754 41356 11767 41402
rect 11813 41356 11826 41402
rect 11754 41286 11826 41356
rect 11754 41240 11767 41286
rect 11813 41240 11826 41286
rect 11754 41170 11826 41240
rect 11290 41067 11362 41124
rect 11754 41124 11767 41170
rect 11813 41124 11826 41170
rect 11754 41067 11826 41124
rect 11290 41054 11826 41067
rect 11290 41008 11303 41054
rect 11349 41008 11419 41054
rect 11465 41008 11535 41054
rect 11581 41008 11651 41054
rect 11697 41008 11767 41054
rect 11813 41008 11826 41054
rect 11290 40995 11826 41008
<< psubdiffcont >>
rect 2353 57156 14713 57202
rect 2353 56240 2399 57038
rect 14667 56240 14713 57038
rect 2353 56076 14713 56122
rect 10764 43582 10810 43628
rect 10878 43582 10924 43628
rect 10992 43582 11038 43628
rect 11106 43582 11152 43628
rect 11220 43582 11266 43628
rect 11334 43582 11380 43628
rect 11448 43582 11494 43628
rect 11562 43582 11608 43628
rect 11676 43582 11722 43628
rect 11790 43582 11836 43628
rect 10764 43468 10810 43514
rect 10878 43468 10924 43514
rect 10992 43468 11038 43514
rect 11106 43468 11152 43514
rect 11220 43468 11266 43514
rect 11334 43468 11380 43514
rect 11448 43468 11494 43514
rect 11562 43468 11608 43514
rect 11676 43468 11722 43514
rect 11790 43468 11836 43514
rect 10764 43354 10810 43400
rect 10878 43354 10924 43400
rect 10992 43354 11038 43400
rect 11106 43354 11152 43400
rect 11220 43354 11266 43400
rect 11334 43354 11380 43400
rect 11448 43354 11494 43400
rect 11562 43354 11608 43400
rect 11676 43354 11722 43400
rect 11790 43354 11836 43400
rect 10764 43240 10810 43286
rect 10878 43240 10924 43286
rect 10992 43240 11038 43286
rect 11106 43240 11152 43286
rect 11220 43240 11266 43286
rect 11334 43240 11380 43286
rect 11448 43240 11494 43286
rect 11562 43240 11608 43286
rect 11676 43240 11722 43286
rect 11790 43240 11836 43286
rect 10764 43126 10810 43172
rect 10878 43126 10924 43172
rect 10992 43126 11038 43172
rect 11106 43126 11152 43172
rect 11220 43126 11266 43172
rect 11334 43126 11380 43172
rect 11448 43126 11494 43172
rect 11562 43126 11608 43172
rect 11676 43126 11722 43172
rect 11790 43126 11836 43172
rect 10764 43012 10810 43058
rect 10878 43012 10924 43058
rect 10992 43012 11038 43058
rect 11106 43012 11152 43058
rect 11220 43012 11266 43058
rect 11334 43012 11380 43058
rect 11448 43012 11494 43058
rect 11562 43012 11608 43058
rect 11676 43012 11722 43058
rect 11790 43012 11836 43058
rect 10764 42898 10810 42944
rect 10878 42898 10924 42944
rect 10992 42898 11038 42944
rect 11106 42898 11152 42944
rect 11220 42898 11266 42944
rect 11334 42898 11380 42944
rect 11448 42898 11494 42944
rect 11562 42898 11608 42944
rect 11676 42898 11722 42944
rect 11790 42898 11836 42944
rect 10764 42784 10810 42830
rect 10878 42784 10924 42830
rect 10992 42784 11038 42830
rect 11106 42784 11152 42830
rect 11220 42784 11266 42830
rect 11334 42784 11380 42830
rect 11448 42784 11494 42830
rect 11562 42784 11608 42830
rect 11676 42784 11722 42830
rect 11790 42784 11836 42830
rect 10764 42670 10810 42716
rect 10878 42670 10924 42716
rect 10992 42670 11038 42716
rect 11106 42670 11152 42716
rect 11220 42670 11266 42716
rect 11334 42670 11380 42716
rect 11448 42670 11494 42716
rect 11562 42670 11608 42716
rect 11676 42670 11722 42716
rect 11790 42670 11836 42716
rect 12075 41087 12121 43577
rect 12182 43531 14484 43577
rect 12182 41087 14484 41133
rect 14592 41087 14638 43577
rect 211 1357 257 10991
rect 14745 1357 14791 10991
rect 287 1160 333 1206
rect 411 1160 457 1206
rect 535 1160 581 1206
rect 659 1160 705 1206
rect 783 1160 829 1206
rect 907 1160 953 1206
rect 1031 1160 1077 1206
rect 1155 1160 1201 1206
rect 1279 1160 1325 1206
rect 1403 1160 1449 1206
rect 1527 1160 1573 1206
rect 1651 1160 1697 1206
rect 1775 1160 1821 1206
rect 1899 1160 1945 1206
rect 2023 1160 2069 1206
rect 2147 1160 2193 1206
rect 2271 1160 2317 1206
rect 2395 1160 2441 1206
rect 2519 1160 2565 1206
rect 2643 1160 2689 1206
rect 2767 1160 2813 1206
rect 2891 1160 2937 1206
rect 3015 1160 3061 1206
rect 3139 1160 3185 1206
rect 3263 1160 3309 1206
rect 3387 1160 3433 1206
rect 3511 1160 3557 1206
rect 3635 1160 3681 1206
rect 3759 1160 3805 1206
rect 3883 1160 3929 1206
rect 4007 1160 4053 1206
rect 4131 1160 4177 1206
rect 4255 1160 4301 1206
rect 4379 1160 4425 1206
rect 4503 1160 4549 1206
rect 4627 1160 4673 1206
rect 4751 1160 4797 1206
rect 4875 1160 4921 1206
rect 4999 1160 5045 1206
rect 5123 1160 5169 1206
rect 5247 1160 5293 1206
rect 5371 1160 5417 1206
rect 5495 1160 5541 1206
rect 5619 1160 5665 1206
rect 5743 1160 5789 1206
rect 5867 1160 5913 1206
rect 5991 1160 6037 1206
rect 6115 1160 6161 1206
rect 6239 1160 6285 1206
rect 6363 1160 6409 1206
rect 6487 1160 6533 1206
rect 6611 1160 6657 1206
rect 6735 1160 6781 1206
rect 6859 1160 6905 1206
rect 6983 1160 7029 1206
rect 7107 1160 7153 1206
rect 7231 1160 7277 1206
rect 7355 1160 7401 1206
rect 7479 1160 7525 1206
rect 7603 1160 7649 1206
rect 7727 1160 7773 1206
rect 7851 1160 7897 1206
rect 7975 1160 8021 1206
rect 8099 1160 8145 1206
rect 8223 1160 8269 1206
rect 8347 1160 8393 1206
rect 8471 1160 8517 1206
rect 8595 1160 8641 1206
rect 8719 1160 8765 1206
rect 8843 1160 8889 1206
rect 8967 1160 9013 1206
rect 9091 1160 9137 1206
rect 9215 1160 9261 1206
rect 9339 1160 9385 1206
rect 9463 1160 9509 1206
rect 9587 1160 9633 1206
rect 9711 1160 9757 1206
rect 9835 1160 9881 1206
rect 9959 1160 10005 1206
rect 10083 1160 10129 1206
rect 10207 1160 10253 1206
rect 10331 1160 10377 1206
rect 10455 1160 10501 1206
rect 10579 1160 10625 1206
rect 10703 1160 10749 1206
rect 10827 1160 10873 1206
rect 10951 1160 10997 1206
rect 11075 1160 11121 1206
rect 11199 1160 11245 1206
rect 11323 1160 11369 1206
rect 11447 1160 11493 1206
rect 11571 1160 11617 1206
rect 11695 1160 11741 1206
rect 11819 1160 11865 1206
rect 11943 1160 11989 1206
rect 12067 1160 12113 1206
rect 12191 1160 12237 1206
rect 12315 1160 12361 1206
rect 12439 1160 12485 1206
rect 12563 1160 12609 1206
rect 12687 1160 12733 1206
rect 12811 1160 12857 1206
rect 12935 1160 12981 1206
rect 13059 1160 13105 1206
rect 13183 1160 13229 1206
rect 13307 1160 13353 1206
rect 13431 1160 13477 1206
rect 13555 1160 13601 1206
rect 13679 1160 13725 1206
rect 13803 1160 13849 1206
rect 13927 1160 13973 1206
rect 14051 1160 14097 1206
rect 14175 1160 14221 1206
rect 14299 1160 14345 1206
rect 14423 1160 14469 1206
rect 14547 1160 14593 1206
rect 14671 1160 14717 1206
rect 287 1036 333 1082
rect 411 1036 457 1082
rect 535 1036 581 1082
rect 659 1036 705 1082
rect 783 1036 829 1082
rect 907 1036 953 1082
rect 1031 1036 1077 1082
rect 1155 1036 1201 1082
rect 1279 1036 1325 1082
rect 1403 1036 1449 1082
rect 1527 1036 1573 1082
rect 1651 1036 1697 1082
rect 1775 1036 1821 1082
rect 1899 1036 1945 1082
rect 2023 1036 2069 1082
rect 2147 1036 2193 1082
rect 2271 1036 2317 1082
rect 2395 1036 2441 1082
rect 2519 1036 2565 1082
rect 2643 1036 2689 1082
rect 2767 1036 2813 1082
rect 2891 1036 2937 1082
rect 3015 1036 3061 1082
rect 3139 1036 3185 1082
rect 3263 1036 3309 1082
rect 3387 1036 3433 1082
rect 3511 1036 3557 1082
rect 3635 1036 3681 1082
rect 3759 1036 3805 1082
rect 3883 1036 3929 1082
rect 4007 1036 4053 1082
rect 4131 1036 4177 1082
rect 4255 1036 4301 1082
rect 4379 1036 4425 1082
rect 4503 1036 4549 1082
rect 4627 1036 4673 1082
rect 4751 1036 4797 1082
rect 4875 1036 4921 1082
rect 4999 1036 5045 1082
rect 5123 1036 5169 1082
rect 5247 1036 5293 1082
rect 5371 1036 5417 1082
rect 5495 1036 5541 1082
rect 5619 1036 5665 1082
rect 5743 1036 5789 1082
rect 5867 1036 5913 1082
rect 5991 1036 6037 1082
rect 6115 1036 6161 1082
rect 6239 1036 6285 1082
rect 6363 1036 6409 1082
rect 6487 1036 6533 1082
rect 6611 1036 6657 1082
rect 6735 1036 6781 1082
rect 6859 1036 6905 1082
rect 6983 1036 7029 1082
rect 7107 1036 7153 1082
rect 7231 1036 7277 1082
rect 7355 1036 7401 1082
rect 7479 1036 7525 1082
rect 7603 1036 7649 1082
rect 7727 1036 7773 1082
rect 7851 1036 7897 1082
rect 7975 1036 8021 1082
rect 8099 1036 8145 1082
rect 8223 1036 8269 1082
rect 8347 1036 8393 1082
rect 8471 1036 8517 1082
rect 8595 1036 8641 1082
rect 8719 1036 8765 1082
rect 8843 1036 8889 1082
rect 8967 1036 9013 1082
rect 9091 1036 9137 1082
rect 9215 1036 9261 1082
rect 9339 1036 9385 1082
rect 9463 1036 9509 1082
rect 9587 1036 9633 1082
rect 9711 1036 9757 1082
rect 9835 1036 9881 1082
rect 9959 1036 10005 1082
rect 10083 1036 10129 1082
rect 10207 1036 10253 1082
rect 10331 1036 10377 1082
rect 10455 1036 10501 1082
rect 10579 1036 10625 1082
rect 10703 1036 10749 1082
rect 10827 1036 10873 1082
rect 10951 1036 10997 1082
rect 11075 1036 11121 1082
rect 11199 1036 11245 1082
rect 11323 1036 11369 1082
rect 11447 1036 11493 1082
rect 11571 1036 11617 1082
rect 11695 1036 11741 1082
rect 11819 1036 11865 1082
rect 11943 1036 11989 1082
rect 12067 1036 12113 1082
rect 12191 1036 12237 1082
rect 12315 1036 12361 1082
rect 12439 1036 12485 1082
rect 12563 1036 12609 1082
rect 12687 1036 12733 1082
rect 12811 1036 12857 1082
rect 12935 1036 12981 1082
rect 13059 1036 13105 1082
rect 13183 1036 13229 1082
rect 13307 1036 13353 1082
rect 13431 1036 13477 1082
rect 13555 1036 13601 1082
rect 13679 1036 13725 1082
rect 13803 1036 13849 1082
rect 13927 1036 13973 1082
rect 14051 1036 14097 1082
rect 14175 1036 14221 1082
rect 14299 1036 14345 1082
rect 14423 1036 14469 1082
rect 14547 1036 14593 1082
rect 14671 1036 14717 1082
<< nsubdiffcont >>
rect 459 56642 975 56688
rect 1305 56642 1539 56688
rect 459 55266 505 56534
rect 1493 56300 1539 56534
rect 1493 55548 1539 56064
rect 1493 55266 1539 55312
rect 459 55112 1539 55158
<< mvnsubdiffcont >>
rect 11303 41936 11349 41982
rect 11419 41936 11465 41982
rect 11535 41936 11581 41982
rect 11651 41936 11697 41982
rect 11767 41936 11813 41982
rect 11303 41820 11349 41866
rect 11303 41704 11349 41750
rect 11303 41588 11349 41634
rect 11767 41820 11813 41866
rect 11767 41704 11813 41750
rect 11767 41588 11813 41634
rect 11303 41472 11349 41518
rect 11419 41472 11465 41518
rect 11535 41472 11581 41518
rect 11651 41472 11697 41518
rect 11767 41472 11813 41518
rect 11303 41356 11349 41402
rect 11303 41240 11349 41286
rect 11303 41124 11349 41170
rect 11767 41356 11813 41402
rect 11767 41240 11813 41286
rect 11767 41124 11813 41170
rect 11303 41008 11349 41054
rect 11419 41008 11465 41054
rect 11535 41008 11581 41054
rect 11651 41008 11697 41054
rect 11767 41008 11813 41054
<< mvnmoscap >>
rect 2760 56489 3760 56789
rect 4260 56489 5260 56789
rect 5760 56489 6760 56789
rect 7260 56489 8260 56789
rect 8760 56489 9760 56789
rect 10260 56489 11260 56789
rect 11760 56489 12760 56789
rect 13260 56489 14260 56789
rect 12482 42516 13082 43116
rect 13622 42516 14222 43116
rect 12482 41548 13082 42148
rect 13622 41548 14222 42148
<< polysilicon >>
rect 779 56372 939 56385
rect 779 56326 836 56372
rect 882 56326 939 56372
rect 779 56283 939 56326
rect 779 55460 939 55503
rect 779 55414 836 55460
rect 882 55414 939 55460
rect 779 55401 939 55414
rect 1059 56372 1219 56385
rect 1059 56326 1116 56372
rect 1162 56326 1219 56372
rect 1059 56283 1219 56326
rect 1059 55460 1219 55503
rect 1059 55414 1116 55460
rect 1162 55414 1219 55460
rect 1059 55401 1219 55414
rect 2668 56736 2760 56789
rect 2668 56690 2681 56736
rect 2727 56690 2760 56736
rect 2668 56588 2760 56690
rect 2668 56542 2681 56588
rect 2727 56542 2760 56588
rect 2668 56489 2760 56542
rect 3760 56736 3852 56789
rect 3760 56690 3793 56736
rect 3839 56690 3852 56736
rect 3760 56588 3852 56690
rect 3760 56542 3793 56588
rect 3839 56542 3852 56588
rect 3760 56489 3852 56542
rect 4168 56736 4260 56789
rect 4168 56690 4181 56736
rect 4227 56690 4260 56736
rect 4168 56588 4260 56690
rect 4168 56542 4181 56588
rect 4227 56542 4260 56588
rect 4168 56489 4260 56542
rect 5260 56736 5352 56789
rect 5260 56690 5293 56736
rect 5339 56690 5352 56736
rect 5260 56588 5352 56690
rect 5260 56542 5293 56588
rect 5339 56542 5352 56588
rect 5260 56489 5352 56542
rect 5668 56736 5760 56789
rect 5668 56690 5681 56736
rect 5727 56690 5760 56736
rect 5668 56588 5760 56690
rect 5668 56542 5681 56588
rect 5727 56542 5760 56588
rect 5668 56489 5760 56542
rect 6760 56736 6852 56789
rect 6760 56690 6793 56736
rect 6839 56690 6852 56736
rect 6760 56588 6852 56690
rect 6760 56542 6793 56588
rect 6839 56542 6852 56588
rect 6760 56489 6852 56542
rect 7168 56736 7260 56789
rect 7168 56690 7181 56736
rect 7227 56690 7260 56736
rect 7168 56588 7260 56690
rect 7168 56542 7181 56588
rect 7227 56542 7260 56588
rect 7168 56489 7260 56542
rect 8260 56736 8352 56789
rect 8260 56690 8293 56736
rect 8339 56690 8352 56736
rect 8260 56588 8352 56690
rect 8260 56542 8293 56588
rect 8339 56542 8352 56588
rect 8260 56489 8352 56542
rect 8668 56736 8760 56789
rect 8668 56690 8681 56736
rect 8727 56690 8760 56736
rect 8668 56588 8760 56690
rect 8668 56542 8681 56588
rect 8727 56542 8760 56588
rect 8668 56489 8760 56542
rect 9760 56736 9852 56789
rect 9760 56690 9793 56736
rect 9839 56690 9852 56736
rect 9760 56588 9852 56690
rect 9760 56542 9793 56588
rect 9839 56542 9852 56588
rect 9760 56489 9852 56542
rect 10168 56736 10260 56789
rect 10168 56690 10181 56736
rect 10227 56690 10260 56736
rect 10168 56588 10260 56690
rect 10168 56542 10181 56588
rect 10227 56542 10260 56588
rect 10168 56489 10260 56542
rect 11260 56736 11352 56789
rect 11260 56690 11293 56736
rect 11339 56690 11352 56736
rect 11260 56588 11352 56690
rect 11260 56542 11293 56588
rect 11339 56542 11352 56588
rect 11260 56489 11352 56542
rect 11668 56736 11760 56789
rect 11668 56690 11681 56736
rect 11727 56690 11760 56736
rect 11668 56588 11760 56690
rect 11668 56542 11681 56588
rect 11727 56542 11760 56588
rect 11668 56489 11760 56542
rect 12760 56736 12852 56789
rect 12760 56690 12793 56736
rect 12839 56690 12852 56736
rect 12760 56588 12852 56690
rect 12760 56542 12793 56588
rect 12839 56542 12852 56588
rect 12760 56489 12852 56542
rect 13168 56736 13260 56789
rect 13168 56690 13181 56736
rect 13227 56690 13260 56736
rect 13168 56588 13260 56690
rect 13168 56542 13181 56588
rect 13227 56542 13260 56588
rect 13168 56489 13260 56542
rect 14260 56736 14352 56789
rect 14260 56690 14293 56736
rect 14339 56690 14352 56736
rect 14260 56588 14352 56690
rect 14260 56542 14293 56588
rect 14339 56542 14352 56588
rect 14260 56489 14352 56542
rect 12390 43063 12482 43116
rect 12390 43017 12403 43063
rect 12449 43017 12482 43063
rect 12390 42951 12482 43017
rect 12390 42905 12403 42951
rect 12449 42905 12482 42951
rect 12390 42839 12482 42905
rect 12390 42793 12403 42839
rect 12449 42793 12482 42839
rect 12390 42727 12482 42793
rect 12390 42681 12403 42727
rect 12449 42681 12482 42727
rect 12390 42615 12482 42681
rect 12390 42569 12403 42615
rect 12449 42569 12482 42615
rect 12390 42516 12482 42569
rect 13082 43063 13174 43116
rect 13082 43017 13115 43063
rect 13161 43017 13174 43063
rect 13082 42951 13174 43017
rect 13082 42905 13115 42951
rect 13161 42905 13174 42951
rect 13082 42839 13174 42905
rect 13082 42793 13115 42839
rect 13161 42793 13174 42839
rect 13082 42727 13174 42793
rect 13082 42681 13115 42727
rect 13161 42681 13174 42727
rect 13082 42615 13174 42681
rect 13082 42569 13115 42615
rect 13161 42569 13174 42615
rect 13082 42516 13174 42569
rect 13530 43063 13622 43116
rect 13530 43017 13543 43063
rect 13589 43017 13622 43063
rect 13530 42951 13622 43017
rect 13530 42905 13543 42951
rect 13589 42905 13622 42951
rect 13530 42839 13622 42905
rect 13530 42793 13543 42839
rect 13589 42793 13622 42839
rect 13530 42727 13622 42793
rect 13530 42681 13543 42727
rect 13589 42681 13622 42727
rect 13530 42615 13622 42681
rect 13530 42569 13543 42615
rect 13589 42569 13622 42615
rect 13530 42516 13622 42569
rect 14222 43063 14314 43116
rect 14222 43017 14255 43063
rect 14301 43017 14314 43063
rect 14222 42951 14314 43017
rect 14222 42905 14255 42951
rect 14301 42905 14314 42951
rect 14222 42839 14314 42905
rect 14222 42793 14255 42839
rect 14301 42793 14314 42839
rect 14222 42727 14314 42793
rect 14222 42681 14255 42727
rect 14301 42681 14314 42727
rect 14222 42615 14314 42681
rect 14222 42569 14255 42615
rect 14301 42569 14314 42615
rect 14222 42516 14314 42569
rect 12390 42095 12482 42148
rect 12390 42049 12403 42095
rect 12449 42049 12482 42095
rect 12390 41983 12482 42049
rect 12390 41937 12403 41983
rect 12449 41937 12482 41983
rect 12390 41871 12482 41937
rect 12390 41825 12403 41871
rect 12449 41825 12482 41871
rect 12390 41759 12482 41825
rect 12390 41713 12403 41759
rect 12449 41713 12482 41759
rect 12390 41647 12482 41713
rect 12390 41601 12403 41647
rect 12449 41601 12482 41647
rect 12390 41548 12482 41601
rect 13082 42095 13174 42148
rect 13082 42049 13115 42095
rect 13161 42049 13174 42095
rect 13082 41983 13174 42049
rect 13082 41937 13115 41983
rect 13161 41937 13174 41983
rect 13082 41871 13174 41937
rect 13082 41825 13115 41871
rect 13161 41825 13174 41871
rect 13082 41759 13174 41825
rect 13082 41713 13115 41759
rect 13161 41713 13174 41759
rect 13082 41647 13174 41713
rect 13082 41601 13115 41647
rect 13161 41601 13174 41647
rect 13082 41548 13174 41601
rect 13530 42095 13622 42148
rect 13530 42049 13543 42095
rect 13589 42049 13622 42095
rect 13530 41983 13622 42049
rect 13530 41937 13543 41983
rect 13589 41937 13622 41983
rect 13530 41871 13622 41937
rect 13530 41825 13543 41871
rect 13589 41825 13622 41871
rect 13530 41759 13622 41825
rect 13530 41713 13543 41759
rect 13589 41713 13622 41759
rect 13530 41647 13622 41713
rect 13530 41601 13543 41647
rect 13589 41601 13622 41647
rect 13530 41548 13622 41601
rect 14222 42095 14314 42148
rect 14222 42049 14255 42095
rect 14301 42049 14314 42095
rect 14222 41983 14314 42049
rect 14222 41937 14255 41983
rect 14301 41937 14314 41983
rect 14222 41871 14314 41937
rect 14222 41825 14255 41871
rect 14301 41825 14314 41871
rect 14222 41759 14314 41825
rect 14222 41713 14255 41759
rect 14301 41713 14314 41759
rect 14222 41647 14314 41713
rect 14222 41601 14255 41647
rect 14301 41601 14314 41647
rect 14222 41548 14314 41601
<< polycontact >>
rect 836 56326 882 56372
rect 836 55414 882 55460
rect 1116 56326 1162 56372
rect 1116 55414 1162 55460
rect 2681 56690 2727 56736
rect 2681 56542 2727 56588
rect 3793 56690 3839 56736
rect 3793 56542 3839 56588
rect 4181 56690 4227 56736
rect 4181 56542 4227 56588
rect 5293 56690 5339 56736
rect 5293 56542 5339 56588
rect 5681 56690 5727 56736
rect 5681 56542 5727 56588
rect 6793 56690 6839 56736
rect 6793 56542 6839 56588
rect 7181 56690 7227 56736
rect 7181 56542 7227 56588
rect 8293 56690 8339 56736
rect 8293 56542 8339 56588
rect 8681 56690 8727 56736
rect 8681 56542 8727 56588
rect 9793 56690 9839 56736
rect 9793 56542 9839 56588
rect 10181 56690 10227 56736
rect 10181 56542 10227 56588
rect 11293 56690 11339 56736
rect 11293 56542 11339 56588
rect 11681 56690 11727 56736
rect 11681 56542 11727 56588
rect 12793 56690 12839 56736
rect 12793 56542 12839 56588
rect 13181 56690 13227 56736
rect 13181 56542 13227 56588
rect 14293 56690 14339 56736
rect 14293 56542 14339 56588
rect 12403 43017 12449 43063
rect 12403 42905 12449 42951
rect 12403 42793 12449 42839
rect 12403 42681 12449 42727
rect 12403 42569 12449 42615
rect 13115 43017 13161 43063
rect 13115 42905 13161 42951
rect 13115 42793 13161 42839
rect 13115 42681 13161 42727
rect 13115 42569 13161 42615
rect 13543 43017 13589 43063
rect 13543 42905 13589 42951
rect 13543 42793 13589 42839
rect 13543 42681 13589 42727
rect 13543 42569 13589 42615
rect 14255 43017 14301 43063
rect 14255 42905 14301 42951
rect 14255 42793 14301 42839
rect 14255 42681 14301 42727
rect 14255 42569 14301 42615
rect 12403 42049 12449 42095
rect 12403 41937 12449 41983
rect 12403 41825 12449 41871
rect 12403 41713 12449 41759
rect 12403 41601 12449 41647
rect 13115 42049 13161 42095
rect 13115 41937 13161 41983
rect 13115 41825 13161 41871
rect 13115 41713 13161 41759
rect 13115 41601 13161 41647
rect 13543 42049 13589 42095
rect 13543 41937 13589 41983
rect 13543 41825 13589 41871
rect 13543 41713 13589 41759
rect 13543 41601 13589 41647
rect 14255 42049 14301 42095
rect 14255 41937 14301 41983
rect 14255 41825 14301 41871
rect 14255 41713 14301 41759
rect 14255 41601 14301 41647
<< ppolyres >>
rect 779 55503 939 56283
rect 1059 55503 1219 56283
<< mvpdiode >>
rect 11458 41814 11658 41827
rect 11458 41768 11471 41814
rect 11517 41768 11599 41814
rect 11645 41768 11658 41814
rect 11458 41686 11658 41768
rect 11458 41640 11471 41686
rect 11517 41640 11599 41686
rect 11645 41640 11658 41686
rect 11458 41627 11658 41640
rect 11458 41350 11658 41363
rect 11458 41304 11471 41350
rect 11517 41304 11599 41350
rect 11645 41304 11658 41350
rect 11458 41222 11658 41304
rect 11458 41176 11471 41222
rect 11517 41176 11599 41222
rect 11645 41176 11658 41222
rect 11458 41163 11658 41176
<< mvpdiodec >>
rect 11471 41768 11517 41814
rect 11599 41768 11645 41814
rect 11471 41640 11517 41686
rect 11599 41640 11645 41686
rect 11471 41304 11517 41350
rect 11599 41304 11645 41350
rect 11471 41176 11517 41222
rect 11599 41176 11645 41222
<< metal1 >>
rect 0 52543 122 57527
rect 704 57327 14134 57339
rect 704 57171 716 57327
rect 768 57275 1486 57327
rect 1642 57275 13822 57327
rect 14082 57275 14134 57327
rect 768 57263 14134 57275
rect 768 57171 780 57263
rect 704 57159 780 57171
rect 448 56688 999 56699
rect 448 56642 459 56688
rect 975 56642 999 56688
rect 448 56631 999 56642
rect 448 56534 516 56631
rect 448 55266 459 56534
rect 505 55471 516 56534
rect 781 56372 937 56383
rect 781 56326 836 56372
rect 882 56326 937 56372
rect 781 56315 937 56326
rect 1061 56372 1217 57263
rect 2342 57202 14724 57213
rect 2342 57156 2353 57202
rect 14713 57156 14724 57202
rect 2342 57108 2522 57156
rect 2574 57108 2646 57156
rect 2698 57108 2770 57156
rect 2822 57108 2894 57156
rect 2946 57108 3018 57156
rect 3070 57108 3142 57156
rect 3194 57108 3266 57156
rect 3318 57108 3390 57156
rect 3442 57108 3514 57156
rect 3566 57108 3638 57156
rect 3690 57108 3762 57156
rect 3814 57108 3886 57156
rect 3938 57108 4010 57156
rect 4062 57108 4134 57156
rect 4186 57108 4258 57156
rect 4310 57108 4382 57156
rect 4434 57108 4506 57156
rect 4558 57108 4630 57156
rect 4682 57108 4754 57156
rect 4806 57108 4878 57156
rect 4930 57108 5002 57156
rect 5054 57108 5126 57156
rect 5178 57108 5250 57156
rect 5302 57108 5374 57156
rect 5426 57108 5498 57156
rect 5550 57108 5622 57156
rect 5674 57108 5746 57156
rect 5798 57108 5870 57156
rect 5922 57108 5994 57156
rect 6046 57108 6118 57156
rect 6170 57108 6242 57156
rect 6294 57108 6366 57156
rect 6418 57108 6490 57156
rect 6542 57108 6614 57156
rect 6666 57108 6738 57156
rect 6790 57108 6862 57156
rect 6914 57108 6986 57156
rect 7038 57108 7110 57156
rect 7162 57108 7234 57156
rect 7286 57108 7358 57156
rect 7410 57108 7482 57156
rect 7534 57108 7606 57156
rect 7658 57108 7730 57156
rect 7782 57108 7854 57156
rect 7906 57108 7978 57156
rect 8030 57108 8102 57156
rect 8154 57108 8226 57156
rect 8278 57108 8350 57156
rect 8402 57108 8474 57156
rect 8526 57108 8598 57156
rect 8650 57108 8722 57156
rect 8774 57108 8846 57156
rect 8898 57108 8970 57156
rect 9022 57108 9094 57156
rect 9146 57108 9218 57156
rect 9270 57108 9342 57156
rect 9394 57108 9466 57156
rect 9518 57108 9590 57156
rect 9642 57108 9714 57156
rect 9766 57108 9838 57156
rect 9890 57108 9962 57156
rect 10014 57108 10086 57156
rect 10138 57108 10210 57156
rect 10262 57108 10334 57156
rect 10386 57108 10458 57156
rect 10510 57108 10582 57156
rect 10634 57108 10706 57156
rect 10758 57108 10830 57156
rect 10882 57108 10954 57156
rect 11006 57108 11078 57156
rect 11130 57108 11202 57156
rect 11254 57108 11326 57156
rect 11378 57108 11450 57156
rect 11502 57108 11574 57156
rect 11626 57108 11698 57156
rect 11750 57108 11822 57156
rect 11874 57108 11946 57156
rect 11998 57108 12070 57156
rect 12122 57108 12194 57156
rect 12246 57108 12318 57156
rect 12370 57108 12442 57156
rect 12494 57108 12566 57156
rect 12618 57108 12690 57156
rect 12742 57108 12814 57156
rect 12866 57108 12938 57156
rect 12990 57108 13062 57156
rect 13114 57108 13186 57156
rect 13238 57108 13310 57156
rect 13362 57108 13434 57156
rect 13486 57108 13558 57156
rect 13610 57108 14724 57156
rect 2342 57038 14724 57108
rect 1273 56688 1550 56699
rect 1273 56642 1305 56688
rect 1539 56642 1550 56688
rect 1273 56631 1550 56642
rect 1061 56326 1116 56372
rect 1162 56326 1217 56372
rect 1061 56315 1217 56326
rect 1482 56534 1550 56631
rect 861 56225 937 56315
rect 1482 56300 1493 56534
rect 1539 56300 1550 56534
rect 1482 56285 1550 56300
rect 2342 56240 2353 57038
rect 2399 57036 14667 57038
rect 2399 56984 2522 57036
rect 2574 56984 2646 57036
rect 2698 56984 2770 57036
rect 2822 56984 2894 57036
rect 2946 56984 3018 57036
rect 3070 56984 3142 57036
rect 3194 56984 3266 57036
rect 3318 56984 3390 57036
rect 3442 56984 3514 57036
rect 3566 56984 3638 57036
rect 3690 56984 3762 57036
rect 3814 56984 3886 57036
rect 3938 56984 4010 57036
rect 4062 56984 4134 57036
rect 4186 56984 4258 57036
rect 4310 56984 4382 57036
rect 4434 56984 4506 57036
rect 4558 56984 4630 57036
rect 4682 56984 4754 57036
rect 4806 56984 4878 57036
rect 4930 56984 5002 57036
rect 5054 56984 5126 57036
rect 5178 56984 5250 57036
rect 5302 56984 5374 57036
rect 5426 56984 5498 57036
rect 5550 56984 5622 57036
rect 5674 56984 5746 57036
rect 5798 56984 5870 57036
rect 5922 56984 5994 57036
rect 6046 56984 6118 57036
rect 6170 56984 6242 57036
rect 6294 56984 6366 57036
rect 6418 56984 6490 57036
rect 6542 56984 6614 57036
rect 6666 56984 6738 57036
rect 6790 56984 6862 57036
rect 6914 56984 6986 57036
rect 7038 56984 7110 57036
rect 7162 56984 7234 57036
rect 7286 56984 7358 57036
rect 7410 56984 7482 57036
rect 7534 56984 7606 57036
rect 7658 56984 7730 57036
rect 7782 56984 7854 57036
rect 7906 56984 7978 57036
rect 8030 56984 8102 57036
rect 8154 56984 8226 57036
rect 8278 56984 8350 57036
rect 8402 56984 8474 57036
rect 8526 56984 8598 57036
rect 8650 56984 8722 57036
rect 8774 56984 8846 57036
rect 8898 56984 8970 57036
rect 9022 56984 9094 57036
rect 9146 56984 9218 57036
rect 9270 56984 9342 57036
rect 9394 56984 9466 57036
rect 9518 56984 9590 57036
rect 9642 56984 9714 57036
rect 9766 56984 9838 57036
rect 9890 56984 9962 57036
rect 10014 56984 10086 57036
rect 10138 56984 10210 57036
rect 10262 56984 10334 57036
rect 10386 56984 10458 57036
rect 10510 56984 10582 57036
rect 10634 56984 10706 57036
rect 10758 56984 10830 57036
rect 10882 56984 10954 57036
rect 11006 56984 11078 57036
rect 11130 56984 11202 57036
rect 11254 56984 11326 57036
rect 11378 56984 11450 57036
rect 11502 56984 11574 57036
rect 11626 56984 11698 57036
rect 11750 56984 11822 57036
rect 11874 56984 11946 57036
rect 11998 56984 12070 57036
rect 12122 56984 12194 57036
rect 12246 56984 12318 57036
rect 12370 56984 12442 57036
rect 12494 56984 12566 57036
rect 12618 56984 12690 57036
rect 12742 56984 12814 57036
rect 12866 56984 12938 57036
rect 12990 56984 13062 57036
rect 13114 56984 13186 57036
rect 13238 56984 13310 57036
rect 13362 56984 13434 57036
rect 13486 56984 13558 57036
rect 13610 56984 14667 57036
rect 2399 56912 14667 56984
rect 2399 56860 2522 56912
rect 2574 56860 2646 56912
rect 2698 56860 2770 56912
rect 2822 56864 2894 56912
rect 2946 56864 3018 56912
rect 3070 56864 3142 56912
rect 3194 56864 3266 56912
rect 3318 56864 3390 56912
rect 3442 56864 3514 56912
rect 3566 56864 3638 56912
rect 3690 56864 3762 56912
rect 3723 56860 3762 56864
rect 3814 56860 3886 56912
rect 3938 56860 4010 56912
rect 4062 56860 4134 56912
rect 4186 56860 4258 56912
rect 4310 56864 4382 56912
rect 4434 56864 4506 56912
rect 4558 56864 4630 56912
rect 4682 56864 4754 56912
rect 4806 56864 4878 56912
rect 4930 56864 5002 56912
rect 5054 56864 5126 56912
rect 5178 56864 5250 56912
rect 5223 56860 5250 56864
rect 5302 56860 5374 56912
rect 5426 56860 5498 56912
rect 5550 56860 5622 56912
rect 5674 56860 5746 56912
rect 5798 56864 5870 56912
rect 5922 56864 5994 56912
rect 6046 56864 6118 56912
rect 6170 56864 6242 56912
rect 6294 56864 6366 56912
rect 6418 56864 6490 56912
rect 6542 56864 6614 56912
rect 6666 56864 6738 56912
rect 6723 56860 6738 56864
rect 6790 56860 6862 56912
rect 6914 56860 6986 56912
rect 7038 56860 7110 56912
rect 7162 56860 7234 56912
rect 7286 56864 7358 56912
rect 7410 56864 7482 56912
rect 7534 56864 7606 56912
rect 7658 56864 7730 56912
rect 7782 56864 7854 56912
rect 7906 56864 7978 56912
rect 8030 56864 8102 56912
rect 8154 56864 8226 56912
rect 7286 56860 7297 56864
rect 8223 56860 8226 56864
rect 8278 56860 8350 56912
rect 8402 56860 8474 56912
rect 8526 56860 8598 56912
rect 8650 56860 8722 56912
rect 8774 56864 8846 56912
rect 8898 56864 8970 56912
rect 9022 56864 9094 56912
rect 9146 56864 9218 56912
rect 9270 56864 9342 56912
rect 9394 56864 9466 56912
rect 9518 56864 9590 56912
rect 9642 56864 9714 56912
rect 8774 56860 8797 56864
rect 9766 56860 9838 56912
rect 9890 56860 9962 56912
rect 10014 56860 10086 56912
rect 10138 56860 10210 56912
rect 10262 56864 10334 56912
rect 10386 56864 10458 56912
rect 10510 56864 10582 56912
rect 10634 56864 10706 56912
rect 10758 56864 10830 56912
rect 10882 56864 10954 56912
rect 11006 56864 11078 56912
rect 11130 56864 11202 56912
rect 10262 56860 10297 56864
rect 11254 56860 11326 56912
rect 11378 56860 11450 56912
rect 11502 56860 11574 56912
rect 11626 56860 11698 56912
rect 11750 56864 11822 56912
rect 11874 56864 11946 56912
rect 11998 56864 12070 56912
rect 12122 56864 12194 56912
rect 12246 56864 12318 56912
rect 12370 56864 12442 56912
rect 12494 56864 12566 56912
rect 12618 56864 12690 56912
rect 11750 56860 11797 56864
rect 12742 56860 12814 56912
rect 12866 56860 12938 56912
rect 12990 56860 13062 56912
rect 13114 56860 13186 56912
rect 13238 56864 13310 56912
rect 13362 56864 13434 56912
rect 13486 56864 13558 56912
rect 13610 56864 14667 56912
rect 13238 56860 13297 56864
rect 2399 56818 2797 56860
rect 3723 56818 4297 56860
rect 5223 56818 5797 56860
rect 6723 56818 7297 56860
rect 8223 56818 8797 56860
rect 9723 56818 10297 56860
rect 11223 56818 11797 56860
rect 12723 56818 13297 56860
rect 14223 56818 14667 56864
rect 2399 56807 14667 56818
rect 2399 56471 2610 56807
rect 2670 56736 3850 56747
rect 2670 56690 2681 56736
rect 2727 56715 3793 56736
rect 2670 56588 2682 56690
rect 2670 56542 2681 56588
rect 2838 56559 3682 56715
rect 3839 56690 3850 56736
rect 3838 56588 3850 56690
rect 2727 56542 3793 56559
rect 3839 56542 3850 56588
rect 2670 56531 3850 56542
rect 3910 56471 4110 56807
rect 4170 56736 5350 56747
rect 4170 56690 4181 56736
rect 4227 56715 5293 56736
rect 4170 56588 4182 56690
rect 4170 56542 4181 56588
rect 4338 56559 5182 56715
rect 5339 56690 5350 56736
rect 5338 56588 5350 56690
rect 4227 56542 5293 56559
rect 5339 56542 5350 56588
rect 4170 56531 5350 56542
rect 5410 56471 5610 56807
rect 5670 56736 6850 56747
rect 5670 56690 5681 56736
rect 5727 56715 6793 56736
rect 5670 56588 5682 56690
rect 5670 56542 5681 56588
rect 5838 56559 6682 56715
rect 6839 56690 6850 56736
rect 6838 56588 6850 56690
rect 5727 56542 6793 56559
rect 6839 56542 6850 56588
rect 5670 56531 6850 56542
rect 6910 56471 7110 56807
rect 7170 56736 8350 56747
rect 7170 56690 7181 56736
rect 7227 56715 8293 56736
rect 7170 56588 7182 56690
rect 7170 56542 7181 56588
rect 7338 56559 8182 56715
rect 8339 56690 8350 56736
rect 8338 56588 8350 56690
rect 7227 56542 8293 56559
rect 8339 56542 8350 56588
rect 7170 56531 8350 56542
rect 8410 56471 8610 56807
rect 8670 56736 9850 56747
rect 8670 56690 8681 56736
rect 8727 56715 9793 56736
rect 8670 56588 8682 56690
rect 8670 56542 8681 56588
rect 8838 56559 9682 56715
rect 9839 56690 9850 56736
rect 9838 56588 9850 56690
rect 8727 56542 9793 56559
rect 9839 56542 9850 56588
rect 8670 56531 9850 56542
rect 9910 56471 10110 56807
rect 10170 56736 11350 56747
rect 10170 56690 10181 56736
rect 10227 56715 11293 56736
rect 10170 56588 10182 56690
rect 10170 56542 10181 56588
rect 10338 56559 11182 56715
rect 11339 56690 11350 56736
rect 11338 56588 11350 56690
rect 10227 56542 11293 56559
rect 11339 56542 11350 56588
rect 10170 56531 11350 56542
rect 11410 56471 11610 56807
rect 11670 56736 12850 56747
rect 11670 56690 11681 56736
rect 11727 56715 12793 56736
rect 11670 56588 11682 56690
rect 11670 56542 11681 56588
rect 11838 56559 12682 56715
rect 12839 56690 12850 56736
rect 12838 56588 12850 56690
rect 11727 56542 12793 56559
rect 12839 56542 12850 56588
rect 11670 56531 12850 56542
rect 12910 56471 13110 56807
rect 13170 56736 14560 56747
rect 13170 56690 13181 56736
rect 13227 56715 14293 56736
rect 13338 56690 14293 56715
rect 14339 56715 14560 56736
rect 14339 56690 14392 56715
rect 13170 56588 13182 56690
rect 13338 56588 14392 56690
rect 13170 56542 13181 56588
rect 13338 56559 14293 56588
rect 13227 56542 14293 56559
rect 14339 56559 14392 56588
rect 14548 56559 14560 56715
rect 14339 56542 14560 56559
rect 13170 56531 14560 56542
rect 14656 56471 14667 56807
rect 2399 56460 14667 56471
rect 2399 56418 2797 56460
rect 3723 56418 4297 56460
rect 5223 56418 5797 56460
rect 6723 56418 7297 56460
rect 8223 56418 8797 56460
rect 9723 56418 10297 56460
rect 11223 56418 11797 56460
rect 12723 56418 13297 56460
rect 2399 56366 2522 56418
rect 2574 56366 2646 56418
rect 2698 56366 2770 56418
rect 3723 56414 3762 56418
rect 2822 56366 2894 56414
rect 2946 56366 3018 56414
rect 3070 56366 3142 56414
rect 3194 56366 3266 56414
rect 3318 56366 3390 56414
rect 3442 56366 3514 56414
rect 3566 56366 3638 56414
rect 3690 56366 3762 56414
rect 3814 56366 3886 56418
rect 3938 56366 4010 56418
rect 4062 56366 4134 56418
rect 4186 56366 4258 56418
rect 5223 56414 5250 56418
rect 4310 56366 4382 56414
rect 4434 56366 4506 56414
rect 4558 56366 4630 56414
rect 4682 56366 4754 56414
rect 4806 56366 4878 56414
rect 4930 56366 5002 56414
rect 5054 56366 5126 56414
rect 5178 56366 5250 56414
rect 5302 56366 5374 56418
rect 5426 56366 5498 56418
rect 5550 56366 5622 56418
rect 5674 56366 5746 56418
rect 6723 56414 6738 56418
rect 5798 56366 5870 56414
rect 5922 56366 5994 56414
rect 6046 56366 6118 56414
rect 6170 56366 6242 56414
rect 6294 56366 6366 56414
rect 6418 56366 6490 56414
rect 6542 56366 6614 56414
rect 6666 56366 6738 56414
rect 6790 56366 6862 56418
rect 6914 56366 6986 56418
rect 7038 56366 7110 56418
rect 7162 56366 7234 56418
rect 7286 56414 7297 56418
rect 8223 56414 8226 56418
rect 7286 56366 7358 56414
rect 7410 56366 7482 56414
rect 7534 56366 7606 56414
rect 7658 56366 7730 56414
rect 7782 56366 7854 56414
rect 7906 56366 7978 56414
rect 8030 56366 8102 56414
rect 8154 56366 8226 56414
rect 8278 56366 8350 56418
rect 8402 56366 8474 56418
rect 8526 56366 8598 56418
rect 8650 56366 8722 56418
rect 8774 56414 8797 56418
rect 8774 56366 8846 56414
rect 8898 56366 8970 56414
rect 9022 56366 9094 56414
rect 9146 56366 9218 56414
rect 9270 56366 9342 56414
rect 9394 56366 9466 56414
rect 9518 56366 9590 56414
rect 9642 56366 9714 56414
rect 9766 56366 9838 56418
rect 9890 56366 9962 56418
rect 10014 56366 10086 56418
rect 10138 56366 10210 56418
rect 10262 56414 10297 56418
rect 10262 56366 10334 56414
rect 10386 56366 10458 56414
rect 10510 56366 10582 56414
rect 10634 56366 10706 56414
rect 10758 56366 10830 56414
rect 10882 56366 10954 56414
rect 11006 56366 11078 56414
rect 11130 56366 11202 56414
rect 11254 56366 11326 56418
rect 11378 56366 11450 56418
rect 11502 56366 11574 56418
rect 11626 56366 11698 56418
rect 11750 56414 11797 56418
rect 11750 56366 11822 56414
rect 11874 56366 11946 56414
rect 11998 56366 12070 56414
rect 12122 56366 12194 56414
rect 12246 56366 12318 56414
rect 12370 56366 12442 56414
rect 12494 56366 12566 56414
rect 12618 56366 12690 56414
rect 12742 56366 12814 56418
rect 12866 56366 12938 56418
rect 12990 56366 13062 56418
rect 13114 56366 13186 56418
rect 13238 56414 13297 56418
rect 14223 56414 14667 56460
rect 13238 56366 13310 56414
rect 13362 56366 13434 56414
rect 13486 56366 13558 56414
rect 13610 56366 14667 56414
rect 2399 56294 14667 56366
rect 2399 56242 2522 56294
rect 2574 56242 2646 56294
rect 2698 56242 2770 56294
rect 2822 56242 2894 56294
rect 2946 56242 3018 56294
rect 3070 56242 3142 56294
rect 3194 56242 3266 56294
rect 3318 56242 3390 56294
rect 3442 56242 3514 56294
rect 3566 56242 3638 56294
rect 3690 56242 3762 56294
rect 3814 56242 3886 56294
rect 3938 56242 4010 56294
rect 4062 56242 4134 56294
rect 4186 56242 4258 56294
rect 4310 56242 4382 56294
rect 4434 56242 4506 56294
rect 4558 56242 4630 56294
rect 4682 56242 4754 56294
rect 4806 56242 4878 56294
rect 4930 56242 5002 56294
rect 5054 56242 5126 56294
rect 5178 56242 5250 56294
rect 5302 56242 5374 56294
rect 5426 56242 5498 56294
rect 5550 56242 5622 56294
rect 5674 56242 5746 56294
rect 5798 56242 5870 56294
rect 5922 56242 5994 56294
rect 6046 56242 6118 56294
rect 6170 56242 6242 56294
rect 6294 56242 6366 56294
rect 6418 56242 6490 56294
rect 6542 56242 6614 56294
rect 6666 56242 6738 56294
rect 6790 56242 6862 56294
rect 6914 56242 6986 56294
rect 7038 56242 7110 56294
rect 7162 56242 7234 56294
rect 7286 56242 7358 56294
rect 7410 56242 7482 56294
rect 7534 56242 7606 56294
rect 7658 56242 7730 56294
rect 7782 56242 7854 56294
rect 7906 56242 7978 56294
rect 8030 56242 8102 56294
rect 8154 56242 8226 56294
rect 8278 56242 8350 56294
rect 8402 56242 8474 56294
rect 8526 56242 8598 56294
rect 8650 56242 8722 56294
rect 8774 56242 8846 56294
rect 8898 56242 8970 56294
rect 9022 56242 9094 56294
rect 9146 56242 9218 56294
rect 9270 56242 9342 56294
rect 9394 56242 9466 56294
rect 9518 56242 9590 56294
rect 9642 56242 9714 56294
rect 9766 56242 9838 56294
rect 9890 56242 9962 56294
rect 10014 56242 10086 56294
rect 10138 56242 10210 56294
rect 10262 56242 10334 56294
rect 10386 56242 10458 56294
rect 10510 56242 10582 56294
rect 10634 56242 10706 56294
rect 10758 56242 10830 56294
rect 10882 56242 10954 56294
rect 11006 56242 11078 56294
rect 11130 56242 11202 56294
rect 11254 56242 11326 56294
rect 11378 56242 11450 56294
rect 11502 56242 11574 56294
rect 11626 56242 11698 56294
rect 11750 56242 11822 56294
rect 11874 56242 11946 56294
rect 11998 56242 12070 56294
rect 12122 56242 12194 56294
rect 12246 56242 12318 56294
rect 12370 56242 12442 56294
rect 12494 56242 12566 56294
rect 12618 56242 12690 56294
rect 12742 56242 12814 56294
rect 12866 56242 12938 56294
rect 12990 56242 13062 56294
rect 13114 56242 13186 56294
rect 13238 56242 13310 56294
rect 13362 56242 13434 56294
rect 13486 56242 13558 56294
rect 13610 56242 14667 56294
rect 2399 56240 14667 56242
rect 14713 56240 14724 57038
rect 861 56149 1827 56225
rect 1482 56064 1550 56089
rect 1482 55548 1493 56064
rect 1539 55548 1550 56064
rect 1751 55723 1827 56149
rect 2342 56170 14724 56240
rect 2342 56122 2522 56170
rect 2574 56122 2646 56170
rect 2698 56122 2770 56170
rect 2822 56122 2894 56170
rect 2946 56122 3018 56170
rect 3070 56122 3142 56170
rect 3194 56122 3266 56170
rect 3318 56122 3390 56170
rect 3442 56122 3514 56170
rect 3566 56122 3638 56170
rect 3690 56122 3762 56170
rect 3814 56122 3886 56170
rect 3938 56122 4010 56170
rect 4062 56122 4134 56170
rect 4186 56122 4258 56170
rect 4310 56122 4382 56170
rect 4434 56122 4506 56170
rect 4558 56122 4630 56170
rect 4682 56122 4754 56170
rect 4806 56122 4878 56170
rect 4930 56122 5002 56170
rect 5054 56122 5126 56170
rect 5178 56122 5250 56170
rect 5302 56122 5374 56170
rect 5426 56122 5498 56170
rect 5550 56122 5622 56170
rect 5674 56122 5746 56170
rect 5798 56122 5870 56170
rect 5922 56122 5994 56170
rect 6046 56122 6118 56170
rect 6170 56122 6242 56170
rect 6294 56122 6366 56170
rect 6418 56122 6490 56170
rect 6542 56122 6614 56170
rect 6666 56122 6738 56170
rect 6790 56122 6862 56170
rect 6914 56122 6986 56170
rect 7038 56122 7110 56170
rect 7162 56122 7234 56170
rect 7286 56122 7358 56170
rect 7410 56122 7482 56170
rect 7534 56122 7606 56170
rect 7658 56122 7730 56170
rect 7782 56122 7854 56170
rect 7906 56122 7978 56170
rect 8030 56122 8102 56170
rect 8154 56122 8226 56170
rect 8278 56122 8350 56170
rect 8402 56122 8474 56170
rect 8526 56122 8598 56170
rect 8650 56122 8722 56170
rect 8774 56122 8846 56170
rect 8898 56122 8970 56170
rect 9022 56122 9094 56170
rect 9146 56122 9218 56170
rect 9270 56122 9342 56170
rect 9394 56122 9466 56170
rect 9518 56122 9590 56170
rect 9642 56122 9714 56170
rect 9766 56122 9838 56170
rect 9890 56122 9962 56170
rect 10014 56122 10086 56170
rect 10138 56122 10210 56170
rect 10262 56122 10334 56170
rect 10386 56122 10458 56170
rect 10510 56122 10582 56170
rect 10634 56122 10706 56170
rect 10758 56122 10830 56170
rect 10882 56122 10954 56170
rect 11006 56122 11078 56170
rect 11130 56122 11202 56170
rect 11254 56122 11326 56170
rect 11378 56122 11450 56170
rect 11502 56122 11574 56170
rect 11626 56122 11698 56170
rect 11750 56122 11822 56170
rect 11874 56122 11946 56170
rect 11998 56122 12070 56170
rect 12122 56122 12194 56170
rect 12246 56122 12318 56170
rect 12370 56122 12442 56170
rect 12494 56122 12566 56170
rect 12618 56122 12690 56170
rect 12742 56122 12814 56170
rect 12866 56122 12938 56170
rect 12990 56122 13062 56170
rect 13114 56122 13186 56170
rect 13238 56122 13310 56170
rect 13362 56122 13434 56170
rect 13486 56122 13558 56170
rect 13610 56122 14724 56170
rect 2342 56076 2353 56122
rect 14713 56076 14724 56122
rect 2342 56065 14724 56076
rect 3500 55837 4096 55849
rect 3500 55785 3512 55837
rect 4084 55785 4096 55837
rect 3500 55773 4096 55785
rect 8030 55829 8106 55841
rect 4938 55758 5014 55770
rect 4750 55729 4826 55741
rect 1751 55711 2385 55723
rect 1751 55647 2321 55711
rect 1482 55520 1550 55548
rect 2309 55555 2321 55647
rect 2373 55555 2385 55711
rect 2309 55543 2385 55555
rect 2593 55471 2773 55475
rect 505 55460 937 55471
rect 505 55414 836 55460
rect 882 55414 937 55460
rect 505 55403 937 55414
rect 1061 55463 2773 55471
rect 1061 55460 2605 55463
rect 1061 55414 1116 55460
rect 1162 55414 2605 55460
rect 1061 55411 2605 55414
rect 2761 55411 2773 55463
rect 1061 55403 2773 55411
rect 505 55266 516 55403
rect 2593 55399 2773 55403
rect 448 55169 516 55266
rect 1482 55312 1550 55345
rect 1482 55266 1493 55312
rect 1539 55266 1550 55312
rect 1482 55169 1550 55266
rect 184 55158 1550 55169
rect 184 55112 459 55158
rect 1539 55112 1550 55158
rect 184 55101 1550 55112
rect 184 55095 921 55101
rect 184 55043 234 55095
rect 286 55043 358 55095
rect 410 55043 482 55095
rect 534 55043 921 55095
rect 184 54971 921 55043
rect 184 54919 234 54971
rect 286 54919 358 54971
rect 410 54919 482 54971
rect 534 54919 921 54971
rect 184 54847 921 54919
rect 184 54795 234 54847
rect 286 54795 358 54847
rect 410 54795 482 54847
rect 534 54795 921 54847
rect 4750 54845 4762 55729
rect 4814 54845 4826 55729
rect 4938 54978 4950 55758
rect 5002 54978 5014 55758
rect 4938 54966 5014 54978
rect 5426 55767 5502 55779
rect 5426 54987 5438 55767
rect 5490 54987 5502 55767
rect 5426 54975 5502 54987
rect 5914 55767 5990 55779
rect 5914 54987 5926 55767
rect 5978 54987 5990 55767
rect 5914 54975 5990 54987
rect 6096 55729 6172 55773
rect 4750 54833 4826 54845
rect 6096 54845 6108 55729
rect 6160 54845 6172 55729
rect 6278 55767 6354 55779
rect 6278 54987 6290 55767
rect 6342 54987 6354 55767
rect 6278 54975 6354 54987
rect 6766 55767 6842 55779
rect 6766 54987 6778 55767
rect 6830 54987 6842 55767
rect 6766 54975 6842 54987
rect 7254 55767 7330 55779
rect 7254 54987 7266 55767
rect 7318 54987 7330 55767
rect 7254 54975 7330 54987
rect 7442 55729 7518 55741
rect 6096 54833 6172 54845
rect 7442 54845 7454 55729
rect 7506 54845 7518 55729
rect 7442 54833 7518 54845
rect 8030 54841 8042 55829
rect 8094 54841 8106 55829
rect 8030 54829 8106 54841
rect 8499 55829 8575 55841
rect 8499 54841 8511 55829
rect 8563 54841 8575 55829
rect 8499 54829 8575 54841
rect 8714 55829 8790 55841
rect 8714 54841 8726 55829
rect 8778 54841 8790 55829
rect 8714 54829 8790 54841
rect 8937 55829 9013 55841
rect 8937 54841 8949 55829
rect 9001 54841 9013 55829
rect 8937 54829 9013 54841
rect 9406 55829 9482 55841
rect 9406 54841 9418 55829
rect 9470 54841 9482 55829
rect 10182 55767 10258 55779
rect 9406 54829 9482 54841
rect 9994 55729 10070 55741
rect 9994 54845 10006 55729
rect 10058 54845 10070 55729
rect 10182 54987 10194 55767
rect 10246 54987 10258 55767
rect 10182 54975 10258 54987
rect 10670 55767 10746 55779
rect 10670 54987 10682 55767
rect 10734 54987 10746 55767
rect 10670 54975 10746 54987
rect 11158 55767 11234 55779
rect 11158 54987 11170 55767
rect 11222 54987 11234 55767
rect 11158 54975 11234 54987
rect 11340 55729 11416 55773
rect 9994 54833 10070 54845
rect 11340 54845 11352 55729
rect 11404 54845 11416 55729
rect 11522 55767 11598 55779
rect 11522 54987 11534 55767
rect 11586 54987 11598 55767
rect 11522 54975 11598 54987
rect 12010 55767 12086 55779
rect 12010 54987 12022 55767
rect 12074 54987 12086 55767
rect 12010 54975 12086 54987
rect 12498 55767 12574 55779
rect 12498 54987 12510 55767
rect 12562 54987 12574 55767
rect 12498 54975 12574 54987
rect 12686 55729 12762 55741
rect 11340 54833 11416 54845
rect 12686 54845 12698 55729
rect 12750 54845 12762 55729
rect 12686 54833 12762 54845
rect 13274 55729 13350 55741
rect 13274 54845 13286 55729
rect 13338 54845 13350 55729
rect 13274 54833 13350 54845
rect 184 54724 921 54795
rect 3470 54371 3546 54383
rect 184 54186 921 54260
rect 184 54134 234 54186
rect 286 54134 358 54186
rect 410 54134 482 54186
rect 534 54134 921 54186
rect 184 54062 921 54134
rect 184 54010 234 54062
rect 286 54010 358 54062
rect 410 54010 482 54062
rect 534 54010 921 54062
rect 184 53938 921 54010
rect 184 53886 234 53938
rect 286 53886 358 53938
rect 410 53886 482 53938
rect 534 53886 921 53938
rect 184 53815 921 53886
rect 3470 53383 3482 54371
rect 3534 53383 3546 54371
rect 8718 54371 8794 54383
rect 6096 54267 6172 54279
rect 3470 53371 3546 53383
rect 4162 54163 4238 54175
rect 4162 53383 4174 54163
rect 4226 53383 4238 54163
rect 4162 53371 4238 53383
rect 4750 54163 4826 54175
rect 4750 53383 4762 54163
rect 4814 53383 4826 54163
rect 4938 54002 5014 54014
rect 4938 53430 4950 54002
rect 5002 53430 5014 54002
rect 4938 53418 5014 53430
rect 5426 54002 5502 54014
rect 5426 53430 5438 54002
rect 5490 53430 5502 54002
rect 5426 53418 5502 53430
rect 5914 54002 5990 54014
rect 5914 53430 5926 54002
rect 5978 53430 5990 54002
rect 5914 53418 5990 53430
rect 4750 53371 4826 53383
rect 6096 53383 6108 54267
rect 6160 53383 6172 54267
rect 7442 54163 7518 54175
rect 6278 54002 6354 54014
rect 6278 53430 6290 54002
rect 6342 53430 6354 54002
rect 6278 53418 6354 53430
rect 6766 54002 6842 54014
rect 6766 53430 6778 54002
rect 6830 53430 6842 54002
rect 6766 53418 6842 53430
rect 7254 54002 7330 54014
rect 7254 53430 7266 54002
rect 7318 53430 7330 54002
rect 7254 53418 7330 53430
rect 6096 53371 6172 53383
rect 7442 53383 7454 54163
rect 7506 53383 7518 54163
rect 7442 53371 7518 53383
rect 8030 54163 8106 54175
rect 8030 53383 8042 54163
rect 8094 53383 8106 54163
rect 8030 53371 8106 53383
rect 8718 53383 8730 54371
rect 8782 53383 8794 54371
rect 11340 54267 11416 54279
rect 8718 53371 8794 53383
rect 9994 54163 10070 54175
rect 9994 53383 10006 54163
rect 10058 53383 10070 54163
rect 10182 54002 10258 54014
rect 10182 53430 10194 54002
rect 10246 53430 10258 54002
rect 10182 53418 10258 53430
rect 10670 54002 10746 54014
rect 10670 53430 10682 54002
rect 10734 53430 10746 54002
rect 10670 53418 10746 53430
rect 11158 54002 11234 54014
rect 11158 53430 11170 54002
rect 11222 53430 11234 54002
rect 11158 53418 11234 53430
rect 9994 53371 10070 53383
rect 11340 53383 11352 54267
rect 11404 53383 11416 54267
rect 12686 54163 12762 54175
rect 11522 54002 11598 54014
rect 11522 53430 11534 54002
rect 11586 53430 11598 54002
rect 11522 53418 11598 53430
rect 12010 54002 12086 54014
rect 12010 53430 12022 54002
rect 12074 53430 12086 54002
rect 12010 53418 12086 53430
rect 12498 54002 12574 54014
rect 12498 53430 12510 54002
rect 12562 53430 12574 54002
rect 12498 53418 12574 53430
rect 11340 53371 11416 53383
rect 12686 53383 12698 54163
rect 12750 53383 12762 54163
rect 12686 53371 12762 53383
rect 13274 54163 13350 54175
rect 13274 53383 13286 54163
rect 13338 53383 13350 54163
rect 13274 53371 13350 53383
rect 704 53007 3863 53019
rect 704 52955 722 53007
rect 1086 52955 3378 53007
rect 3534 52955 3695 53007
rect 3851 52955 3863 53007
rect 704 52943 3863 52955
rect 4734 52679 5226 52691
rect 4734 52627 4746 52679
rect 5214 52627 5226 52679
rect 4734 52615 5226 52627
rect 6438 52679 6930 52691
rect 6438 52627 6450 52679
rect 6918 52627 6930 52679
rect 6438 52615 6930 52627
rect 7254 52679 7434 52691
rect 7254 52627 7266 52679
rect 7422 52627 7434 52679
rect 7254 52615 7434 52627
rect 0 51243 58 52543
rect 110 51243 122 52543
rect 0 38143 122 51243
rect 14942 52491 15064 57557
rect 14942 51295 14954 52491
rect 15006 51295 15064 52491
rect 1852 50269 6816 50281
rect 1852 50217 1864 50269
rect 6804 50217 6816 50269
rect 1852 50205 6816 50217
rect 7720 50269 8108 50281
rect 7720 50217 7732 50269
rect 8096 50217 8108 50269
rect 7720 50205 8108 50217
rect 8422 50269 8810 50281
rect 8422 50217 8434 50269
rect 8798 50217 8810 50269
rect 8422 50205 8810 50217
rect 4632 49424 4956 49436
rect 4632 49372 4644 49424
rect 4696 49372 4768 49424
rect 4820 49372 4892 49424
rect 4944 49372 4956 49424
rect 4632 49300 4956 49372
rect 4632 49248 4644 49300
rect 4696 49248 4768 49300
rect 4820 49248 4892 49300
rect 4944 49248 4956 49300
rect 4632 49176 4956 49248
rect 4632 49124 4644 49176
rect 4696 49124 4768 49176
rect 4820 49124 4892 49176
rect 4944 49124 4956 49176
rect 5519 49398 5907 49410
rect 5519 49138 5531 49398
rect 5895 49138 5907 49398
rect 5519 49126 5907 49138
rect 6422 49398 6810 49410
rect 6422 49138 6434 49398
rect 6798 49138 6810 49398
rect 6422 49126 6810 49138
rect 7720 49398 8108 49410
rect 7720 49138 7732 49398
rect 8096 49138 8108 49398
rect 7720 49126 8108 49138
rect 8422 49398 8810 49410
rect 8422 49138 8434 49398
rect 8798 49138 8810 49398
rect 8422 49126 8810 49138
rect 10782 49360 10858 49372
rect 4632 49052 4956 49124
rect 4632 49000 4644 49052
rect 4696 49000 4768 49052
rect 4820 49000 4892 49052
rect 4944 49000 4956 49052
rect 4632 48928 4956 49000
rect 4632 48876 4644 48928
rect 4696 48876 4768 48928
rect 4820 48876 4892 48928
rect 4944 48876 4956 48928
rect 4632 48804 4956 48876
rect 4632 48752 4644 48804
rect 4696 48752 4768 48804
rect 4820 48752 4892 48804
rect 4944 48752 4956 48804
rect 4632 48680 4956 48752
rect 4632 48628 4644 48680
rect 4696 48628 4768 48680
rect 4820 48628 4892 48680
rect 4944 48628 4956 48680
rect 4632 48556 4956 48628
rect 4632 48504 4644 48556
rect 4696 48504 4768 48556
rect 4820 48504 4892 48556
rect 4944 48504 4956 48556
rect 4632 48432 4956 48504
rect 4632 48380 4644 48432
rect 4696 48380 4768 48432
rect 4820 48380 4892 48432
rect 4944 48380 4956 48432
rect 4632 48308 4956 48380
rect 10782 48372 10794 49360
rect 10846 48372 10858 49360
rect 14408 49316 14564 49320
rect 14380 49304 14564 49316
rect 14380 49252 14392 49304
rect 14444 49252 14500 49304
rect 14552 49252 14564 49304
rect 14380 49196 14564 49252
rect 14380 49144 14392 49196
rect 14444 49144 14500 49196
rect 14552 49144 14564 49196
rect 14380 49088 14564 49144
rect 14380 49036 14392 49088
rect 14444 49036 14500 49088
rect 14552 49036 14564 49088
rect 14380 48980 14564 49036
rect 14380 48928 14392 48980
rect 14444 48928 14500 48980
rect 14552 48928 14564 48980
rect 14380 48872 14564 48928
rect 14380 48820 14392 48872
rect 14444 48820 14500 48872
rect 14552 48820 14564 48872
rect 14380 48808 14564 48820
rect 14408 48804 14564 48808
rect 10782 48360 10858 48372
rect 14408 48348 14564 48352
rect 4632 48256 4644 48308
rect 4696 48256 4768 48308
rect 4820 48256 4892 48308
rect 4944 48256 4956 48308
rect 4632 48184 4956 48256
rect 4632 48132 4644 48184
rect 4696 48132 4768 48184
rect 4820 48132 4892 48184
rect 4944 48132 4956 48184
rect 4632 48060 4956 48132
rect 4632 48008 4644 48060
rect 4696 48008 4768 48060
rect 4820 48008 4892 48060
rect 4944 48008 4956 48060
rect 4632 47936 4956 48008
rect 14380 48336 14564 48348
rect 14380 48284 14392 48336
rect 14444 48284 14500 48336
rect 14552 48284 14564 48336
rect 14380 48228 14564 48284
rect 14380 48176 14392 48228
rect 14444 48176 14500 48228
rect 14552 48176 14564 48228
rect 14380 48120 14564 48176
rect 14380 48068 14392 48120
rect 14444 48068 14500 48120
rect 14552 48068 14564 48120
rect 14380 48012 14564 48068
rect 14380 47960 14392 48012
rect 14444 47960 14500 48012
rect 14552 47960 14564 48012
rect 4632 47884 4644 47936
rect 4696 47884 4768 47936
rect 4820 47884 4892 47936
rect 4944 47884 4956 47936
rect 4632 47872 4956 47884
rect 11589 47942 11742 47954
rect 3608 47788 3684 47800
rect 3608 46696 3620 47788
rect 3672 46696 3684 47788
rect 11589 47786 11630 47942
rect 11682 47786 11742 47942
rect 14380 47904 14564 47960
rect 14380 47852 14392 47904
rect 14444 47852 14500 47904
rect 14552 47852 14564 47904
rect 14380 47840 14564 47852
rect 14408 47836 14564 47840
rect 11001 47718 11077 47730
rect 11001 47146 11013 47718
rect 11065 47146 11077 47718
rect 11001 47134 11077 47146
rect 3608 46684 3684 46696
rect 3185 46504 3365 46520
rect 3185 46036 3197 46504
rect 3353 46036 3365 46504
rect 11589 46426 11742 47786
rect 12260 46966 12660 46978
rect 12260 46957 12272 46966
rect 12241 46914 12272 46957
rect 12324 46914 12380 46966
rect 12432 46914 12488 46966
rect 12540 46914 12596 46966
rect 12648 46957 12660 46966
rect 12648 46914 13567 46957
rect 12241 46467 13567 46914
rect 3185 46024 3365 46036
rect 14204 45993 14280 46005
rect 14204 45837 14216 45993
rect 14268 45837 14280 45993
rect 14204 45825 14280 45837
rect 3608 44543 3684 44555
rect 3608 43243 3620 44543
rect 3672 43243 3684 44543
rect 12422 44053 12602 44065
rect 12422 44001 12434 44053
rect 12590 44001 12602 44053
rect 12422 43989 12602 44001
rect 3608 43231 3684 43243
rect 10470 43628 11847 43639
rect 10470 43582 10764 43628
rect 10810 43582 10878 43628
rect 10924 43582 10992 43628
rect 11038 43582 11106 43628
rect 11152 43582 11220 43628
rect 11266 43582 11334 43628
rect 11380 43582 11448 43628
rect 11494 43582 11562 43628
rect 11608 43582 11676 43628
rect 11722 43582 11790 43628
rect 11836 43588 11847 43628
rect 11836 43582 14677 43588
rect 10470 43577 14677 43582
rect 10470 43514 12075 43577
rect 10470 43468 10764 43514
rect 10810 43468 10878 43514
rect 10924 43468 10992 43514
rect 11038 43468 11106 43514
rect 11152 43468 11220 43514
rect 11266 43468 11334 43514
rect 11380 43468 11448 43514
rect 11494 43468 11562 43514
rect 11608 43468 11676 43514
rect 11722 43468 11790 43514
rect 11836 43468 12075 43514
rect 10470 43400 12075 43468
rect 10470 43354 10764 43400
rect 10810 43354 10878 43400
rect 10924 43354 10992 43400
rect 11038 43354 11106 43400
rect 11152 43354 11220 43400
rect 11266 43354 11334 43400
rect 11380 43354 11448 43400
rect 11494 43354 11562 43400
rect 11608 43354 11676 43400
rect 11722 43354 11790 43400
rect 11836 43354 12075 43400
rect 10470 43286 12075 43354
rect 10470 43240 10764 43286
rect 10810 43240 10878 43286
rect 10924 43240 10992 43286
rect 11038 43240 11106 43286
rect 11152 43240 11220 43286
rect 11266 43240 11334 43286
rect 11380 43240 11448 43286
rect 11494 43240 11562 43286
rect 11608 43240 11676 43286
rect 11722 43240 11790 43286
rect 11836 43240 12075 43286
rect 10470 43172 12075 43240
rect 10470 43143 10764 43172
rect 10753 43126 10764 43143
rect 10810 43126 10878 43172
rect 10924 43126 10992 43172
rect 11038 43126 11106 43172
rect 11152 43126 11220 43172
rect 11266 43126 11334 43172
rect 11380 43126 11448 43172
rect 11494 43126 11562 43172
rect 11608 43126 11676 43172
rect 11722 43126 11790 43172
rect 11836 43126 12075 43172
rect 10753 43058 12075 43126
rect 10753 43012 10764 43058
rect 10810 43012 10878 43058
rect 10924 43012 10992 43058
rect 11038 43012 11106 43058
rect 11152 43012 11220 43058
rect 11266 43012 11334 43058
rect 11380 43012 11448 43058
rect 11494 43012 11562 43058
rect 11608 43012 11676 43058
rect 11722 43012 11790 43058
rect 11836 43012 12075 43058
rect 3608 42943 3684 42955
rect 3608 41643 3620 42943
rect 3672 41643 3684 42943
rect 10753 42944 12075 43012
rect 10753 42898 10764 42944
rect 10810 42898 10878 42944
rect 10924 42898 10992 42944
rect 11038 42898 11106 42944
rect 11152 42898 11220 42944
rect 11266 42898 11334 42944
rect 11380 42898 11448 42944
rect 11494 42898 11562 42944
rect 11608 42898 11676 42944
rect 11722 42898 11790 42944
rect 11836 42898 12075 42944
rect 10753 42830 12075 42898
rect 10753 42784 10764 42830
rect 10810 42784 10878 42830
rect 10924 42784 10992 42830
rect 11038 42784 11106 42830
rect 11152 42784 11220 42830
rect 11266 42784 11334 42830
rect 11380 42784 11448 42830
rect 11494 42784 11562 42830
rect 11608 42784 11676 42830
rect 11722 42784 11790 42830
rect 11836 42784 12075 42830
rect 10753 42716 12075 42784
rect 10753 42670 10764 42716
rect 10810 42670 10878 42716
rect 10924 42670 10992 42716
rect 11038 42670 11106 42716
rect 11152 42670 11220 42716
rect 11266 42670 11334 42716
rect 11380 42670 11448 42716
rect 11494 42670 11562 42716
rect 11608 42670 11676 42716
rect 11722 42670 11790 42716
rect 11836 42670 12075 42716
rect 10753 42659 12075 42670
rect 3608 41631 3684 41643
rect 11290 41982 11826 41995
rect 11290 41936 11303 41982
rect 11349 41936 11419 41982
rect 11465 41936 11535 41982
rect 11581 41936 11651 41982
rect 11697 41936 11767 41982
rect 11813 41936 11826 41982
rect 11290 41923 11826 41936
rect 11290 41866 11362 41923
rect 11290 41820 11303 41866
rect 11349 41820 11362 41866
rect 11754 41866 11826 41923
rect 11290 41750 11362 41820
rect 11290 41704 11303 41750
rect 11349 41704 11362 41750
rect 11290 41634 11362 41704
rect 11290 41588 11303 41634
rect 11349 41588 11362 41634
rect 11458 41815 11658 41827
rect 11458 41814 11583 41815
rect 11635 41814 11658 41815
rect 11458 41768 11471 41814
rect 11517 41768 11583 41814
rect 11645 41768 11658 41814
rect 11458 41686 11583 41768
rect 11635 41686 11658 41768
rect 11458 41640 11471 41686
rect 11517 41659 11583 41686
rect 11517 41640 11599 41659
rect 11645 41640 11658 41686
rect 11458 41627 11658 41640
rect 11754 41820 11767 41866
rect 11813 41820 11826 41866
rect 11754 41750 11826 41820
rect 11754 41704 11767 41750
rect 11813 41704 11826 41750
rect 11754 41634 11826 41704
rect 11290 41531 11362 41588
rect 11754 41588 11767 41634
rect 11813 41588 11826 41634
rect 11754 41531 11826 41588
rect 11290 41518 11826 41531
rect 11290 41472 11303 41518
rect 11349 41472 11419 41518
rect 11465 41472 11535 41518
rect 11581 41472 11651 41518
rect 11697 41472 11767 41518
rect 11813 41472 11826 41518
rect 11290 41459 11826 41472
rect 11290 41402 11362 41459
rect 11290 41356 11303 41402
rect 11349 41356 11362 41402
rect 11754 41402 11826 41459
rect 11290 41286 11362 41356
rect 11290 41240 11303 41286
rect 11349 41240 11362 41286
rect 11290 41175 11362 41240
rect 11286 41170 11362 41175
rect 11286 41163 11303 41170
rect 11349 41163 11362 41170
rect 11458 41350 11658 41363
rect 11458 41304 11471 41350
rect 11517 41341 11599 41350
rect 11517 41304 11583 41341
rect 11645 41304 11658 41350
rect 11458 41222 11583 41304
rect 11635 41222 11658 41304
rect 11458 41176 11471 41222
rect 11517 41185 11583 41222
rect 11517 41176 11599 41185
rect 11645 41176 11658 41222
rect 11458 41163 11658 41176
rect 11754 41356 11767 41402
rect 11813 41356 11826 41402
rect 11754 41286 11826 41356
rect 11754 41240 11767 41286
rect 11813 41240 11826 41286
rect 11754 41170 11826 41240
rect 1836 41070 3680 41082
rect 1836 41018 1848 41070
rect 3668 41018 3680 41070
rect 1836 41006 3680 41018
rect 11286 41007 11298 41163
rect 11350 41067 11362 41163
rect 11754 41124 11767 41170
rect 11813 41124 11826 41170
rect 11754 41067 11826 41124
rect 12064 41087 12075 42659
rect 12121 43531 12182 43577
rect 14484 43531 14592 43577
rect 12121 43191 14592 43531
rect 12121 43145 12519 43191
rect 13045 43145 13659 43191
rect 14185 43145 14592 43191
rect 12121 43134 14592 43145
rect 12121 42498 12332 43134
rect 12392 43063 13172 43074
rect 12392 43017 12403 43063
rect 12449 43017 13115 43063
rect 13161 43017 13172 43063
rect 12392 42951 13172 43017
rect 12392 42905 12403 42951
rect 12449 42905 13115 42951
rect 13161 42905 13172 42951
rect 12392 42868 13172 42905
rect 12392 42839 13108 42868
rect 13160 42839 13172 42868
rect 12392 42793 12403 42839
rect 12449 42793 13108 42839
rect 13161 42793 13172 42839
rect 12392 42727 13108 42793
rect 13160 42727 13172 42793
rect 12392 42681 12403 42727
rect 12449 42712 13108 42727
rect 12449 42681 13115 42712
rect 13161 42681 13172 42727
rect 12392 42615 13172 42681
rect 12392 42569 12403 42615
rect 12449 42569 13115 42615
rect 13161 42569 13172 42615
rect 12392 42558 13172 42569
rect 13272 42498 13472 43134
rect 13532 43063 14312 43074
rect 13532 43017 13543 43063
rect 13589 43017 14255 43063
rect 14301 43017 14312 43063
rect 13532 42951 14312 43017
rect 13532 42905 13543 42951
rect 13589 42905 14255 42951
rect 14301 42905 14312 42951
rect 13532 42868 14312 42905
rect 13532 42839 13544 42868
rect 13596 42839 14312 42868
rect 13532 42793 13543 42839
rect 13596 42793 14255 42839
rect 14301 42793 14312 42839
rect 13532 42727 13544 42793
rect 13596 42727 14312 42793
rect 13532 42681 13543 42727
rect 13596 42712 14255 42727
rect 13589 42681 14255 42712
rect 14301 42681 14312 42727
rect 13532 42615 14312 42681
rect 13532 42569 13543 42615
rect 13589 42569 14255 42615
rect 14301 42569 14312 42615
rect 13532 42558 14312 42569
rect 12121 42487 13082 42498
rect 12121 42441 12519 42487
rect 13045 42441 13082 42487
rect 12121 42223 13082 42441
rect 12121 42177 12519 42223
rect 13045 42177 13082 42223
rect 12121 42166 13082 42177
rect 13272 42487 14222 42498
rect 13272 42441 13659 42487
rect 14185 42441 14222 42487
rect 13272 42223 14222 42441
rect 13272 42177 13659 42223
rect 14185 42177 14222 42223
rect 13272 42166 14222 42177
rect 12121 41530 12332 42166
rect 12392 42095 13172 42106
rect 12392 42049 12403 42095
rect 12449 42049 13115 42095
rect 13161 42049 13172 42095
rect 12392 41983 13172 42049
rect 12392 41937 12403 41983
rect 12449 41941 13115 41983
rect 12449 41937 13108 41941
rect 13161 41937 13172 41983
rect 12392 41871 13108 41937
rect 13160 41871 13172 41937
rect 12392 41825 12403 41871
rect 12449 41825 13108 41871
rect 13161 41825 13172 41871
rect 12392 41785 13108 41825
rect 13160 41785 13172 41825
rect 12392 41759 13172 41785
rect 12392 41713 12403 41759
rect 12449 41713 13115 41759
rect 13161 41713 13172 41759
rect 12392 41647 13172 41713
rect 12392 41601 12403 41647
rect 12449 41601 13115 41647
rect 13161 41601 13172 41647
rect 12392 41590 13172 41601
rect 13272 41530 13472 42166
rect 13532 42095 14312 42106
rect 13532 42049 13543 42095
rect 13589 42049 14255 42095
rect 14301 42049 14312 42095
rect 13532 41983 14312 42049
rect 13532 41937 13543 41983
rect 13589 41941 14255 41983
rect 13596 41937 14255 41941
rect 14301 41937 14312 41983
rect 13532 41871 13544 41937
rect 13596 41871 14312 41937
rect 13532 41825 13543 41871
rect 13596 41825 14255 41871
rect 14301 41825 14312 41871
rect 13532 41785 13544 41825
rect 13596 41785 14312 41825
rect 13532 41759 14312 41785
rect 13532 41713 13543 41759
rect 13589 41713 14255 41759
rect 14301 41713 14312 41759
rect 13532 41647 14312 41713
rect 13532 41601 13543 41647
rect 13589 41601 14255 41647
rect 14301 41601 14312 41647
rect 13532 41590 14312 41601
rect 12121 41529 13082 41530
rect 13272 41529 14222 41530
rect 14581 41529 14592 43134
rect 12121 41519 14592 41529
rect 12121 41473 12519 41519
rect 13045 41473 13659 41519
rect 14185 41473 14592 41519
rect 12121 41133 14592 41473
rect 12121 41087 12182 41133
rect 14484 41087 14592 41133
rect 14638 43134 14677 43577
rect 14638 41529 14649 43134
rect 14638 41087 14677 41529
rect 12064 41075 14677 41087
rect 11350 41054 11826 41067
rect 11350 41008 11419 41054
rect 11465 41008 11535 41054
rect 11581 41008 11651 41054
rect 11697 41008 11767 41054
rect 11813 41008 11826 41054
rect 11350 41007 11826 41008
rect 11286 40995 11826 41007
rect 11017 40972 11093 40984
rect 11017 40816 11029 40972
rect 11081 40910 11093 40972
rect 11081 40883 11890 40910
rect 11081 40831 11714 40883
rect 11870 40831 11890 40883
rect 11081 40816 11890 40831
rect 11017 40804 11890 40816
rect 14058 40838 14134 40850
rect 14058 40746 14070 40838
rect 1913 40734 14070 40746
rect 1913 40682 1925 40734
rect 2081 40682 4849 40734
rect 5005 40682 7065 40734
rect 7221 40682 10900 40734
rect 11056 40682 14070 40734
rect 14122 40682 14134 40838
rect 1913 40670 14134 40682
rect 11416 40598 13842 40610
rect 1596 40568 5746 40580
rect 1596 40516 1608 40568
rect 1764 40516 5578 40568
rect 5734 40516 5746 40568
rect 11416 40546 11428 40598
rect 11584 40546 13674 40598
rect 13830 40546 13842 40598
rect 11416 40534 13842 40546
rect 1596 40504 5746 40516
rect 10644 40462 13988 40474
rect 10644 40410 10656 40462
rect 10812 40410 11996 40462
rect 12152 40410 13820 40462
rect 13976 40410 13988 40462
rect 10644 40398 13988 40410
rect 184 40306 954 40318
rect 184 40254 202 40306
rect 566 40254 954 40306
rect 184 40250 954 40254
rect 2433 40314 4485 40326
rect 2433 40262 2445 40314
rect 4473 40262 4485 40314
rect 2433 40250 4485 40262
rect 7888 40314 9732 40326
rect 7888 40262 7900 40314
rect 9720 40262 9732 40314
rect 7888 40250 9732 40262
rect 12772 40314 13784 40326
rect 12772 40262 12784 40314
rect 13772 40262 13784 40314
rect 12772 40250 13784 40262
rect 190 40242 578 40250
rect 1771 39788 1847 39800
rect 1771 39216 1783 39788
rect 1835 39216 1847 39788
rect 10327 39788 10403 39800
rect 1771 39204 1847 39216
rect 5083 39758 5159 39770
rect 5083 39186 5095 39758
rect 5147 39186 5159 39758
rect 5083 39174 5159 39186
rect 6049 39758 6125 39770
rect 6049 38770 6061 39758
rect 6113 38770 6125 39758
rect 7015 39758 7091 39770
rect 6306 39057 6382 39459
rect 7015 39186 7027 39758
rect 7079 39186 7091 39758
rect 7015 39174 7091 39186
rect 6306 38877 6504 39057
rect 10327 38800 10339 39788
rect 10391 38800 10403 39788
rect 11200 39788 11276 39800
rect 10644 39046 10720 39058
rect 10644 38890 10656 39046
rect 10708 38890 10720 39046
rect 10644 38878 10720 38890
rect 10888 39046 10964 39058
rect 10888 38890 10900 39046
rect 10952 38890 10964 39046
rect 10888 38878 10964 38890
rect 10327 38788 10403 38800
rect 11200 38800 11212 39788
rect 11264 38800 11276 39788
rect 11200 38788 11276 38800
rect 6049 38758 6125 38770
rect 8293 38688 8369 38700
rect 8293 38532 8305 38688
rect 8357 38532 8369 38688
rect 0 36843 58 38143
rect 110 36843 122 38143
rect 805 38512 881 38524
rect 805 37524 817 38512
rect 869 37524 881 38512
rect 3427 38512 3503 38524
rect 2707 37939 2783 37951
rect 2707 37783 2719 37939
rect 2771 37783 2783 37939
rect 2707 37771 2783 37783
rect 3195 37939 3271 37951
rect 3195 37783 3207 37939
rect 3259 37783 3271 37939
rect 3195 37771 3271 37783
rect 805 37512 881 37524
rect 3427 37524 3439 38512
rect 3491 37524 3503 38512
rect 6049 38512 6125 38524
rect 8293 38520 8369 38532
rect 11520 38685 11596 38697
rect 11520 38529 11532 38685
rect 11584 38529 11596 38685
rect 3659 37939 3735 37951
rect 3659 37783 3671 37939
rect 3723 37783 3735 37939
rect 3659 37771 3735 37783
rect 4147 37939 4223 37951
rect 4147 37783 4159 37939
rect 4211 37783 4223 37939
rect 4147 37771 4223 37783
rect 3427 37512 3503 37524
rect 6049 37524 6061 38512
rect 6113 37524 6125 38512
rect 8671 38512 8747 38524
rect 11520 38517 11596 38529
rect 13303 38675 13379 38687
rect 13303 38519 13315 38675
rect 13367 38519 13379 38675
rect 8439 37939 8515 37951
rect 8439 37783 8451 37939
rect 8503 37783 8515 37939
rect 8439 37771 8515 37783
rect 6049 37512 6125 37524
rect 8671 37524 8683 38512
rect 8735 37524 8747 38512
rect 13303 38507 13379 38519
rect 13439 38023 13515 38035
rect 8895 37939 8971 37951
rect 8895 37783 8907 37939
rect 8959 37783 8971 37939
rect 13439 37867 13451 38023
rect 13503 37867 13515 38023
rect 13439 37855 13515 37867
rect 8895 37771 8971 37783
rect 8671 37512 8747 37524
rect 10331 37568 11551 37580
rect 10331 37516 10343 37568
rect 11539 37516 11551 37568
rect 10331 37504 11551 37516
rect 0 11002 122 36843
rect 8439 37002 8515 37014
rect 8439 36846 8451 37002
rect 8503 36910 8515 37002
rect 8503 36898 13242 36910
rect 8503 36846 13074 36898
rect 13230 36846 13242 36898
rect 8439 36834 13242 36846
rect 8293 36762 13102 36774
rect 8293 36710 8305 36762
rect 8461 36710 12934 36762
rect 13090 36710 13102 36762
rect 8293 36698 13102 36710
rect 2066 36626 2469 36638
rect 2066 36574 2088 36626
rect 2452 36574 2469 36626
rect 2066 36562 2469 36574
rect 4461 36626 9150 36638
rect 4461 36574 4473 36626
rect 4629 36574 5822 36626
rect 5978 36574 8982 36626
rect 9138 36574 9150 36626
rect 4461 36562 9150 36574
rect 1822 36490 3271 36502
rect 1822 36438 1834 36490
rect 1990 36438 3103 36490
rect 3259 36438 3271 36490
rect 1822 36426 3271 36438
rect 3659 36490 9010 36502
rect 3659 36438 3671 36490
rect 3827 36438 6066 36490
rect 6222 36438 8842 36490
rect 8998 36438 9010 36490
rect 3659 36426 9010 36438
rect 2482 36354 12686 36366
rect 2482 36302 2494 36354
rect 2650 36302 5406 36354
rect 5562 36302 9502 36354
rect 9658 36302 12518 36354
rect 12674 36302 12686 36354
rect 2482 36290 12686 36302
rect 1310 36218 13754 36230
rect 1310 36166 1322 36218
rect 1478 36166 6578 36218
rect 6734 36166 8330 36218
rect 8486 36166 13586 36218
rect 13742 36166 13754 36218
rect 1310 36154 13754 36166
rect 3386 36082 13515 36094
rect 3386 36030 3398 36082
rect 3554 36030 4502 36082
rect 4658 36030 10406 36082
rect 10562 36030 11510 36082
rect 11666 36030 13347 36082
rect 13503 36030 13515 36082
rect 3386 36018 13515 36030
rect 486 35946 562 35958
rect 486 34126 498 35946
rect 550 34126 562 35946
rect 724 35946 800 35958
rect 724 34542 736 35946
rect 788 34542 800 35946
rect 724 34530 800 34542
rect 3092 35946 3168 35958
rect 3092 34542 3104 35946
rect 3156 34542 3168 35946
rect 3092 34530 3168 34542
rect 3990 35946 4066 35958
rect 1822 34435 1898 34447
rect 1822 34279 1834 34435
rect 1886 34279 1898 34435
rect 1822 34267 1898 34279
rect 2066 34435 2142 34447
rect 2066 34279 2078 34435
rect 2130 34279 2142 34435
rect 2066 34267 2142 34279
rect 2482 34435 2558 34447
rect 2482 34279 2494 34435
rect 2546 34279 2558 34435
rect 2482 34267 2558 34279
rect 486 34114 562 34126
rect 486 33851 562 33863
rect 486 30055 498 33851
rect 550 30055 562 33851
rect 3990 33294 4002 35946
rect 4054 33294 4066 35946
rect 4888 35946 4964 35958
rect 4888 34542 4900 35946
rect 4952 34542 4964 35946
rect 8567 35946 8747 35958
rect 8567 35894 8579 35946
rect 8735 35894 8747 35946
rect 8567 35882 8747 35894
rect 10100 35946 10176 35958
rect 4888 34530 4964 34542
rect 10100 34542 10112 35946
rect 10164 34542 10176 35946
rect 10100 34530 10176 34542
rect 10998 35946 11074 35958
rect 5498 34435 5574 34447
rect 5498 34279 5510 34435
rect 5562 34279 5574 34435
rect 5498 34267 5574 34279
rect 5914 34435 5990 34447
rect 5914 34279 5926 34435
rect 5978 34279 5990 34435
rect 5914 34267 5990 34279
rect 6158 34435 6234 34447
rect 6158 34279 6170 34435
rect 6222 34279 6234 34435
rect 6158 34267 6234 34279
rect 8830 34435 8906 34447
rect 8830 34279 8842 34435
rect 8894 34279 8906 34435
rect 8830 34267 8906 34279
rect 9074 34435 9150 34447
rect 9074 34279 9086 34435
rect 9138 34279 9150 34435
rect 9074 34267 9150 34279
rect 9490 34435 9566 34447
rect 9490 34279 9502 34435
rect 9554 34279 9566 34435
rect 9490 34267 9566 34279
rect 3990 33282 4066 33294
rect 10998 33294 11010 35946
rect 11062 33294 11074 35946
rect 11896 35946 11972 35958
rect 11896 34542 11908 35946
rect 11960 34542 11972 35946
rect 13919 35890 14119 38520
rect 14942 38143 15064 51295
rect 14942 36843 14954 38143
rect 15006 36843 15064 38143
rect 11896 34530 11972 34542
rect 12506 34435 12582 34447
rect 12506 34279 12518 34435
rect 12570 34279 12582 34435
rect 12506 34267 12582 34279
rect 12922 34435 12998 34447
rect 12922 34279 12934 34435
rect 12986 34279 12998 34435
rect 12922 34267 12998 34279
rect 13166 34435 13242 34447
rect 13166 34279 13178 34435
rect 13230 34279 13242 34435
rect 13166 34267 13242 34279
rect 10998 33282 11074 33294
rect 14502 33851 14578 33863
rect 3990 32825 4066 32837
rect 968 32690 1044 32702
rect 968 30454 980 32690
rect 1032 30454 1044 32690
rect 2360 32690 2436 32702
rect 968 30442 1044 30454
rect 1456 30678 1532 30690
rect 1456 30314 1468 30678
rect 1520 30314 1532 30678
rect 1456 30302 1532 30314
rect 1700 30678 1776 30690
rect 1700 30314 1712 30678
rect 1764 30314 1776 30678
rect 2360 30454 2372 32690
rect 2424 30454 2436 32690
rect 2360 30442 2436 30454
rect 2776 32690 2852 32702
rect 2776 30454 2788 32690
rect 2840 30454 2852 32690
rect 3264 32690 3340 32702
rect 3264 31078 3276 32690
rect 3328 31078 3340 32690
rect 3264 31066 3340 31078
rect 3752 32640 3828 32652
rect 3752 31028 3764 32640
rect 3816 31028 3828 32640
rect 3752 31016 3828 31028
rect 3990 31005 4002 32825
rect 4054 31005 4066 32825
rect 10998 32825 11074 32837
rect 4716 32690 4792 32702
rect 4228 32640 4304 32652
rect 4228 31028 4240 32640
rect 4292 31028 4304 32640
rect 4716 31078 4728 32690
rect 4780 31078 4792 32690
rect 4716 31066 4792 31078
rect 5204 32690 5280 32702
rect 5204 31078 5216 32690
rect 5268 31078 5280 32690
rect 5204 31066 5280 31078
rect 5620 32690 5696 32702
rect 5620 31078 5632 32690
rect 5684 31078 5696 32690
rect 5620 31066 5696 31078
rect 7012 32690 7088 32702
rect 4228 31016 4304 31028
rect 3990 30993 4066 31005
rect 3020 30858 3096 30870
rect 3020 30494 3032 30858
rect 3084 30494 3096 30858
rect 4472 30858 4548 30870
rect 3020 30482 3096 30494
rect 3508 30678 3584 30690
rect 2776 30442 2852 30454
rect 1700 30302 1776 30314
rect 3508 30314 3520 30678
rect 3572 30314 3584 30678
rect 4472 30494 4484 30858
rect 4536 30494 4548 30858
rect 4472 30482 4548 30494
rect 4960 30678 5036 30690
rect 3508 30302 3584 30314
rect 4960 30314 4972 30678
rect 5024 30314 5036 30678
rect 4960 30302 5036 30314
rect 6524 30678 6600 30690
rect 6524 30314 6536 30678
rect 6588 30314 6600 30678
rect 6524 30302 6600 30314
rect 6768 30678 6844 30690
rect 6768 30314 6780 30678
rect 6832 30314 6844 30678
rect 7012 30454 7024 32690
rect 7076 30454 7088 32690
rect 7012 30442 7088 30454
rect 7976 32690 8052 32702
rect 7976 30454 7988 32690
rect 8040 30454 8052 32690
rect 9368 32690 9444 32702
rect 9368 31078 9380 32690
rect 9432 31078 9444 32690
rect 9368 31066 9444 31078
rect 9784 32690 9860 32702
rect 9784 31078 9796 32690
rect 9848 31078 9860 32690
rect 9784 31066 9860 31078
rect 10272 32690 10348 32702
rect 10272 31078 10284 32690
rect 10336 31078 10348 32690
rect 10272 31066 10348 31078
rect 10760 32640 10836 32652
rect 10760 31028 10772 32640
rect 10824 31028 10836 32640
rect 10760 31016 10836 31028
rect 10998 31005 11010 32825
rect 11062 31005 11074 32825
rect 11724 32690 11800 32702
rect 11236 32640 11312 32652
rect 11236 31028 11248 32640
rect 11300 31028 11312 32640
rect 11724 31078 11736 32690
rect 11788 31078 11800 32690
rect 11724 31066 11800 31078
rect 12212 32690 12288 32702
rect 11236 31016 11312 31028
rect 10998 30993 11074 31005
rect 10516 30858 10592 30870
rect 7976 30442 8052 30454
rect 8464 30678 8540 30690
rect 6768 30302 6844 30314
rect 8464 30314 8476 30678
rect 8528 30314 8540 30678
rect 8464 30302 8540 30314
rect 8708 30678 8784 30690
rect 8708 30314 8720 30678
rect 8772 30314 8784 30678
rect 8708 30302 8784 30314
rect 10028 30678 10104 30690
rect 10028 30314 10040 30678
rect 10092 30314 10104 30678
rect 10516 30494 10528 30858
rect 10580 30494 10592 30858
rect 11968 30858 12044 30870
rect 10516 30482 10592 30494
rect 11480 30678 11556 30690
rect 10028 30302 10104 30314
rect 11480 30314 11492 30678
rect 11544 30314 11556 30678
rect 11968 30494 11980 30858
rect 12032 30494 12044 30858
rect 11968 30482 12044 30494
rect 12212 30454 12224 32690
rect 12276 30454 12288 32690
rect 12212 30442 12288 30454
rect 12628 32690 12704 32702
rect 12628 30454 12640 32690
rect 12692 30454 12704 32690
rect 14020 32690 14096 32702
rect 12628 30442 12704 30454
rect 13532 30678 13608 30690
rect 11480 30302 11556 30314
rect 13532 30314 13544 30678
rect 13596 30314 13608 30678
rect 13532 30302 13608 30314
rect 13776 30678 13852 30690
rect 13776 30314 13788 30678
rect 13840 30314 13852 30678
rect 14020 30454 14032 32690
rect 14084 30454 14096 32690
rect 14020 30442 14096 30454
rect 13776 30302 13852 30314
rect 486 30043 562 30055
rect 2000 30107 3324 30119
rect 2000 30055 2012 30107
rect 3312 30055 3324 30107
rect 2000 30043 3324 30055
rect 11937 30107 13261 30119
rect 11937 30055 11949 30107
rect 13249 30055 13261 30107
rect 11937 30043 13261 30055
rect 14502 30055 14514 33851
rect 14566 30055 14578 33851
rect 14502 30043 14578 30055
rect 1367 29817 6612 29841
rect 1367 29765 1379 29817
rect 1535 29765 6444 29817
rect 6600 29765 6612 29817
rect 1367 29741 6612 29765
rect 8696 29817 13699 29841
rect 8696 29765 8708 29817
rect 8864 29765 13531 29817
rect 13687 29765 13699 29817
rect 8696 29741 13699 29765
rect 1547 29637 6856 29661
rect 1547 29585 1559 29637
rect 1715 29585 6688 29637
rect 6844 29585 6856 29637
rect 1547 29561 6856 29585
rect 8452 29637 13519 29661
rect 8452 29585 8464 29637
rect 8620 29585 13351 29637
rect 13507 29585 13519 29637
rect 8452 29561 13519 29585
rect 2340 29430 3888 29481
rect 2340 29378 3508 29430
rect 3664 29378 3888 29430
rect 2340 29319 3888 29378
rect 2340 24880 2502 29319
rect 3726 24880 3888 29319
rect 4112 29469 4274 29481
rect 4112 29313 4167 29469
rect 4219 29313 4274 29469
rect 4112 24880 4274 29313
rect 4960 29469 5648 29481
rect 4960 29313 4972 29469
rect 5024 29319 5648 29469
rect 5024 29313 5036 29319
rect 4960 29301 5036 29313
rect 5486 24880 5648 29319
rect 5877 29469 7420 29481
rect 5877 29313 5926 29469
rect 5978 29319 7420 29469
rect 5978 29313 6039 29319
rect 5877 24880 6039 29313
rect 7258 24880 7420 29319
rect 7646 29469 9190 29481
rect 7646 29319 9088 29469
rect 7646 24880 7808 29319
rect 9028 29313 9088 29319
rect 9140 29313 9190 29469
rect 9028 24880 9190 29313
rect 9415 29469 10106 29481
rect 9415 29319 10042 29469
rect 9415 24880 9577 29319
rect 10030 29313 10042 29319
rect 10094 29313 10106 29469
rect 10030 29301 10106 29313
rect 10794 29469 10956 29481
rect 10794 29313 10847 29469
rect 10899 29313 10956 29469
rect 10794 24880 10956 29313
rect 11181 29430 12729 29481
rect 11181 29378 11402 29430
rect 11558 29378 12729 29430
rect 11181 29319 12729 29378
rect 11181 24880 11343 29319
rect 12567 24880 12729 29319
rect 14942 11002 15064 36843
rect 0 10991 268 11002
rect 0 1357 211 10991
rect 257 1357 268 10991
rect 0 1217 268 1357
rect 14734 10991 15064 11002
rect 14734 1357 14745 10991
rect 14791 1357 15064 10991
rect 14734 1217 15064 1357
rect 0 1206 15064 1217
rect 0 1160 287 1206
rect 333 1160 411 1206
rect 457 1160 535 1206
rect 581 1160 659 1206
rect 705 1160 783 1206
rect 829 1160 907 1206
rect 953 1160 1031 1206
rect 1077 1160 1155 1206
rect 1201 1160 1279 1206
rect 1325 1160 1403 1206
rect 1449 1160 1527 1206
rect 1573 1160 1651 1206
rect 1697 1160 1775 1206
rect 1821 1160 1899 1206
rect 1945 1160 2023 1206
rect 2069 1160 2147 1206
rect 2193 1160 2271 1206
rect 2317 1160 2395 1206
rect 2441 1160 2519 1206
rect 2565 1160 2643 1206
rect 2689 1160 2767 1206
rect 2813 1160 2891 1206
rect 2937 1160 3015 1206
rect 3061 1160 3139 1206
rect 3185 1160 3263 1206
rect 3309 1160 3387 1206
rect 3433 1160 3511 1206
rect 3557 1160 3635 1206
rect 3681 1160 3759 1206
rect 3805 1160 3883 1206
rect 3929 1160 4007 1206
rect 4053 1160 4131 1206
rect 4177 1160 4255 1206
rect 4301 1160 4379 1206
rect 4425 1160 4503 1206
rect 4549 1160 4627 1206
rect 4673 1160 4751 1206
rect 4797 1160 4875 1206
rect 4921 1160 4999 1206
rect 5045 1160 5123 1206
rect 5169 1160 5247 1206
rect 5293 1160 5371 1206
rect 5417 1160 5495 1206
rect 5541 1160 5619 1206
rect 5665 1160 5743 1206
rect 5789 1160 5867 1206
rect 5913 1160 5991 1206
rect 6037 1160 6115 1206
rect 6161 1160 6239 1206
rect 6285 1160 6363 1206
rect 6409 1160 6487 1206
rect 6533 1160 6611 1206
rect 6657 1160 6735 1206
rect 6781 1160 6859 1206
rect 6905 1160 6983 1206
rect 7029 1160 7107 1206
rect 7153 1160 7231 1206
rect 7277 1160 7355 1206
rect 7401 1160 7479 1206
rect 7525 1160 7603 1206
rect 7649 1160 7727 1206
rect 7773 1160 7851 1206
rect 7897 1160 7975 1206
rect 8021 1160 8099 1206
rect 8145 1160 8223 1206
rect 8269 1160 8347 1206
rect 8393 1160 8471 1206
rect 8517 1160 8595 1206
rect 8641 1160 8719 1206
rect 8765 1160 8843 1206
rect 8889 1160 8967 1206
rect 9013 1160 9091 1206
rect 9137 1160 9215 1206
rect 9261 1160 9339 1206
rect 9385 1160 9463 1206
rect 9509 1160 9587 1206
rect 9633 1160 9711 1206
rect 9757 1160 9835 1206
rect 9881 1160 9959 1206
rect 10005 1160 10083 1206
rect 10129 1160 10207 1206
rect 10253 1160 10331 1206
rect 10377 1160 10455 1206
rect 10501 1160 10579 1206
rect 10625 1160 10703 1206
rect 10749 1160 10827 1206
rect 10873 1160 10951 1206
rect 10997 1160 11075 1206
rect 11121 1160 11199 1206
rect 11245 1160 11323 1206
rect 11369 1160 11447 1206
rect 11493 1160 11571 1206
rect 11617 1160 11695 1206
rect 11741 1160 11819 1206
rect 11865 1160 11943 1206
rect 11989 1160 12067 1206
rect 12113 1160 12191 1206
rect 12237 1160 12315 1206
rect 12361 1160 12439 1206
rect 12485 1160 12563 1206
rect 12609 1160 12687 1206
rect 12733 1160 12811 1206
rect 12857 1160 12935 1206
rect 12981 1160 13059 1206
rect 13105 1160 13183 1206
rect 13229 1160 13307 1206
rect 13353 1160 13431 1206
rect 13477 1160 13555 1206
rect 13601 1160 13679 1206
rect 13725 1160 13803 1206
rect 13849 1160 13927 1206
rect 13973 1160 14051 1206
rect 14097 1160 14175 1206
rect 14221 1160 14299 1206
rect 14345 1160 14423 1206
rect 14469 1160 14547 1206
rect 14593 1160 14671 1206
rect 14717 1160 15064 1206
rect 0 1082 15064 1160
rect 0 1036 287 1082
rect 333 1036 411 1082
rect 457 1036 535 1082
rect 581 1036 659 1082
rect 705 1036 783 1082
rect 829 1036 907 1082
rect 953 1036 1031 1082
rect 1077 1036 1155 1082
rect 1201 1036 1279 1082
rect 1325 1036 1403 1082
rect 1449 1036 1527 1082
rect 1573 1036 1651 1082
rect 1697 1036 1775 1082
rect 1821 1036 1899 1082
rect 1945 1036 2023 1082
rect 2069 1036 2147 1082
rect 2193 1036 2271 1082
rect 2317 1036 2395 1082
rect 2441 1036 2519 1082
rect 2565 1036 2643 1082
rect 2689 1036 2767 1082
rect 2813 1036 2891 1082
rect 2937 1036 3015 1082
rect 3061 1036 3139 1082
rect 3185 1036 3263 1082
rect 3309 1036 3387 1082
rect 3433 1036 3511 1082
rect 3557 1036 3635 1082
rect 3681 1036 3759 1082
rect 3805 1036 3883 1082
rect 3929 1036 4007 1082
rect 4053 1036 4131 1082
rect 4177 1036 4255 1082
rect 4301 1036 4379 1082
rect 4425 1036 4503 1082
rect 4549 1036 4627 1082
rect 4673 1036 4751 1082
rect 4797 1036 4875 1082
rect 4921 1036 4999 1082
rect 5045 1036 5123 1082
rect 5169 1036 5247 1082
rect 5293 1036 5371 1082
rect 5417 1036 5495 1082
rect 5541 1036 5619 1082
rect 5665 1036 5743 1082
rect 5789 1036 5867 1082
rect 5913 1036 5991 1082
rect 6037 1036 6115 1082
rect 6161 1036 6239 1082
rect 6285 1036 6363 1082
rect 6409 1036 6487 1082
rect 6533 1036 6611 1082
rect 6657 1036 6735 1082
rect 6781 1036 6859 1082
rect 6905 1036 6983 1082
rect 7029 1036 7107 1082
rect 7153 1036 7231 1082
rect 7277 1036 7355 1082
rect 7401 1036 7479 1082
rect 7525 1036 7603 1082
rect 7649 1036 7727 1082
rect 7773 1036 7851 1082
rect 7897 1036 7975 1082
rect 8021 1036 8099 1082
rect 8145 1036 8223 1082
rect 8269 1036 8347 1082
rect 8393 1036 8471 1082
rect 8517 1036 8595 1082
rect 8641 1036 8719 1082
rect 8765 1036 8843 1082
rect 8889 1036 8967 1082
rect 9013 1036 9091 1082
rect 9137 1036 9215 1082
rect 9261 1036 9339 1082
rect 9385 1036 9463 1082
rect 9509 1036 9587 1082
rect 9633 1036 9711 1082
rect 9757 1036 9835 1082
rect 9881 1036 9959 1082
rect 10005 1036 10083 1082
rect 10129 1036 10207 1082
rect 10253 1036 10331 1082
rect 10377 1036 10455 1082
rect 10501 1036 10579 1082
rect 10625 1036 10703 1082
rect 10749 1036 10827 1082
rect 10873 1036 10951 1082
rect 10997 1036 11075 1082
rect 11121 1036 11199 1082
rect 11245 1036 11323 1082
rect 11369 1036 11447 1082
rect 11493 1036 11571 1082
rect 11617 1036 11695 1082
rect 11741 1036 11819 1082
rect 11865 1036 11943 1082
rect 11989 1036 12067 1082
rect 12113 1036 12191 1082
rect 12237 1036 12315 1082
rect 12361 1036 12439 1082
rect 12485 1036 12563 1082
rect 12609 1036 12687 1082
rect 12733 1036 12811 1082
rect 12857 1036 12935 1082
rect 12981 1036 13059 1082
rect 13105 1036 13183 1082
rect 13229 1036 13307 1082
rect 13353 1036 13431 1082
rect 13477 1036 13555 1082
rect 13601 1036 13679 1082
rect 13725 1036 13803 1082
rect 13849 1036 13927 1082
rect 13973 1036 14051 1082
rect 14097 1036 14175 1082
rect 14221 1036 14299 1082
rect 14345 1036 14423 1082
rect 14469 1036 14547 1082
rect 14593 1036 14671 1082
rect 14717 1036 15064 1082
rect 0 846 15064 1036
rect 0 708 122 846
rect 14942 708 15064 846
<< via1 >>
rect 716 57171 768 57327
rect 1486 57275 1642 57327
rect 13822 57275 14082 57327
rect 2522 57156 2574 57160
rect 2646 57156 2698 57160
rect 2770 57156 2822 57160
rect 2894 57156 2946 57160
rect 3018 57156 3070 57160
rect 3142 57156 3194 57160
rect 3266 57156 3318 57160
rect 3390 57156 3442 57160
rect 3514 57156 3566 57160
rect 3638 57156 3690 57160
rect 3762 57156 3814 57160
rect 3886 57156 3938 57160
rect 4010 57156 4062 57160
rect 4134 57156 4186 57160
rect 4258 57156 4310 57160
rect 4382 57156 4434 57160
rect 4506 57156 4558 57160
rect 4630 57156 4682 57160
rect 4754 57156 4806 57160
rect 4878 57156 4930 57160
rect 5002 57156 5054 57160
rect 5126 57156 5178 57160
rect 5250 57156 5302 57160
rect 5374 57156 5426 57160
rect 5498 57156 5550 57160
rect 5622 57156 5674 57160
rect 5746 57156 5798 57160
rect 5870 57156 5922 57160
rect 5994 57156 6046 57160
rect 6118 57156 6170 57160
rect 6242 57156 6294 57160
rect 6366 57156 6418 57160
rect 6490 57156 6542 57160
rect 6614 57156 6666 57160
rect 6738 57156 6790 57160
rect 6862 57156 6914 57160
rect 6986 57156 7038 57160
rect 7110 57156 7162 57160
rect 7234 57156 7286 57160
rect 7358 57156 7410 57160
rect 7482 57156 7534 57160
rect 7606 57156 7658 57160
rect 7730 57156 7782 57160
rect 7854 57156 7906 57160
rect 7978 57156 8030 57160
rect 8102 57156 8154 57160
rect 8226 57156 8278 57160
rect 8350 57156 8402 57160
rect 8474 57156 8526 57160
rect 8598 57156 8650 57160
rect 8722 57156 8774 57160
rect 8846 57156 8898 57160
rect 8970 57156 9022 57160
rect 9094 57156 9146 57160
rect 9218 57156 9270 57160
rect 9342 57156 9394 57160
rect 9466 57156 9518 57160
rect 9590 57156 9642 57160
rect 9714 57156 9766 57160
rect 9838 57156 9890 57160
rect 9962 57156 10014 57160
rect 10086 57156 10138 57160
rect 10210 57156 10262 57160
rect 10334 57156 10386 57160
rect 10458 57156 10510 57160
rect 10582 57156 10634 57160
rect 10706 57156 10758 57160
rect 10830 57156 10882 57160
rect 10954 57156 11006 57160
rect 11078 57156 11130 57160
rect 11202 57156 11254 57160
rect 11326 57156 11378 57160
rect 11450 57156 11502 57160
rect 11574 57156 11626 57160
rect 11698 57156 11750 57160
rect 11822 57156 11874 57160
rect 11946 57156 11998 57160
rect 12070 57156 12122 57160
rect 12194 57156 12246 57160
rect 12318 57156 12370 57160
rect 12442 57156 12494 57160
rect 12566 57156 12618 57160
rect 12690 57156 12742 57160
rect 12814 57156 12866 57160
rect 12938 57156 12990 57160
rect 13062 57156 13114 57160
rect 13186 57156 13238 57160
rect 13310 57156 13362 57160
rect 13434 57156 13486 57160
rect 13558 57156 13610 57160
rect 2522 57108 2574 57156
rect 2646 57108 2698 57156
rect 2770 57108 2822 57156
rect 2894 57108 2946 57156
rect 3018 57108 3070 57156
rect 3142 57108 3194 57156
rect 3266 57108 3318 57156
rect 3390 57108 3442 57156
rect 3514 57108 3566 57156
rect 3638 57108 3690 57156
rect 3762 57108 3814 57156
rect 3886 57108 3938 57156
rect 4010 57108 4062 57156
rect 4134 57108 4186 57156
rect 4258 57108 4310 57156
rect 4382 57108 4434 57156
rect 4506 57108 4558 57156
rect 4630 57108 4682 57156
rect 4754 57108 4806 57156
rect 4878 57108 4930 57156
rect 5002 57108 5054 57156
rect 5126 57108 5178 57156
rect 5250 57108 5302 57156
rect 5374 57108 5426 57156
rect 5498 57108 5550 57156
rect 5622 57108 5674 57156
rect 5746 57108 5798 57156
rect 5870 57108 5922 57156
rect 5994 57108 6046 57156
rect 6118 57108 6170 57156
rect 6242 57108 6294 57156
rect 6366 57108 6418 57156
rect 6490 57108 6542 57156
rect 6614 57108 6666 57156
rect 6738 57108 6790 57156
rect 6862 57108 6914 57156
rect 6986 57108 7038 57156
rect 7110 57108 7162 57156
rect 7234 57108 7286 57156
rect 7358 57108 7410 57156
rect 7482 57108 7534 57156
rect 7606 57108 7658 57156
rect 7730 57108 7782 57156
rect 7854 57108 7906 57156
rect 7978 57108 8030 57156
rect 8102 57108 8154 57156
rect 8226 57108 8278 57156
rect 8350 57108 8402 57156
rect 8474 57108 8526 57156
rect 8598 57108 8650 57156
rect 8722 57108 8774 57156
rect 8846 57108 8898 57156
rect 8970 57108 9022 57156
rect 9094 57108 9146 57156
rect 9218 57108 9270 57156
rect 9342 57108 9394 57156
rect 9466 57108 9518 57156
rect 9590 57108 9642 57156
rect 9714 57108 9766 57156
rect 9838 57108 9890 57156
rect 9962 57108 10014 57156
rect 10086 57108 10138 57156
rect 10210 57108 10262 57156
rect 10334 57108 10386 57156
rect 10458 57108 10510 57156
rect 10582 57108 10634 57156
rect 10706 57108 10758 57156
rect 10830 57108 10882 57156
rect 10954 57108 11006 57156
rect 11078 57108 11130 57156
rect 11202 57108 11254 57156
rect 11326 57108 11378 57156
rect 11450 57108 11502 57156
rect 11574 57108 11626 57156
rect 11698 57108 11750 57156
rect 11822 57108 11874 57156
rect 11946 57108 11998 57156
rect 12070 57108 12122 57156
rect 12194 57108 12246 57156
rect 12318 57108 12370 57156
rect 12442 57108 12494 57156
rect 12566 57108 12618 57156
rect 12690 57108 12742 57156
rect 12814 57108 12866 57156
rect 12938 57108 12990 57156
rect 13062 57108 13114 57156
rect 13186 57108 13238 57156
rect 13310 57108 13362 57156
rect 13434 57108 13486 57156
rect 13558 57108 13610 57156
rect 2522 56984 2574 57036
rect 2646 56984 2698 57036
rect 2770 56984 2822 57036
rect 2894 56984 2946 57036
rect 3018 56984 3070 57036
rect 3142 56984 3194 57036
rect 3266 56984 3318 57036
rect 3390 56984 3442 57036
rect 3514 56984 3566 57036
rect 3638 56984 3690 57036
rect 3762 56984 3814 57036
rect 3886 56984 3938 57036
rect 4010 56984 4062 57036
rect 4134 56984 4186 57036
rect 4258 56984 4310 57036
rect 4382 56984 4434 57036
rect 4506 56984 4558 57036
rect 4630 56984 4682 57036
rect 4754 56984 4806 57036
rect 4878 56984 4930 57036
rect 5002 56984 5054 57036
rect 5126 56984 5178 57036
rect 5250 56984 5302 57036
rect 5374 56984 5426 57036
rect 5498 56984 5550 57036
rect 5622 56984 5674 57036
rect 5746 56984 5798 57036
rect 5870 56984 5922 57036
rect 5994 56984 6046 57036
rect 6118 56984 6170 57036
rect 6242 56984 6294 57036
rect 6366 56984 6418 57036
rect 6490 56984 6542 57036
rect 6614 56984 6666 57036
rect 6738 56984 6790 57036
rect 6862 56984 6914 57036
rect 6986 56984 7038 57036
rect 7110 56984 7162 57036
rect 7234 56984 7286 57036
rect 7358 56984 7410 57036
rect 7482 56984 7534 57036
rect 7606 56984 7658 57036
rect 7730 56984 7782 57036
rect 7854 56984 7906 57036
rect 7978 56984 8030 57036
rect 8102 56984 8154 57036
rect 8226 56984 8278 57036
rect 8350 56984 8402 57036
rect 8474 56984 8526 57036
rect 8598 56984 8650 57036
rect 8722 56984 8774 57036
rect 8846 56984 8898 57036
rect 8970 56984 9022 57036
rect 9094 56984 9146 57036
rect 9218 56984 9270 57036
rect 9342 56984 9394 57036
rect 9466 56984 9518 57036
rect 9590 56984 9642 57036
rect 9714 56984 9766 57036
rect 9838 56984 9890 57036
rect 9962 56984 10014 57036
rect 10086 56984 10138 57036
rect 10210 56984 10262 57036
rect 10334 56984 10386 57036
rect 10458 56984 10510 57036
rect 10582 56984 10634 57036
rect 10706 56984 10758 57036
rect 10830 56984 10882 57036
rect 10954 56984 11006 57036
rect 11078 56984 11130 57036
rect 11202 56984 11254 57036
rect 11326 56984 11378 57036
rect 11450 56984 11502 57036
rect 11574 56984 11626 57036
rect 11698 56984 11750 57036
rect 11822 56984 11874 57036
rect 11946 56984 11998 57036
rect 12070 56984 12122 57036
rect 12194 56984 12246 57036
rect 12318 56984 12370 57036
rect 12442 56984 12494 57036
rect 12566 56984 12618 57036
rect 12690 56984 12742 57036
rect 12814 56984 12866 57036
rect 12938 56984 12990 57036
rect 13062 56984 13114 57036
rect 13186 56984 13238 57036
rect 13310 56984 13362 57036
rect 13434 56984 13486 57036
rect 13558 56984 13610 57036
rect 2522 56860 2574 56912
rect 2646 56860 2698 56912
rect 2770 56864 2822 56912
rect 2894 56864 2946 56912
rect 3018 56864 3070 56912
rect 3142 56864 3194 56912
rect 3266 56864 3318 56912
rect 3390 56864 3442 56912
rect 3514 56864 3566 56912
rect 3638 56864 3690 56912
rect 2770 56860 2797 56864
rect 2797 56860 2822 56864
rect 2894 56860 2946 56864
rect 3018 56860 3070 56864
rect 3142 56860 3194 56864
rect 3266 56860 3318 56864
rect 3390 56860 3442 56864
rect 3514 56860 3566 56864
rect 3638 56860 3690 56864
rect 3762 56860 3814 56912
rect 3886 56860 3938 56912
rect 4010 56860 4062 56912
rect 4134 56860 4186 56912
rect 4258 56864 4310 56912
rect 4382 56864 4434 56912
rect 4506 56864 4558 56912
rect 4630 56864 4682 56912
rect 4754 56864 4806 56912
rect 4878 56864 4930 56912
rect 5002 56864 5054 56912
rect 5126 56864 5178 56912
rect 4258 56860 4297 56864
rect 4297 56860 4310 56864
rect 4382 56860 4434 56864
rect 4506 56860 4558 56864
rect 4630 56860 4682 56864
rect 4754 56860 4806 56864
rect 4878 56860 4930 56864
rect 5002 56860 5054 56864
rect 5126 56860 5178 56864
rect 5250 56860 5302 56912
rect 5374 56860 5426 56912
rect 5498 56860 5550 56912
rect 5622 56860 5674 56912
rect 5746 56864 5798 56912
rect 5870 56864 5922 56912
rect 5994 56864 6046 56912
rect 6118 56864 6170 56912
rect 6242 56864 6294 56912
rect 6366 56864 6418 56912
rect 6490 56864 6542 56912
rect 6614 56864 6666 56912
rect 5746 56860 5797 56864
rect 5797 56860 5798 56864
rect 5870 56860 5922 56864
rect 5994 56860 6046 56864
rect 6118 56860 6170 56864
rect 6242 56860 6294 56864
rect 6366 56860 6418 56864
rect 6490 56860 6542 56864
rect 6614 56860 6666 56864
rect 6738 56860 6790 56912
rect 6862 56860 6914 56912
rect 6986 56860 7038 56912
rect 7110 56860 7162 56912
rect 7234 56860 7286 56912
rect 7358 56864 7410 56912
rect 7482 56864 7534 56912
rect 7606 56864 7658 56912
rect 7730 56864 7782 56912
rect 7854 56864 7906 56912
rect 7978 56864 8030 56912
rect 8102 56864 8154 56912
rect 7358 56860 7410 56864
rect 7482 56860 7534 56864
rect 7606 56860 7658 56864
rect 7730 56860 7782 56864
rect 7854 56860 7906 56864
rect 7978 56860 8030 56864
rect 8102 56860 8154 56864
rect 8226 56860 8278 56912
rect 8350 56860 8402 56912
rect 8474 56860 8526 56912
rect 8598 56860 8650 56912
rect 8722 56860 8774 56912
rect 8846 56864 8898 56912
rect 8970 56864 9022 56912
rect 9094 56864 9146 56912
rect 9218 56864 9270 56912
rect 9342 56864 9394 56912
rect 9466 56864 9518 56912
rect 9590 56864 9642 56912
rect 9714 56864 9766 56912
rect 8846 56860 8898 56864
rect 8970 56860 9022 56864
rect 9094 56860 9146 56864
rect 9218 56860 9270 56864
rect 9342 56860 9394 56864
rect 9466 56860 9518 56864
rect 9590 56860 9642 56864
rect 9714 56860 9723 56864
rect 9723 56860 9766 56864
rect 9838 56860 9890 56912
rect 9962 56860 10014 56912
rect 10086 56860 10138 56912
rect 10210 56860 10262 56912
rect 10334 56864 10386 56912
rect 10458 56864 10510 56912
rect 10582 56864 10634 56912
rect 10706 56864 10758 56912
rect 10830 56864 10882 56912
rect 10954 56864 11006 56912
rect 11078 56864 11130 56912
rect 11202 56864 11254 56912
rect 10334 56860 10386 56864
rect 10458 56860 10510 56864
rect 10582 56860 10634 56864
rect 10706 56860 10758 56864
rect 10830 56860 10882 56864
rect 10954 56860 11006 56864
rect 11078 56860 11130 56864
rect 11202 56860 11223 56864
rect 11223 56860 11254 56864
rect 11326 56860 11378 56912
rect 11450 56860 11502 56912
rect 11574 56860 11626 56912
rect 11698 56860 11750 56912
rect 11822 56864 11874 56912
rect 11946 56864 11998 56912
rect 12070 56864 12122 56912
rect 12194 56864 12246 56912
rect 12318 56864 12370 56912
rect 12442 56864 12494 56912
rect 12566 56864 12618 56912
rect 12690 56864 12742 56912
rect 11822 56860 11874 56864
rect 11946 56860 11998 56864
rect 12070 56860 12122 56864
rect 12194 56860 12246 56864
rect 12318 56860 12370 56864
rect 12442 56860 12494 56864
rect 12566 56860 12618 56864
rect 12690 56860 12723 56864
rect 12723 56860 12742 56864
rect 12814 56860 12866 56912
rect 12938 56860 12990 56912
rect 13062 56860 13114 56912
rect 13186 56860 13238 56912
rect 13310 56864 13362 56912
rect 13434 56864 13486 56912
rect 13558 56864 13610 56912
rect 13310 56860 13362 56864
rect 13434 56860 13486 56864
rect 13558 56860 13610 56864
rect 2682 56690 2727 56715
rect 2727 56690 2838 56715
rect 2682 56588 2838 56690
rect 2682 56559 2727 56588
rect 2727 56559 2838 56588
rect 3682 56690 3793 56715
rect 3793 56690 3838 56715
rect 3682 56588 3838 56690
rect 3682 56559 3793 56588
rect 3793 56559 3838 56588
rect 4182 56690 4227 56715
rect 4227 56690 4338 56715
rect 4182 56588 4338 56690
rect 4182 56559 4227 56588
rect 4227 56559 4338 56588
rect 5182 56690 5293 56715
rect 5293 56690 5338 56715
rect 5182 56588 5338 56690
rect 5182 56559 5293 56588
rect 5293 56559 5338 56588
rect 5682 56690 5727 56715
rect 5727 56690 5838 56715
rect 5682 56588 5838 56690
rect 5682 56559 5727 56588
rect 5727 56559 5838 56588
rect 6682 56690 6793 56715
rect 6793 56690 6838 56715
rect 6682 56588 6838 56690
rect 6682 56559 6793 56588
rect 6793 56559 6838 56588
rect 7182 56690 7227 56715
rect 7227 56690 7338 56715
rect 7182 56588 7338 56690
rect 7182 56559 7227 56588
rect 7227 56559 7338 56588
rect 8182 56690 8293 56715
rect 8293 56690 8338 56715
rect 8182 56588 8338 56690
rect 8182 56559 8293 56588
rect 8293 56559 8338 56588
rect 8682 56690 8727 56715
rect 8727 56690 8838 56715
rect 8682 56588 8838 56690
rect 8682 56559 8727 56588
rect 8727 56559 8838 56588
rect 9682 56690 9793 56715
rect 9793 56690 9838 56715
rect 9682 56588 9838 56690
rect 9682 56559 9793 56588
rect 9793 56559 9838 56588
rect 10182 56690 10227 56715
rect 10227 56690 10338 56715
rect 10182 56588 10338 56690
rect 10182 56559 10227 56588
rect 10227 56559 10338 56588
rect 11182 56690 11293 56715
rect 11293 56690 11338 56715
rect 11182 56588 11338 56690
rect 11182 56559 11293 56588
rect 11293 56559 11338 56588
rect 11682 56690 11727 56715
rect 11727 56690 11838 56715
rect 11682 56588 11838 56690
rect 11682 56559 11727 56588
rect 11727 56559 11838 56588
rect 12682 56690 12793 56715
rect 12793 56690 12838 56715
rect 12682 56588 12838 56690
rect 12682 56559 12793 56588
rect 12793 56559 12838 56588
rect 13182 56690 13227 56715
rect 13227 56690 13338 56715
rect 13182 56588 13338 56690
rect 13182 56559 13227 56588
rect 13227 56559 13338 56588
rect 14392 56559 14548 56715
rect 2522 56366 2574 56418
rect 2646 56366 2698 56418
rect 2770 56414 2797 56418
rect 2797 56414 2822 56418
rect 2894 56414 2946 56418
rect 3018 56414 3070 56418
rect 3142 56414 3194 56418
rect 3266 56414 3318 56418
rect 3390 56414 3442 56418
rect 3514 56414 3566 56418
rect 3638 56414 3690 56418
rect 2770 56366 2822 56414
rect 2894 56366 2946 56414
rect 3018 56366 3070 56414
rect 3142 56366 3194 56414
rect 3266 56366 3318 56414
rect 3390 56366 3442 56414
rect 3514 56366 3566 56414
rect 3638 56366 3690 56414
rect 3762 56366 3814 56418
rect 3886 56366 3938 56418
rect 4010 56366 4062 56418
rect 4134 56366 4186 56418
rect 4258 56414 4297 56418
rect 4297 56414 4310 56418
rect 4382 56414 4434 56418
rect 4506 56414 4558 56418
rect 4630 56414 4682 56418
rect 4754 56414 4806 56418
rect 4878 56414 4930 56418
rect 5002 56414 5054 56418
rect 5126 56414 5178 56418
rect 4258 56366 4310 56414
rect 4382 56366 4434 56414
rect 4506 56366 4558 56414
rect 4630 56366 4682 56414
rect 4754 56366 4806 56414
rect 4878 56366 4930 56414
rect 5002 56366 5054 56414
rect 5126 56366 5178 56414
rect 5250 56366 5302 56418
rect 5374 56366 5426 56418
rect 5498 56366 5550 56418
rect 5622 56366 5674 56418
rect 5746 56414 5797 56418
rect 5797 56414 5798 56418
rect 5870 56414 5922 56418
rect 5994 56414 6046 56418
rect 6118 56414 6170 56418
rect 6242 56414 6294 56418
rect 6366 56414 6418 56418
rect 6490 56414 6542 56418
rect 6614 56414 6666 56418
rect 5746 56366 5798 56414
rect 5870 56366 5922 56414
rect 5994 56366 6046 56414
rect 6118 56366 6170 56414
rect 6242 56366 6294 56414
rect 6366 56366 6418 56414
rect 6490 56366 6542 56414
rect 6614 56366 6666 56414
rect 6738 56366 6790 56418
rect 6862 56366 6914 56418
rect 6986 56366 7038 56418
rect 7110 56366 7162 56418
rect 7234 56366 7286 56418
rect 7358 56414 7410 56418
rect 7482 56414 7534 56418
rect 7606 56414 7658 56418
rect 7730 56414 7782 56418
rect 7854 56414 7906 56418
rect 7978 56414 8030 56418
rect 8102 56414 8154 56418
rect 7358 56366 7410 56414
rect 7482 56366 7534 56414
rect 7606 56366 7658 56414
rect 7730 56366 7782 56414
rect 7854 56366 7906 56414
rect 7978 56366 8030 56414
rect 8102 56366 8154 56414
rect 8226 56366 8278 56418
rect 8350 56366 8402 56418
rect 8474 56366 8526 56418
rect 8598 56366 8650 56418
rect 8722 56366 8774 56418
rect 8846 56414 8898 56418
rect 8970 56414 9022 56418
rect 9094 56414 9146 56418
rect 9218 56414 9270 56418
rect 9342 56414 9394 56418
rect 9466 56414 9518 56418
rect 9590 56414 9642 56418
rect 9714 56414 9723 56418
rect 9723 56414 9766 56418
rect 8846 56366 8898 56414
rect 8970 56366 9022 56414
rect 9094 56366 9146 56414
rect 9218 56366 9270 56414
rect 9342 56366 9394 56414
rect 9466 56366 9518 56414
rect 9590 56366 9642 56414
rect 9714 56366 9766 56414
rect 9838 56366 9890 56418
rect 9962 56366 10014 56418
rect 10086 56366 10138 56418
rect 10210 56366 10262 56418
rect 10334 56414 10386 56418
rect 10458 56414 10510 56418
rect 10582 56414 10634 56418
rect 10706 56414 10758 56418
rect 10830 56414 10882 56418
rect 10954 56414 11006 56418
rect 11078 56414 11130 56418
rect 11202 56414 11223 56418
rect 11223 56414 11254 56418
rect 10334 56366 10386 56414
rect 10458 56366 10510 56414
rect 10582 56366 10634 56414
rect 10706 56366 10758 56414
rect 10830 56366 10882 56414
rect 10954 56366 11006 56414
rect 11078 56366 11130 56414
rect 11202 56366 11254 56414
rect 11326 56366 11378 56418
rect 11450 56366 11502 56418
rect 11574 56366 11626 56418
rect 11698 56366 11750 56418
rect 11822 56414 11874 56418
rect 11946 56414 11998 56418
rect 12070 56414 12122 56418
rect 12194 56414 12246 56418
rect 12318 56414 12370 56418
rect 12442 56414 12494 56418
rect 12566 56414 12618 56418
rect 12690 56414 12723 56418
rect 12723 56414 12742 56418
rect 11822 56366 11874 56414
rect 11946 56366 11998 56414
rect 12070 56366 12122 56414
rect 12194 56366 12246 56414
rect 12318 56366 12370 56414
rect 12442 56366 12494 56414
rect 12566 56366 12618 56414
rect 12690 56366 12742 56414
rect 12814 56366 12866 56418
rect 12938 56366 12990 56418
rect 13062 56366 13114 56418
rect 13186 56366 13238 56418
rect 13310 56414 13362 56418
rect 13434 56414 13486 56418
rect 13558 56414 13610 56418
rect 13310 56366 13362 56414
rect 13434 56366 13486 56414
rect 13558 56366 13610 56414
rect 2522 56242 2574 56294
rect 2646 56242 2698 56294
rect 2770 56242 2822 56294
rect 2894 56242 2946 56294
rect 3018 56242 3070 56294
rect 3142 56242 3194 56294
rect 3266 56242 3318 56294
rect 3390 56242 3442 56294
rect 3514 56242 3566 56294
rect 3638 56242 3690 56294
rect 3762 56242 3814 56294
rect 3886 56242 3938 56294
rect 4010 56242 4062 56294
rect 4134 56242 4186 56294
rect 4258 56242 4310 56294
rect 4382 56242 4434 56294
rect 4506 56242 4558 56294
rect 4630 56242 4682 56294
rect 4754 56242 4806 56294
rect 4878 56242 4930 56294
rect 5002 56242 5054 56294
rect 5126 56242 5178 56294
rect 5250 56242 5302 56294
rect 5374 56242 5426 56294
rect 5498 56242 5550 56294
rect 5622 56242 5674 56294
rect 5746 56242 5798 56294
rect 5870 56242 5922 56294
rect 5994 56242 6046 56294
rect 6118 56242 6170 56294
rect 6242 56242 6294 56294
rect 6366 56242 6418 56294
rect 6490 56242 6542 56294
rect 6614 56242 6666 56294
rect 6738 56242 6790 56294
rect 6862 56242 6914 56294
rect 6986 56242 7038 56294
rect 7110 56242 7162 56294
rect 7234 56242 7286 56294
rect 7358 56242 7410 56294
rect 7482 56242 7534 56294
rect 7606 56242 7658 56294
rect 7730 56242 7782 56294
rect 7854 56242 7906 56294
rect 7978 56242 8030 56294
rect 8102 56242 8154 56294
rect 8226 56242 8278 56294
rect 8350 56242 8402 56294
rect 8474 56242 8526 56294
rect 8598 56242 8650 56294
rect 8722 56242 8774 56294
rect 8846 56242 8898 56294
rect 8970 56242 9022 56294
rect 9094 56242 9146 56294
rect 9218 56242 9270 56294
rect 9342 56242 9394 56294
rect 9466 56242 9518 56294
rect 9590 56242 9642 56294
rect 9714 56242 9766 56294
rect 9838 56242 9890 56294
rect 9962 56242 10014 56294
rect 10086 56242 10138 56294
rect 10210 56242 10262 56294
rect 10334 56242 10386 56294
rect 10458 56242 10510 56294
rect 10582 56242 10634 56294
rect 10706 56242 10758 56294
rect 10830 56242 10882 56294
rect 10954 56242 11006 56294
rect 11078 56242 11130 56294
rect 11202 56242 11254 56294
rect 11326 56242 11378 56294
rect 11450 56242 11502 56294
rect 11574 56242 11626 56294
rect 11698 56242 11750 56294
rect 11822 56242 11874 56294
rect 11946 56242 11998 56294
rect 12070 56242 12122 56294
rect 12194 56242 12246 56294
rect 12318 56242 12370 56294
rect 12442 56242 12494 56294
rect 12566 56242 12618 56294
rect 12690 56242 12742 56294
rect 12814 56242 12866 56294
rect 12938 56242 12990 56294
rect 13062 56242 13114 56294
rect 13186 56242 13238 56294
rect 13310 56242 13362 56294
rect 13434 56242 13486 56294
rect 13558 56242 13610 56294
rect 2522 56122 2574 56170
rect 2646 56122 2698 56170
rect 2770 56122 2822 56170
rect 2894 56122 2946 56170
rect 3018 56122 3070 56170
rect 3142 56122 3194 56170
rect 3266 56122 3318 56170
rect 3390 56122 3442 56170
rect 3514 56122 3566 56170
rect 3638 56122 3690 56170
rect 3762 56122 3814 56170
rect 3886 56122 3938 56170
rect 4010 56122 4062 56170
rect 4134 56122 4186 56170
rect 4258 56122 4310 56170
rect 4382 56122 4434 56170
rect 4506 56122 4558 56170
rect 4630 56122 4682 56170
rect 4754 56122 4806 56170
rect 4878 56122 4930 56170
rect 5002 56122 5054 56170
rect 5126 56122 5178 56170
rect 5250 56122 5302 56170
rect 5374 56122 5426 56170
rect 5498 56122 5550 56170
rect 5622 56122 5674 56170
rect 5746 56122 5798 56170
rect 5870 56122 5922 56170
rect 5994 56122 6046 56170
rect 6118 56122 6170 56170
rect 6242 56122 6294 56170
rect 6366 56122 6418 56170
rect 6490 56122 6542 56170
rect 6614 56122 6666 56170
rect 6738 56122 6790 56170
rect 6862 56122 6914 56170
rect 6986 56122 7038 56170
rect 7110 56122 7162 56170
rect 7234 56122 7286 56170
rect 7358 56122 7410 56170
rect 7482 56122 7534 56170
rect 7606 56122 7658 56170
rect 7730 56122 7782 56170
rect 7854 56122 7906 56170
rect 7978 56122 8030 56170
rect 8102 56122 8154 56170
rect 8226 56122 8278 56170
rect 8350 56122 8402 56170
rect 8474 56122 8526 56170
rect 8598 56122 8650 56170
rect 8722 56122 8774 56170
rect 8846 56122 8898 56170
rect 8970 56122 9022 56170
rect 9094 56122 9146 56170
rect 9218 56122 9270 56170
rect 9342 56122 9394 56170
rect 9466 56122 9518 56170
rect 9590 56122 9642 56170
rect 9714 56122 9766 56170
rect 9838 56122 9890 56170
rect 9962 56122 10014 56170
rect 10086 56122 10138 56170
rect 10210 56122 10262 56170
rect 10334 56122 10386 56170
rect 10458 56122 10510 56170
rect 10582 56122 10634 56170
rect 10706 56122 10758 56170
rect 10830 56122 10882 56170
rect 10954 56122 11006 56170
rect 11078 56122 11130 56170
rect 11202 56122 11254 56170
rect 11326 56122 11378 56170
rect 11450 56122 11502 56170
rect 11574 56122 11626 56170
rect 11698 56122 11750 56170
rect 11822 56122 11874 56170
rect 11946 56122 11998 56170
rect 12070 56122 12122 56170
rect 12194 56122 12246 56170
rect 12318 56122 12370 56170
rect 12442 56122 12494 56170
rect 12566 56122 12618 56170
rect 12690 56122 12742 56170
rect 12814 56122 12866 56170
rect 12938 56122 12990 56170
rect 13062 56122 13114 56170
rect 13186 56122 13238 56170
rect 13310 56122 13362 56170
rect 13434 56122 13486 56170
rect 13558 56122 13610 56170
rect 2522 56118 2574 56122
rect 2646 56118 2698 56122
rect 2770 56118 2822 56122
rect 2894 56118 2946 56122
rect 3018 56118 3070 56122
rect 3142 56118 3194 56122
rect 3266 56118 3318 56122
rect 3390 56118 3442 56122
rect 3514 56118 3566 56122
rect 3638 56118 3690 56122
rect 3762 56118 3814 56122
rect 3886 56118 3938 56122
rect 4010 56118 4062 56122
rect 4134 56118 4186 56122
rect 4258 56118 4310 56122
rect 4382 56118 4434 56122
rect 4506 56118 4558 56122
rect 4630 56118 4682 56122
rect 4754 56118 4806 56122
rect 4878 56118 4930 56122
rect 5002 56118 5054 56122
rect 5126 56118 5178 56122
rect 5250 56118 5302 56122
rect 5374 56118 5426 56122
rect 5498 56118 5550 56122
rect 5622 56118 5674 56122
rect 5746 56118 5798 56122
rect 5870 56118 5922 56122
rect 5994 56118 6046 56122
rect 6118 56118 6170 56122
rect 6242 56118 6294 56122
rect 6366 56118 6418 56122
rect 6490 56118 6542 56122
rect 6614 56118 6666 56122
rect 6738 56118 6790 56122
rect 6862 56118 6914 56122
rect 6986 56118 7038 56122
rect 7110 56118 7162 56122
rect 7234 56118 7286 56122
rect 7358 56118 7410 56122
rect 7482 56118 7534 56122
rect 7606 56118 7658 56122
rect 7730 56118 7782 56122
rect 7854 56118 7906 56122
rect 7978 56118 8030 56122
rect 8102 56118 8154 56122
rect 8226 56118 8278 56122
rect 8350 56118 8402 56122
rect 8474 56118 8526 56122
rect 8598 56118 8650 56122
rect 8722 56118 8774 56122
rect 8846 56118 8898 56122
rect 8970 56118 9022 56122
rect 9094 56118 9146 56122
rect 9218 56118 9270 56122
rect 9342 56118 9394 56122
rect 9466 56118 9518 56122
rect 9590 56118 9642 56122
rect 9714 56118 9766 56122
rect 9838 56118 9890 56122
rect 9962 56118 10014 56122
rect 10086 56118 10138 56122
rect 10210 56118 10262 56122
rect 10334 56118 10386 56122
rect 10458 56118 10510 56122
rect 10582 56118 10634 56122
rect 10706 56118 10758 56122
rect 10830 56118 10882 56122
rect 10954 56118 11006 56122
rect 11078 56118 11130 56122
rect 11202 56118 11254 56122
rect 11326 56118 11378 56122
rect 11450 56118 11502 56122
rect 11574 56118 11626 56122
rect 11698 56118 11750 56122
rect 11822 56118 11874 56122
rect 11946 56118 11998 56122
rect 12070 56118 12122 56122
rect 12194 56118 12246 56122
rect 12318 56118 12370 56122
rect 12442 56118 12494 56122
rect 12566 56118 12618 56122
rect 12690 56118 12742 56122
rect 12814 56118 12866 56122
rect 12938 56118 12990 56122
rect 13062 56118 13114 56122
rect 13186 56118 13238 56122
rect 13310 56118 13362 56122
rect 13434 56118 13486 56122
rect 13558 56118 13610 56122
rect 3512 55785 4084 55837
rect 2321 55555 2373 55711
rect 2605 55411 2761 55463
rect 234 55043 286 55095
rect 358 55043 410 55095
rect 482 55043 534 55095
rect 234 54919 286 54971
rect 358 54919 410 54971
rect 482 54919 534 54971
rect 234 54795 286 54847
rect 358 54795 410 54847
rect 482 54795 534 54847
rect 4762 54845 4814 55729
rect 4950 54978 5002 55758
rect 5438 54987 5490 55767
rect 5926 54987 5978 55767
rect 6108 54845 6160 55729
rect 6290 54987 6342 55767
rect 6778 54987 6830 55767
rect 7266 54987 7318 55767
rect 7454 54845 7506 55729
rect 8042 54841 8094 55829
rect 8511 54841 8563 55829
rect 8726 54841 8778 55829
rect 8949 54841 9001 55829
rect 9418 54841 9470 55829
rect 10006 54845 10058 55729
rect 10194 54987 10246 55767
rect 10682 54987 10734 55767
rect 11170 54987 11222 55767
rect 11352 54845 11404 55729
rect 11534 54987 11586 55767
rect 12022 54987 12074 55767
rect 12510 54987 12562 55767
rect 12698 54845 12750 55729
rect 13286 54845 13338 55729
rect 234 54134 286 54186
rect 358 54134 410 54186
rect 482 54134 534 54186
rect 234 54010 286 54062
rect 358 54010 410 54062
rect 482 54010 534 54062
rect 234 53886 286 53938
rect 358 53886 410 53938
rect 482 53886 534 53938
rect 3482 53383 3534 54371
rect 4174 53383 4226 54163
rect 4762 53383 4814 54163
rect 4950 53430 5002 54002
rect 5438 53430 5490 54002
rect 5926 53430 5978 54002
rect 6108 53383 6160 54267
rect 6290 53430 6342 54002
rect 6778 53430 6830 54002
rect 7266 53430 7318 54002
rect 7454 53383 7506 54163
rect 8042 53383 8094 54163
rect 8730 53383 8782 54371
rect 10006 53383 10058 54163
rect 10194 53430 10246 54002
rect 10682 53430 10734 54002
rect 11170 53430 11222 54002
rect 11352 53383 11404 54267
rect 11534 53430 11586 54002
rect 12022 53430 12074 54002
rect 12510 53430 12562 54002
rect 12698 53383 12750 54163
rect 13286 53383 13338 54163
rect 722 52955 1086 53007
rect 3378 52955 3534 53007
rect 3695 52955 3851 53007
rect 4746 52627 5214 52679
rect 6450 52627 6918 52679
rect 7266 52627 7422 52679
rect 58 51243 110 52543
rect 14954 51295 15006 52491
rect 1864 50217 6804 50269
rect 7732 50217 8096 50269
rect 8434 50217 8798 50269
rect 4644 49372 4696 49424
rect 4768 49372 4820 49424
rect 4892 49372 4944 49424
rect 4644 49248 4696 49300
rect 4768 49248 4820 49300
rect 4892 49248 4944 49300
rect 4644 49124 4696 49176
rect 4768 49124 4820 49176
rect 4892 49124 4944 49176
rect 5531 49138 5895 49398
rect 6434 49138 6798 49398
rect 7732 49138 8096 49398
rect 8434 49138 8798 49398
rect 4644 49000 4696 49052
rect 4768 49000 4820 49052
rect 4892 49000 4944 49052
rect 4644 48876 4696 48928
rect 4768 48876 4820 48928
rect 4892 48876 4944 48928
rect 4644 48752 4696 48804
rect 4768 48752 4820 48804
rect 4892 48752 4944 48804
rect 4644 48628 4696 48680
rect 4768 48628 4820 48680
rect 4892 48628 4944 48680
rect 4644 48504 4696 48556
rect 4768 48504 4820 48556
rect 4892 48504 4944 48556
rect 4644 48380 4696 48432
rect 4768 48380 4820 48432
rect 4892 48380 4944 48432
rect 10794 48372 10846 49360
rect 14392 49252 14444 49304
rect 14500 49252 14552 49304
rect 14392 49144 14444 49196
rect 14500 49144 14552 49196
rect 14392 49036 14444 49088
rect 14500 49036 14552 49088
rect 14392 48928 14444 48980
rect 14500 48928 14552 48980
rect 14392 48820 14444 48872
rect 14500 48820 14552 48872
rect 4644 48256 4696 48308
rect 4768 48256 4820 48308
rect 4892 48256 4944 48308
rect 4644 48132 4696 48184
rect 4768 48132 4820 48184
rect 4892 48132 4944 48184
rect 4644 48008 4696 48060
rect 4768 48008 4820 48060
rect 4892 48008 4944 48060
rect 14392 48284 14444 48336
rect 14500 48284 14552 48336
rect 14392 48176 14444 48228
rect 14500 48176 14552 48228
rect 14392 48068 14444 48120
rect 14500 48068 14552 48120
rect 14392 47960 14444 48012
rect 14500 47960 14552 48012
rect 4644 47884 4696 47936
rect 4768 47884 4820 47936
rect 4892 47884 4944 47936
rect 3620 46696 3672 47788
rect 11630 47786 11682 47942
rect 14392 47852 14444 47904
rect 14500 47852 14552 47904
rect 11013 47146 11065 47718
rect 3197 46036 3353 46504
rect 12272 46914 12324 46966
rect 12380 46914 12432 46966
rect 12488 46914 12540 46966
rect 12596 46914 12648 46966
rect 14216 45837 14268 45993
rect 3620 43243 3672 44543
rect 12434 44001 12590 44053
rect 3620 41643 3672 42943
rect 11583 41814 11635 41815
rect 11583 41768 11599 41814
rect 11599 41768 11635 41814
rect 11583 41686 11635 41768
rect 11583 41659 11599 41686
rect 11599 41659 11635 41686
rect 11583 41304 11599 41341
rect 11599 41304 11635 41341
rect 11583 41222 11635 41304
rect 11583 41185 11599 41222
rect 11599 41185 11635 41222
rect 1848 41018 3668 41070
rect 11298 41124 11303 41163
rect 11303 41124 11349 41163
rect 11349 41124 11350 41163
rect 11298 41054 11350 41124
rect 13108 42839 13160 42868
rect 13108 42793 13115 42839
rect 13115 42793 13160 42839
rect 13108 42727 13160 42793
rect 13108 42712 13115 42727
rect 13115 42712 13160 42727
rect 13544 42839 13596 42868
rect 13544 42793 13589 42839
rect 13589 42793 13596 42839
rect 13544 42727 13596 42793
rect 13544 42712 13589 42727
rect 13589 42712 13596 42727
rect 13108 41937 13115 41941
rect 13115 41937 13160 41941
rect 13108 41871 13160 41937
rect 13108 41825 13115 41871
rect 13115 41825 13160 41871
rect 13108 41785 13160 41825
rect 13544 41937 13589 41941
rect 13589 41937 13596 41941
rect 13544 41871 13596 41937
rect 13544 41825 13589 41871
rect 13589 41825 13596 41871
rect 13544 41785 13596 41825
rect 11298 41008 11303 41054
rect 11303 41008 11349 41054
rect 11349 41008 11350 41054
rect 11298 41007 11350 41008
rect 11029 40816 11081 40972
rect 11714 40831 11870 40883
rect 1925 40682 2081 40734
rect 4849 40682 5005 40734
rect 7065 40682 7221 40734
rect 10900 40682 11056 40734
rect 14070 40682 14122 40838
rect 1608 40516 1764 40568
rect 5578 40516 5734 40568
rect 11428 40546 11584 40598
rect 13674 40546 13830 40598
rect 10656 40410 10812 40462
rect 11996 40410 12152 40462
rect 13820 40410 13976 40462
rect 202 40254 566 40306
rect 2445 40262 4473 40314
rect 7900 40262 9720 40314
rect 12784 40262 13772 40314
rect 1783 39216 1835 39788
rect 5095 39186 5147 39758
rect 6061 38770 6113 39758
rect 7027 39186 7079 39758
rect 10339 38800 10391 39788
rect 10656 38890 10708 39046
rect 10900 38890 10952 39046
rect 11212 38800 11264 39788
rect 8305 38532 8357 38688
rect 58 36843 110 38143
rect 817 37524 869 38512
rect 2719 37783 2771 37939
rect 3207 37783 3259 37939
rect 3439 37524 3491 38512
rect 11532 38529 11584 38685
rect 3671 37783 3723 37939
rect 4159 37783 4211 37939
rect 6061 37524 6113 38512
rect 13315 38519 13367 38675
rect 8451 37783 8503 37939
rect 8683 37524 8735 38512
rect 8907 37783 8959 37939
rect 13451 37867 13503 38023
rect 10343 37516 11539 37568
rect 8451 36846 8503 37002
rect 13074 36846 13230 36898
rect 8305 36710 8461 36762
rect 12934 36710 13090 36762
rect 2088 36574 2452 36626
rect 4473 36574 4629 36626
rect 5822 36574 5978 36626
rect 8982 36574 9138 36626
rect 1834 36438 1990 36490
rect 3103 36438 3259 36490
rect 3671 36438 3827 36490
rect 6066 36438 6222 36490
rect 8842 36438 8998 36490
rect 2494 36302 2650 36354
rect 5406 36302 5562 36354
rect 9502 36302 9658 36354
rect 12518 36302 12674 36354
rect 1322 36166 1478 36218
rect 6578 36166 6734 36218
rect 8330 36166 8486 36218
rect 13586 36166 13742 36218
rect 3398 36030 3554 36082
rect 4502 36030 4658 36082
rect 10406 36030 10562 36082
rect 11510 36030 11666 36082
rect 13347 36030 13503 36082
rect 498 34126 550 35946
rect 736 34542 788 35946
rect 3104 34542 3156 35946
rect 1834 34279 1886 34435
rect 2078 34279 2130 34435
rect 2494 34279 2546 34435
rect 498 30055 550 33851
rect 4002 33294 4054 35946
rect 4900 34542 4952 35946
rect 8579 35894 8735 35946
rect 10112 34542 10164 35946
rect 5510 34279 5562 34435
rect 5926 34279 5978 34435
rect 6170 34279 6222 34435
rect 8842 34279 8894 34435
rect 9086 34279 9138 34435
rect 9502 34279 9554 34435
rect 11010 33294 11062 35946
rect 11908 34542 11960 35946
rect 14954 36843 15006 38143
rect 12518 34279 12570 34435
rect 12934 34279 12986 34435
rect 13178 34279 13230 34435
rect 980 30454 1032 32690
rect 1468 30314 1520 30678
rect 1712 30314 1764 30678
rect 2372 30454 2424 32690
rect 2788 30454 2840 32690
rect 3276 31078 3328 32690
rect 3764 31028 3816 32640
rect 4002 31005 4054 32825
rect 4240 31028 4292 32640
rect 4728 31078 4780 32690
rect 5216 31078 5268 32690
rect 5632 31078 5684 32690
rect 3032 30494 3084 30858
rect 3520 30314 3572 30678
rect 4484 30494 4536 30858
rect 4972 30314 5024 30678
rect 6536 30314 6588 30678
rect 6780 30314 6832 30678
rect 7024 30454 7076 32690
rect 7988 30454 8040 32690
rect 9380 31078 9432 32690
rect 9796 31078 9848 32690
rect 10284 31078 10336 32690
rect 10772 31028 10824 32640
rect 11010 31005 11062 32825
rect 11248 31028 11300 32640
rect 11736 31078 11788 32690
rect 8476 30314 8528 30678
rect 8720 30314 8772 30678
rect 10040 30314 10092 30678
rect 10528 30494 10580 30858
rect 11492 30314 11544 30678
rect 11980 30494 12032 30858
rect 12224 30454 12276 32690
rect 12640 30454 12692 32690
rect 13544 30314 13596 30678
rect 13788 30314 13840 30678
rect 14032 30454 14084 32690
rect 2012 30055 3312 30107
rect 11949 30055 13249 30107
rect 14514 30055 14566 33851
rect 1379 29765 1535 29817
rect 6444 29765 6600 29817
rect 8708 29765 8864 29817
rect 13531 29765 13687 29817
rect 1559 29585 1715 29637
rect 6688 29585 6844 29637
rect 8464 29585 8620 29637
rect 13351 29585 13507 29637
rect 3508 29378 3664 29430
rect 4167 29313 4219 29469
rect 4972 29313 5024 29469
rect 5926 29313 5978 29469
rect 9088 29313 9140 29469
rect 10042 29313 10094 29469
rect 10847 29313 10899 29469
rect 11402 29378 11558 29430
<< metal2 >>
rect 704 57327 780 57339
rect 704 57171 716 57327
rect 768 57171 780 57327
rect 704 55400 780 57171
rect 1225 55400 1301 57600
rect 1454 57327 1672 57339
rect 1454 57275 1486 57327
rect 1642 57275 1672 57327
rect 1454 57263 1672 57275
rect 184 55095 584 55169
rect 184 55043 234 55095
rect 286 55043 358 55095
rect 410 55043 482 55095
rect 534 55043 584 55095
rect 184 54971 584 55043
rect 184 54919 234 54971
rect 286 54919 358 54971
rect 410 54919 482 54971
rect 534 54919 584 54971
rect 184 54847 584 54919
rect 184 54795 234 54847
rect 286 54795 358 54847
rect 410 54795 482 54847
rect 534 54795 584 54847
rect 184 54186 584 54795
rect 184 54134 234 54186
rect 286 54134 358 54186
rect 410 54134 482 54186
rect 534 54134 584 54186
rect 184 54062 584 54134
rect 184 54010 234 54062
rect 286 54010 358 54062
rect 410 54010 482 54062
rect 534 54010 584 54062
rect 184 53938 584 54010
rect 184 53886 234 53938
rect 286 53886 358 53938
rect 410 53886 482 53938
rect 534 53886 584 53938
rect 32 52567 122 52600
rect 32 52511 56 52567
rect 112 52511 122 52567
rect 32 52425 58 52511
rect 110 52425 122 52511
rect 32 52369 56 52425
rect 112 52369 122 52425
rect 32 52283 58 52369
rect 110 52283 122 52369
rect 32 52227 56 52283
rect 112 52227 122 52283
rect 32 52141 58 52227
rect 110 52141 122 52227
rect 32 52085 56 52141
rect 112 52085 122 52141
rect 32 51999 58 52085
rect 110 51999 122 52085
rect 32 51943 56 51999
rect 112 51943 122 51999
rect 32 51857 58 51943
rect 110 51857 122 51943
rect 32 51801 56 51857
rect 112 51801 122 51857
rect 32 51715 58 51801
rect 110 51715 122 51801
rect 32 51659 56 51715
rect 112 51659 122 51715
rect 32 51573 58 51659
rect 110 51573 122 51659
rect 32 51517 56 51573
rect 112 51517 122 51573
rect 32 51431 58 51517
rect 110 51431 122 51517
rect 32 51375 56 51431
rect 112 51375 122 51431
rect 32 51289 58 51375
rect 110 51289 122 51375
rect 32 51233 56 51289
rect 112 51233 122 51289
rect 32 51200 122 51233
rect 184 50960 584 53886
rect 184 50904 214 50960
rect 270 50904 356 50960
rect 412 50904 498 50960
rect 554 50904 584 50960
rect 184 50818 584 50904
rect 184 50762 214 50818
rect 270 50762 356 50818
rect 412 50762 498 50818
rect 554 50762 584 50818
rect 184 50676 584 50762
rect 184 50620 214 50676
rect 270 50620 356 50676
rect 412 50620 498 50676
rect 554 50620 584 50676
rect 184 50534 584 50620
rect 184 50478 214 50534
rect 270 50478 356 50534
rect 412 50478 498 50534
rect 554 50478 584 50534
rect 184 50392 584 50478
rect 184 50336 214 50392
rect 270 50336 356 50392
rect 412 50336 498 50392
rect 554 50336 584 50392
rect 184 50250 584 50336
rect 184 50194 214 50250
rect 270 50194 356 50250
rect 412 50194 498 50250
rect 554 50194 584 50250
rect 184 50108 584 50194
rect 184 50052 214 50108
rect 270 50052 356 50108
rect 412 50052 498 50108
rect 554 50052 584 50108
rect 184 49966 584 50052
rect 184 49910 214 49966
rect 270 49910 356 49966
rect 412 49910 498 49966
rect 554 49910 584 49966
rect 184 49824 584 49910
rect 184 49768 214 49824
rect 270 49768 356 49824
rect 412 49768 498 49824
rect 554 49768 584 49824
rect 184 49682 584 49768
rect 184 49626 214 49682
rect 270 49626 356 49682
rect 412 49626 498 49682
rect 554 49626 584 49682
rect 184 40306 584 49626
rect 184 40254 202 40306
rect 566 40254 584 40306
rect 184 39760 584 40254
rect 184 39704 214 39760
rect 270 39704 356 39760
rect 412 39704 498 39760
rect 554 39704 584 39760
rect 184 39618 584 39704
rect 184 39562 214 39618
rect 270 39562 356 39618
rect 412 39562 498 39618
rect 554 39562 584 39618
rect 184 39476 584 39562
rect 184 39420 214 39476
rect 270 39420 356 39476
rect 412 39420 498 39476
rect 554 39420 584 39476
rect 184 39334 584 39420
rect 184 39278 214 39334
rect 270 39278 356 39334
rect 412 39278 498 39334
rect 554 39278 584 39334
rect 184 39192 584 39278
rect 184 39136 214 39192
rect 270 39136 356 39192
rect 412 39136 498 39192
rect 554 39136 584 39192
rect 184 39050 584 39136
rect 184 38994 214 39050
rect 270 38994 356 39050
rect 412 38994 498 39050
rect 554 38994 584 39050
rect 184 38908 584 38994
rect 184 38852 214 38908
rect 270 38852 356 38908
rect 412 38852 498 38908
rect 554 38852 584 38908
rect 184 38766 584 38852
rect 184 38710 214 38766
rect 270 38710 356 38766
rect 412 38710 498 38766
rect 554 38710 584 38766
rect 184 38624 584 38710
rect 184 38568 214 38624
rect 270 38568 356 38624
rect 412 38568 498 38624
rect 554 38568 584 38624
rect 184 38482 584 38568
rect 184 38426 214 38482
rect 270 38426 356 38482
rect 412 38426 498 38482
rect 554 38426 584 38482
rect 184 38400 584 38426
rect 704 53007 1104 53019
rect 704 52955 722 53007
rect 1086 52955 1104 53007
rect 704 52560 1104 52955
rect 704 52504 734 52560
rect 790 52504 876 52560
rect 932 52504 1018 52560
rect 1074 52504 1104 52560
rect 704 52418 1104 52504
rect 704 52362 734 52418
rect 790 52362 876 52418
rect 932 52362 1018 52418
rect 1074 52362 1104 52418
rect 704 52276 1104 52362
rect 704 52220 734 52276
rect 790 52220 876 52276
rect 932 52220 1018 52276
rect 1074 52220 1104 52276
rect 704 52134 1104 52220
rect 704 52078 734 52134
rect 790 52078 876 52134
rect 932 52078 1018 52134
rect 1074 52078 1104 52134
rect 704 51992 1104 52078
rect 704 51936 734 51992
rect 790 51936 876 51992
rect 932 51936 1018 51992
rect 1074 51936 1104 51992
rect 704 51850 1104 51936
rect 704 51794 734 51850
rect 790 51794 876 51850
rect 932 51794 1018 51850
rect 1074 51794 1104 51850
rect 704 51708 1104 51794
rect 704 51652 734 51708
rect 790 51652 876 51708
rect 932 51652 1018 51708
rect 1074 51652 1104 51708
rect 704 51566 1104 51652
rect 704 51510 734 51566
rect 790 51510 876 51566
rect 932 51510 1018 51566
rect 1074 51510 1104 51566
rect 704 51424 1104 51510
rect 704 51368 734 51424
rect 790 51368 876 51424
rect 932 51368 1018 51424
rect 1074 51368 1104 51424
rect 704 51282 1104 51368
rect 704 51226 734 51282
rect 790 51226 876 51282
rect 932 51226 1018 51282
rect 1074 51226 1104 51282
rect 704 38512 1104 51226
rect 1454 40579 1530 57263
rect 1184 40503 1530 40579
rect 1596 40580 1672 57263
rect 1886 57235 1962 57245
rect 1886 57179 1896 57235
rect 1952 57179 1962 57235
rect 1886 57093 1962 57179
rect 1886 57037 1896 57093
rect 1952 57037 1962 57093
rect 1886 56951 1962 57037
rect 1886 56895 1896 56951
rect 1952 56895 1962 56951
rect 1886 56809 1962 56895
rect 1886 56753 1896 56809
rect 1952 56753 1962 56809
rect 1886 56667 1962 56753
rect 1886 56611 1896 56667
rect 1952 56611 1962 56667
rect 1886 56525 1962 56611
rect 1886 56469 1896 56525
rect 1952 56469 1962 56525
rect 1886 56383 1962 56469
rect 1886 56327 1896 56383
rect 1952 56327 1962 56383
rect 1886 56241 1962 56327
rect 1886 56185 1896 56241
rect 1952 56185 1962 56241
rect 1886 56099 1962 56185
rect 1886 56043 1896 56099
rect 1952 56043 1962 56099
rect 1886 54160 1962 56043
rect 1886 54104 1896 54160
rect 1952 54104 1962 54160
rect 1886 54018 1962 54104
rect 1886 53962 1896 54018
rect 1952 53962 1962 54018
rect 1886 53876 1962 53962
rect 1886 53820 1896 53876
rect 1952 53820 1962 53876
rect 1886 53734 1962 53820
rect 1886 53678 1896 53734
rect 1952 53678 1962 53734
rect 1886 53592 1962 53678
rect 1886 53536 1896 53592
rect 1952 53536 1962 53592
rect 2098 53666 2174 57600
rect 13766 57327 14134 57339
rect 13766 57275 13822 57327
rect 14082 57275 14134 57327
rect 13766 57263 14134 57275
rect 2490 57180 13642 57190
rect 2490 57124 2500 57180
rect 2556 57160 2642 57180
rect 2698 57160 2784 57180
rect 2840 57160 2926 57180
rect 2982 57160 3068 57180
rect 3124 57160 3210 57180
rect 2574 57124 2642 57160
rect 2490 57108 2522 57124
rect 2574 57108 2646 57124
rect 2698 57108 2770 57160
rect 2840 57124 2894 57160
rect 2982 57124 3018 57160
rect 3124 57124 3142 57160
rect 2822 57108 2894 57124
rect 2946 57108 3018 57124
rect 3070 57108 3142 57124
rect 3194 57124 3210 57160
rect 3266 57160 3352 57180
rect 3408 57160 3494 57180
rect 3550 57160 3636 57180
rect 3692 57160 3778 57180
rect 3834 57160 3920 57180
rect 3976 57160 4062 57180
rect 3194 57108 3266 57124
rect 3318 57124 3352 57160
rect 3442 57124 3494 57160
rect 3566 57124 3636 57160
rect 3692 57124 3762 57160
rect 3834 57124 3886 57160
rect 3976 57124 4010 57160
rect 3318 57108 3390 57124
rect 3442 57108 3514 57124
rect 3566 57108 3638 57124
rect 3690 57108 3762 57124
rect 3814 57108 3886 57124
rect 3938 57108 4010 57124
rect 4118 57160 4204 57180
rect 4260 57160 4346 57180
rect 4402 57160 4488 57180
rect 4544 57160 4630 57180
rect 4686 57160 4772 57180
rect 4828 57160 4914 57180
rect 4970 57160 5056 57180
rect 4118 57124 4134 57160
rect 4062 57108 4134 57124
rect 4186 57124 4204 57160
rect 4310 57124 4346 57160
rect 4434 57124 4488 57160
rect 4186 57108 4258 57124
rect 4310 57108 4382 57124
rect 4434 57108 4506 57124
rect 4558 57108 4630 57160
rect 4686 57124 4754 57160
rect 4828 57124 4878 57160
rect 4970 57124 5002 57160
rect 4682 57108 4754 57124
rect 4806 57108 4878 57124
rect 4930 57108 5002 57124
rect 5054 57124 5056 57160
rect 5112 57160 5198 57180
rect 5254 57160 5340 57180
rect 5396 57160 5482 57180
rect 5538 57160 5624 57180
rect 5680 57160 5766 57180
rect 5822 57160 5908 57180
rect 5964 57160 6050 57180
rect 5112 57124 5126 57160
rect 5054 57108 5126 57124
rect 5178 57124 5198 57160
rect 5302 57124 5340 57160
rect 5426 57124 5482 57160
rect 5178 57108 5250 57124
rect 5302 57108 5374 57124
rect 5426 57108 5498 57124
rect 5550 57108 5622 57160
rect 5680 57124 5746 57160
rect 5822 57124 5870 57160
rect 5964 57124 5994 57160
rect 5674 57108 5746 57124
rect 5798 57108 5870 57124
rect 5922 57108 5994 57124
rect 6046 57124 6050 57160
rect 6106 57160 6192 57180
rect 6248 57160 6334 57180
rect 6390 57160 6476 57180
rect 6532 57160 6618 57180
rect 6674 57160 6760 57180
rect 6816 57160 6902 57180
rect 6958 57160 7044 57180
rect 6106 57124 6118 57160
rect 6046 57108 6118 57124
rect 6170 57124 6192 57160
rect 6294 57124 6334 57160
rect 6418 57124 6476 57160
rect 6170 57108 6242 57124
rect 6294 57108 6366 57124
rect 6418 57108 6490 57124
rect 6542 57108 6614 57160
rect 6674 57124 6738 57160
rect 6816 57124 6862 57160
rect 6958 57124 6986 57160
rect 6666 57108 6738 57124
rect 6790 57108 6862 57124
rect 6914 57108 6986 57124
rect 7038 57124 7044 57160
rect 7100 57160 7186 57180
rect 7242 57160 7328 57180
rect 7384 57160 7470 57180
rect 7526 57160 7612 57180
rect 7668 57160 7754 57180
rect 7810 57160 7896 57180
rect 7952 57160 8038 57180
rect 7100 57124 7110 57160
rect 7038 57108 7110 57124
rect 7162 57124 7186 57160
rect 7286 57124 7328 57160
rect 7410 57124 7470 57160
rect 7162 57108 7234 57124
rect 7286 57108 7358 57124
rect 7410 57108 7482 57124
rect 7534 57108 7606 57160
rect 7668 57124 7730 57160
rect 7810 57124 7854 57160
rect 7952 57124 7978 57160
rect 7658 57108 7730 57124
rect 7782 57108 7854 57124
rect 7906 57108 7978 57124
rect 8030 57124 8038 57160
rect 8094 57160 8180 57180
rect 8236 57160 8322 57180
rect 8378 57160 8464 57180
rect 8520 57160 8606 57180
rect 8662 57160 8748 57180
rect 8804 57160 8890 57180
rect 8946 57160 9032 57180
rect 8094 57124 8102 57160
rect 8030 57108 8102 57124
rect 8154 57124 8180 57160
rect 8278 57124 8322 57160
rect 8402 57124 8464 57160
rect 8154 57108 8226 57124
rect 8278 57108 8350 57124
rect 8402 57108 8474 57124
rect 8526 57108 8598 57160
rect 8662 57124 8722 57160
rect 8804 57124 8846 57160
rect 8946 57124 8970 57160
rect 8650 57108 8722 57124
rect 8774 57108 8846 57124
rect 8898 57108 8970 57124
rect 9022 57124 9032 57160
rect 9088 57160 9174 57180
rect 9230 57160 9316 57180
rect 9372 57160 9458 57180
rect 9514 57160 9600 57180
rect 9656 57160 9742 57180
rect 9798 57160 9884 57180
rect 9940 57160 10026 57180
rect 9088 57124 9094 57160
rect 9022 57108 9094 57124
rect 9146 57124 9174 57160
rect 9270 57124 9316 57160
rect 9394 57124 9458 57160
rect 9146 57108 9218 57124
rect 9270 57108 9342 57124
rect 9394 57108 9466 57124
rect 9518 57108 9590 57160
rect 9656 57124 9714 57160
rect 9798 57124 9838 57160
rect 9940 57124 9962 57160
rect 9642 57108 9714 57124
rect 9766 57108 9838 57124
rect 9890 57108 9962 57124
rect 10014 57124 10026 57160
rect 10082 57160 10168 57180
rect 10224 57160 10310 57180
rect 10366 57160 10452 57180
rect 10508 57160 10594 57180
rect 10650 57160 10736 57180
rect 10792 57160 10878 57180
rect 10934 57160 11020 57180
rect 10082 57124 10086 57160
rect 10014 57108 10086 57124
rect 10138 57124 10168 57160
rect 10262 57124 10310 57160
rect 10386 57124 10452 57160
rect 10138 57108 10210 57124
rect 10262 57108 10334 57124
rect 10386 57108 10458 57124
rect 10510 57108 10582 57160
rect 10650 57124 10706 57160
rect 10792 57124 10830 57160
rect 10934 57124 10954 57160
rect 10634 57108 10706 57124
rect 10758 57108 10830 57124
rect 10882 57108 10954 57124
rect 11006 57124 11020 57160
rect 11076 57160 11162 57180
rect 11218 57160 11304 57180
rect 11360 57160 11446 57180
rect 11502 57160 11588 57180
rect 11644 57160 11730 57180
rect 11786 57160 11872 57180
rect 11928 57160 12014 57180
rect 11076 57124 11078 57160
rect 11006 57108 11078 57124
rect 11130 57124 11162 57160
rect 11254 57124 11304 57160
rect 11378 57124 11446 57160
rect 11130 57108 11202 57124
rect 11254 57108 11326 57124
rect 11378 57108 11450 57124
rect 11502 57108 11574 57160
rect 11644 57124 11698 57160
rect 11786 57124 11822 57160
rect 11928 57124 11946 57160
rect 11626 57108 11698 57124
rect 11750 57108 11822 57124
rect 11874 57108 11946 57124
rect 11998 57124 12014 57160
rect 12070 57160 12156 57180
rect 12212 57160 12298 57180
rect 12354 57160 12440 57180
rect 12496 57160 12582 57180
rect 12638 57160 12724 57180
rect 12780 57160 12866 57180
rect 11998 57108 12070 57124
rect 12122 57124 12156 57160
rect 12246 57124 12298 57160
rect 12370 57124 12440 57160
rect 12496 57124 12566 57160
rect 12638 57124 12690 57160
rect 12780 57124 12814 57160
rect 12122 57108 12194 57124
rect 12246 57108 12318 57124
rect 12370 57108 12442 57124
rect 12494 57108 12566 57124
rect 12618 57108 12690 57124
rect 12742 57108 12814 57124
rect 12922 57160 13008 57180
rect 13064 57160 13150 57180
rect 13206 57160 13292 57180
rect 13348 57160 13434 57180
rect 13490 57160 13576 57180
rect 12922 57124 12938 57160
rect 12866 57108 12938 57124
rect 12990 57124 13008 57160
rect 13114 57124 13150 57160
rect 13238 57124 13292 57160
rect 12990 57108 13062 57124
rect 13114 57108 13186 57124
rect 13238 57108 13310 57124
rect 13362 57108 13434 57160
rect 13490 57124 13558 57160
rect 13632 57124 13642 57180
rect 13486 57108 13558 57124
rect 13610 57108 13642 57124
rect 2490 57038 13642 57108
rect 2490 56982 2500 57038
rect 2556 57036 2642 57038
rect 2698 57036 2784 57038
rect 2840 57036 2926 57038
rect 2982 57036 3068 57038
rect 3124 57036 3210 57038
rect 2574 56984 2642 57036
rect 2698 56984 2770 57036
rect 2840 56984 2894 57036
rect 2982 56984 3018 57036
rect 3124 56984 3142 57036
rect 3194 56984 3210 57036
rect 2556 56982 2642 56984
rect 2698 56982 2784 56984
rect 2840 56982 2926 56984
rect 2982 56982 3068 56984
rect 3124 56982 3210 56984
rect 3266 57036 3352 57038
rect 3408 57036 3494 57038
rect 3550 57036 3636 57038
rect 3692 57036 3778 57038
rect 3834 57036 3920 57038
rect 3976 57036 4062 57038
rect 3318 56984 3352 57036
rect 3442 56984 3494 57036
rect 3566 56984 3636 57036
rect 3692 56984 3762 57036
rect 3834 56984 3886 57036
rect 3976 56984 4010 57036
rect 3266 56982 3352 56984
rect 3408 56982 3494 56984
rect 3550 56982 3636 56984
rect 3692 56982 3778 56984
rect 3834 56982 3920 56984
rect 3976 56982 4062 56984
rect 4118 57036 4204 57038
rect 4260 57036 4346 57038
rect 4402 57036 4488 57038
rect 4544 57036 4630 57038
rect 4686 57036 4772 57038
rect 4828 57036 4914 57038
rect 4970 57036 5056 57038
rect 4118 56984 4134 57036
rect 4186 56984 4204 57036
rect 4310 56984 4346 57036
rect 4434 56984 4488 57036
rect 4558 56984 4630 57036
rect 4686 56984 4754 57036
rect 4828 56984 4878 57036
rect 4970 56984 5002 57036
rect 5054 56984 5056 57036
rect 4118 56982 4204 56984
rect 4260 56982 4346 56984
rect 4402 56982 4488 56984
rect 4544 56982 4630 56984
rect 4686 56982 4772 56984
rect 4828 56982 4914 56984
rect 4970 56982 5056 56984
rect 5112 57036 5198 57038
rect 5254 57036 5340 57038
rect 5396 57036 5482 57038
rect 5538 57036 5624 57038
rect 5680 57036 5766 57038
rect 5822 57036 5908 57038
rect 5964 57036 6050 57038
rect 5112 56984 5126 57036
rect 5178 56984 5198 57036
rect 5302 56984 5340 57036
rect 5426 56984 5482 57036
rect 5550 56984 5622 57036
rect 5680 56984 5746 57036
rect 5822 56984 5870 57036
rect 5964 56984 5994 57036
rect 6046 56984 6050 57036
rect 5112 56982 5198 56984
rect 5254 56982 5340 56984
rect 5396 56982 5482 56984
rect 5538 56982 5624 56984
rect 5680 56982 5766 56984
rect 5822 56982 5908 56984
rect 5964 56982 6050 56984
rect 6106 57036 6192 57038
rect 6248 57036 6334 57038
rect 6390 57036 6476 57038
rect 6532 57036 6618 57038
rect 6674 57036 6760 57038
rect 6816 57036 6902 57038
rect 6958 57036 7044 57038
rect 6106 56984 6118 57036
rect 6170 56984 6192 57036
rect 6294 56984 6334 57036
rect 6418 56984 6476 57036
rect 6542 56984 6614 57036
rect 6674 56984 6738 57036
rect 6816 56984 6862 57036
rect 6958 56984 6986 57036
rect 7038 56984 7044 57036
rect 6106 56982 6192 56984
rect 6248 56982 6334 56984
rect 6390 56982 6476 56984
rect 6532 56982 6618 56984
rect 6674 56982 6760 56984
rect 6816 56982 6902 56984
rect 6958 56982 7044 56984
rect 7100 57036 7186 57038
rect 7242 57036 7328 57038
rect 7384 57036 7470 57038
rect 7526 57036 7612 57038
rect 7668 57036 7754 57038
rect 7810 57036 7896 57038
rect 7952 57036 8038 57038
rect 7100 56984 7110 57036
rect 7162 56984 7186 57036
rect 7286 56984 7328 57036
rect 7410 56984 7470 57036
rect 7534 56984 7606 57036
rect 7668 56984 7730 57036
rect 7810 56984 7854 57036
rect 7952 56984 7978 57036
rect 8030 56984 8038 57036
rect 7100 56982 7186 56984
rect 7242 56982 7328 56984
rect 7384 56982 7470 56984
rect 7526 56982 7612 56984
rect 7668 56982 7754 56984
rect 7810 56982 7896 56984
rect 7952 56982 8038 56984
rect 8094 57036 8180 57038
rect 8236 57036 8322 57038
rect 8378 57036 8464 57038
rect 8520 57036 8606 57038
rect 8662 57036 8748 57038
rect 8804 57036 8890 57038
rect 8946 57036 9032 57038
rect 8094 56984 8102 57036
rect 8154 56984 8180 57036
rect 8278 56984 8322 57036
rect 8402 56984 8464 57036
rect 8526 56984 8598 57036
rect 8662 56984 8722 57036
rect 8804 56984 8846 57036
rect 8946 56984 8970 57036
rect 9022 56984 9032 57036
rect 8094 56982 8180 56984
rect 8236 56982 8322 56984
rect 8378 56982 8464 56984
rect 8520 56982 8606 56984
rect 8662 56982 8748 56984
rect 8804 56982 8890 56984
rect 8946 56982 9032 56984
rect 9088 57036 9174 57038
rect 9230 57036 9316 57038
rect 9372 57036 9458 57038
rect 9514 57036 9600 57038
rect 9656 57036 9742 57038
rect 9798 57036 9884 57038
rect 9940 57036 10026 57038
rect 9088 56984 9094 57036
rect 9146 56984 9174 57036
rect 9270 56984 9316 57036
rect 9394 56984 9458 57036
rect 9518 56984 9590 57036
rect 9656 56984 9714 57036
rect 9798 56984 9838 57036
rect 9940 56984 9962 57036
rect 10014 56984 10026 57036
rect 9088 56982 9174 56984
rect 9230 56982 9316 56984
rect 9372 56982 9458 56984
rect 9514 56982 9600 56984
rect 9656 56982 9742 56984
rect 9798 56982 9884 56984
rect 9940 56982 10026 56984
rect 10082 57036 10168 57038
rect 10224 57036 10310 57038
rect 10366 57036 10452 57038
rect 10508 57036 10594 57038
rect 10650 57036 10736 57038
rect 10792 57036 10878 57038
rect 10934 57036 11020 57038
rect 10082 56984 10086 57036
rect 10138 56984 10168 57036
rect 10262 56984 10310 57036
rect 10386 56984 10452 57036
rect 10510 56984 10582 57036
rect 10650 56984 10706 57036
rect 10792 56984 10830 57036
rect 10934 56984 10954 57036
rect 11006 56984 11020 57036
rect 10082 56982 10168 56984
rect 10224 56982 10310 56984
rect 10366 56982 10452 56984
rect 10508 56982 10594 56984
rect 10650 56982 10736 56984
rect 10792 56982 10878 56984
rect 10934 56982 11020 56984
rect 11076 57036 11162 57038
rect 11218 57036 11304 57038
rect 11360 57036 11446 57038
rect 11502 57036 11588 57038
rect 11644 57036 11730 57038
rect 11786 57036 11872 57038
rect 11928 57036 12014 57038
rect 11076 56984 11078 57036
rect 11130 56984 11162 57036
rect 11254 56984 11304 57036
rect 11378 56984 11446 57036
rect 11502 56984 11574 57036
rect 11644 56984 11698 57036
rect 11786 56984 11822 57036
rect 11928 56984 11946 57036
rect 11998 56984 12014 57036
rect 11076 56982 11162 56984
rect 11218 56982 11304 56984
rect 11360 56982 11446 56984
rect 11502 56982 11588 56984
rect 11644 56982 11730 56984
rect 11786 56982 11872 56984
rect 11928 56982 12014 56984
rect 12070 57036 12156 57038
rect 12212 57036 12298 57038
rect 12354 57036 12440 57038
rect 12496 57036 12582 57038
rect 12638 57036 12724 57038
rect 12780 57036 12866 57038
rect 12122 56984 12156 57036
rect 12246 56984 12298 57036
rect 12370 56984 12440 57036
rect 12496 56984 12566 57036
rect 12638 56984 12690 57036
rect 12780 56984 12814 57036
rect 12070 56982 12156 56984
rect 12212 56982 12298 56984
rect 12354 56982 12440 56984
rect 12496 56982 12582 56984
rect 12638 56982 12724 56984
rect 12780 56982 12866 56984
rect 12922 57036 13008 57038
rect 13064 57036 13150 57038
rect 13206 57036 13292 57038
rect 13348 57036 13434 57038
rect 13490 57036 13576 57038
rect 12922 56984 12938 57036
rect 12990 56984 13008 57036
rect 13114 56984 13150 57036
rect 13238 56984 13292 57036
rect 13362 56984 13434 57036
rect 13490 56984 13558 57036
rect 12922 56982 13008 56984
rect 13064 56982 13150 56984
rect 13206 56982 13292 56984
rect 13348 56982 13434 56984
rect 13490 56982 13576 56984
rect 13632 56982 13642 57038
rect 2490 56912 13642 56982
rect 2490 56896 2522 56912
rect 2574 56896 2646 56912
rect 2490 56840 2500 56896
rect 2574 56860 2642 56896
rect 2698 56860 2770 56912
rect 2822 56896 2894 56912
rect 2946 56896 3018 56912
rect 3070 56896 3142 56912
rect 2840 56860 2894 56896
rect 2982 56860 3018 56896
rect 3124 56860 3142 56896
rect 3194 56896 3266 56912
rect 3194 56860 3210 56896
rect 2556 56840 2642 56860
rect 2698 56840 2784 56860
rect 2840 56840 2926 56860
rect 2982 56840 3068 56860
rect 3124 56840 3210 56860
rect 3318 56896 3390 56912
rect 3442 56896 3514 56912
rect 3566 56896 3638 56912
rect 3690 56896 3762 56912
rect 3814 56896 3886 56912
rect 3938 56896 4010 56912
rect 3318 56860 3352 56896
rect 3442 56860 3494 56896
rect 3566 56860 3636 56896
rect 3692 56860 3762 56896
rect 3834 56860 3886 56896
rect 3976 56860 4010 56896
rect 4062 56896 4134 56912
rect 3266 56840 3352 56860
rect 3408 56840 3494 56860
rect 3550 56840 3636 56860
rect 3692 56840 3778 56860
rect 3834 56840 3920 56860
rect 3976 56840 4062 56860
rect 4118 56860 4134 56896
rect 4186 56896 4258 56912
rect 4310 56896 4382 56912
rect 4434 56896 4506 56912
rect 4186 56860 4204 56896
rect 4310 56860 4346 56896
rect 4434 56860 4488 56896
rect 4558 56860 4630 56912
rect 4682 56896 4754 56912
rect 4806 56896 4878 56912
rect 4930 56896 5002 56912
rect 4686 56860 4754 56896
rect 4828 56860 4878 56896
rect 4970 56860 5002 56896
rect 5054 56896 5126 56912
rect 5054 56860 5056 56896
rect 4118 56840 4204 56860
rect 4260 56840 4346 56860
rect 4402 56840 4488 56860
rect 4544 56840 4630 56860
rect 4686 56840 4772 56860
rect 4828 56840 4914 56860
rect 4970 56840 5056 56860
rect 5112 56860 5126 56896
rect 5178 56896 5250 56912
rect 5302 56896 5374 56912
rect 5426 56896 5498 56912
rect 5178 56860 5198 56896
rect 5302 56860 5340 56896
rect 5426 56860 5482 56896
rect 5550 56860 5622 56912
rect 5674 56896 5746 56912
rect 5798 56896 5870 56912
rect 5922 56896 5994 56912
rect 5680 56860 5746 56896
rect 5822 56860 5870 56896
rect 5964 56860 5994 56896
rect 6046 56896 6118 56912
rect 6046 56860 6050 56896
rect 5112 56840 5198 56860
rect 5254 56840 5340 56860
rect 5396 56840 5482 56860
rect 5538 56840 5624 56860
rect 5680 56840 5766 56860
rect 5822 56840 5908 56860
rect 5964 56840 6050 56860
rect 6106 56860 6118 56896
rect 6170 56896 6242 56912
rect 6294 56896 6366 56912
rect 6418 56896 6490 56912
rect 6170 56860 6192 56896
rect 6294 56860 6334 56896
rect 6418 56860 6476 56896
rect 6542 56860 6614 56912
rect 6666 56896 6738 56912
rect 6790 56896 6862 56912
rect 6914 56896 6986 56912
rect 6674 56860 6738 56896
rect 6816 56860 6862 56896
rect 6958 56860 6986 56896
rect 7038 56896 7110 56912
rect 7038 56860 7044 56896
rect 6106 56840 6192 56860
rect 6248 56840 6334 56860
rect 6390 56840 6476 56860
rect 6532 56840 6618 56860
rect 6674 56840 6760 56860
rect 6816 56840 6902 56860
rect 6958 56840 7044 56860
rect 7100 56860 7110 56896
rect 7162 56896 7234 56912
rect 7286 56896 7358 56912
rect 7410 56896 7482 56912
rect 7162 56860 7186 56896
rect 7286 56860 7328 56896
rect 7410 56860 7470 56896
rect 7534 56860 7606 56912
rect 7658 56896 7730 56912
rect 7782 56896 7854 56912
rect 7906 56896 7978 56912
rect 7668 56860 7730 56896
rect 7810 56860 7854 56896
rect 7952 56860 7978 56896
rect 8030 56896 8102 56912
rect 8030 56860 8038 56896
rect 7100 56840 7186 56860
rect 7242 56840 7328 56860
rect 7384 56840 7470 56860
rect 7526 56840 7612 56860
rect 7668 56840 7754 56860
rect 7810 56840 7896 56860
rect 7952 56840 8038 56860
rect 8094 56860 8102 56896
rect 8154 56896 8226 56912
rect 8278 56896 8350 56912
rect 8402 56896 8474 56912
rect 8154 56860 8180 56896
rect 8278 56860 8322 56896
rect 8402 56860 8464 56896
rect 8526 56860 8598 56912
rect 8650 56896 8722 56912
rect 8774 56896 8846 56912
rect 8898 56896 8970 56912
rect 8662 56860 8722 56896
rect 8804 56860 8846 56896
rect 8946 56860 8970 56896
rect 9022 56896 9094 56912
rect 9022 56860 9032 56896
rect 8094 56840 8180 56860
rect 8236 56840 8322 56860
rect 8378 56840 8464 56860
rect 8520 56840 8606 56860
rect 8662 56840 8748 56860
rect 8804 56840 8890 56860
rect 8946 56840 9032 56860
rect 9088 56860 9094 56896
rect 9146 56896 9218 56912
rect 9270 56896 9342 56912
rect 9394 56896 9466 56912
rect 9146 56860 9174 56896
rect 9270 56860 9316 56896
rect 9394 56860 9458 56896
rect 9518 56860 9590 56912
rect 9642 56896 9714 56912
rect 9766 56896 9838 56912
rect 9890 56896 9962 56912
rect 9656 56860 9714 56896
rect 9798 56860 9838 56896
rect 9940 56860 9962 56896
rect 10014 56896 10086 56912
rect 10014 56860 10026 56896
rect 9088 56840 9174 56860
rect 9230 56840 9316 56860
rect 9372 56840 9458 56860
rect 9514 56840 9600 56860
rect 9656 56840 9742 56860
rect 9798 56840 9884 56860
rect 9940 56840 10026 56860
rect 10082 56860 10086 56896
rect 10138 56896 10210 56912
rect 10262 56896 10334 56912
rect 10386 56896 10458 56912
rect 10138 56860 10168 56896
rect 10262 56860 10310 56896
rect 10386 56860 10452 56896
rect 10510 56860 10582 56912
rect 10634 56896 10706 56912
rect 10758 56896 10830 56912
rect 10882 56896 10954 56912
rect 10650 56860 10706 56896
rect 10792 56860 10830 56896
rect 10934 56860 10954 56896
rect 11006 56896 11078 56912
rect 11006 56860 11020 56896
rect 10082 56840 10168 56860
rect 10224 56840 10310 56860
rect 10366 56840 10452 56860
rect 10508 56840 10594 56860
rect 10650 56840 10736 56860
rect 10792 56840 10878 56860
rect 10934 56840 11020 56860
rect 11076 56860 11078 56896
rect 11130 56896 11202 56912
rect 11254 56896 11326 56912
rect 11378 56896 11450 56912
rect 11130 56860 11162 56896
rect 11254 56860 11304 56896
rect 11378 56860 11446 56896
rect 11502 56860 11574 56912
rect 11626 56896 11698 56912
rect 11750 56896 11822 56912
rect 11874 56896 11946 56912
rect 11644 56860 11698 56896
rect 11786 56860 11822 56896
rect 11928 56860 11946 56896
rect 11998 56896 12070 56912
rect 11998 56860 12014 56896
rect 11076 56840 11162 56860
rect 11218 56840 11304 56860
rect 11360 56840 11446 56860
rect 11502 56840 11588 56860
rect 11644 56840 11730 56860
rect 11786 56840 11872 56860
rect 11928 56840 12014 56860
rect 12122 56896 12194 56912
rect 12246 56896 12318 56912
rect 12370 56896 12442 56912
rect 12494 56896 12566 56912
rect 12618 56896 12690 56912
rect 12742 56896 12814 56912
rect 12122 56860 12156 56896
rect 12246 56860 12298 56896
rect 12370 56860 12440 56896
rect 12496 56860 12566 56896
rect 12638 56860 12690 56896
rect 12780 56860 12814 56896
rect 12866 56896 12938 56912
rect 12070 56840 12156 56860
rect 12212 56840 12298 56860
rect 12354 56840 12440 56860
rect 12496 56840 12582 56860
rect 12638 56840 12724 56860
rect 12780 56840 12866 56860
rect 12922 56860 12938 56896
rect 12990 56896 13062 56912
rect 13114 56896 13186 56912
rect 13238 56896 13310 56912
rect 12990 56860 13008 56896
rect 13114 56860 13150 56896
rect 13238 56860 13292 56896
rect 13362 56860 13434 56912
rect 13486 56896 13558 56912
rect 13610 56896 13642 56912
rect 13490 56860 13558 56896
rect 12922 56840 13008 56860
rect 13064 56840 13150 56860
rect 13206 56840 13292 56860
rect 13348 56840 13434 56860
rect 13490 56840 13576 56860
rect 13632 56840 13642 56896
rect 2490 56830 13642 56840
rect 2670 56715 13350 56747
rect 2670 56559 2682 56715
rect 2838 56559 3682 56715
rect 3838 56559 4182 56715
rect 4338 56559 5182 56715
rect 5338 56559 5682 56715
rect 5838 56559 6682 56715
rect 6838 56559 7182 56715
rect 7338 56559 8182 56715
rect 8338 56559 8682 56715
rect 8838 56559 9682 56715
rect 9838 56559 10182 56715
rect 10338 56559 11182 56715
rect 11338 56559 11682 56715
rect 11838 56559 12682 56715
rect 12838 56559 13182 56715
rect 13338 56559 13350 56715
rect 2670 56531 13350 56559
rect 2490 56438 13642 56448
rect 2490 56382 2500 56438
rect 2556 56418 2642 56438
rect 2698 56418 2784 56438
rect 2840 56418 2926 56438
rect 2982 56418 3068 56438
rect 3124 56418 3210 56438
rect 2574 56382 2642 56418
rect 2490 56366 2522 56382
rect 2574 56366 2646 56382
rect 2698 56366 2770 56418
rect 2840 56382 2894 56418
rect 2982 56382 3018 56418
rect 3124 56382 3142 56418
rect 2822 56366 2894 56382
rect 2946 56366 3018 56382
rect 3070 56366 3142 56382
rect 3194 56382 3210 56418
rect 3266 56418 3352 56438
rect 3408 56418 3494 56438
rect 3550 56418 3636 56438
rect 3692 56418 3778 56438
rect 3834 56418 3920 56438
rect 3976 56418 4062 56438
rect 3194 56366 3266 56382
rect 3318 56382 3352 56418
rect 3442 56382 3494 56418
rect 3566 56382 3636 56418
rect 3692 56382 3762 56418
rect 3834 56382 3886 56418
rect 3976 56382 4010 56418
rect 3318 56366 3390 56382
rect 3442 56366 3514 56382
rect 3566 56366 3638 56382
rect 3690 56366 3762 56382
rect 3814 56366 3886 56382
rect 3938 56366 4010 56382
rect 4118 56418 4204 56438
rect 4260 56418 4346 56438
rect 4402 56418 4488 56438
rect 4544 56418 4630 56438
rect 4686 56418 4772 56438
rect 4828 56418 4914 56438
rect 4970 56418 5056 56438
rect 4118 56382 4134 56418
rect 4062 56366 4134 56382
rect 4186 56382 4204 56418
rect 4310 56382 4346 56418
rect 4434 56382 4488 56418
rect 4186 56366 4258 56382
rect 4310 56366 4382 56382
rect 4434 56366 4506 56382
rect 4558 56366 4630 56418
rect 4686 56382 4754 56418
rect 4828 56382 4878 56418
rect 4970 56382 5002 56418
rect 4682 56366 4754 56382
rect 4806 56366 4878 56382
rect 4930 56366 5002 56382
rect 5054 56382 5056 56418
rect 5112 56418 5198 56438
rect 5254 56418 5340 56438
rect 5396 56418 5482 56438
rect 5538 56418 5624 56438
rect 5680 56418 5766 56438
rect 5822 56418 5908 56438
rect 5964 56418 6050 56438
rect 5112 56382 5126 56418
rect 5054 56366 5126 56382
rect 5178 56382 5198 56418
rect 5302 56382 5340 56418
rect 5426 56382 5482 56418
rect 5178 56366 5250 56382
rect 5302 56366 5374 56382
rect 5426 56366 5498 56382
rect 5550 56366 5622 56418
rect 5680 56382 5746 56418
rect 5822 56382 5870 56418
rect 5964 56382 5994 56418
rect 5674 56366 5746 56382
rect 5798 56366 5870 56382
rect 5922 56366 5994 56382
rect 6046 56382 6050 56418
rect 6106 56418 6192 56438
rect 6248 56418 6334 56438
rect 6390 56418 6476 56438
rect 6532 56418 6618 56438
rect 6674 56418 6760 56438
rect 6816 56418 6902 56438
rect 6958 56418 7044 56438
rect 6106 56382 6118 56418
rect 6046 56366 6118 56382
rect 6170 56382 6192 56418
rect 6294 56382 6334 56418
rect 6418 56382 6476 56418
rect 6170 56366 6242 56382
rect 6294 56366 6366 56382
rect 6418 56366 6490 56382
rect 6542 56366 6614 56418
rect 6674 56382 6738 56418
rect 6816 56382 6862 56418
rect 6958 56382 6986 56418
rect 6666 56366 6738 56382
rect 6790 56366 6862 56382
rect 6914 56366 6986 56382
rect 7038 56382 7044 56418
rect 7100 56418 7186 56438
rect 7242 56418 7328 56438
rect 7384 56418 7470 56438
rect 7526 56418 7612 56438
rect 7668 56418 7754 56438
rect 7810 56418 7896 56438
rect 7952 56418 8038 56438
rect 7100 56382 7110 56418
rect 7038 56366 7110 56382
rect 7162 56382 7186 56418
rect 7286 56382 7328 56418
rect 7410 56382 7470 56418
rect 7162 56366 7234 56382
rect 7286 56366 7358 56382
rect 7410 56366 7482 56382
rect 7534 56366 7606 56418
rect 7668 56382 7730 56418
rect 7810 56382 7854 56418
rect 7952 56382 7978 56418
rect 7658 56366 7730 56382
rect 7782 56366 7854 56382
rect 7906 56366 7978 56382
rect 8030 56382 8038 56418
rect 8094 56418 8180 56438
rect 8236 56418 8322 56438
rect 8378 56418 8464 56438
rect 8520 56418 8606 56438
rect 8662 56418 8748 56438
rect 8804 56418 8890 56438
rect 8946 56418 9032 56438
rect 8094 56382 8102 56418
rect 8030 56366 8102 56382
rect 8154 56382 8180 56418
rect 8278 56382 8322 56418
rect 8402 56382 8464 56418
rect 8154 56366 8226 56382
rect 8278 56366 8350 56382
rect 8402 56366 8474 56382
rect 8526 56366 8598 56418
rect 8662 56382 8722 56418
rect 8804 56382 8846 56418
rect 8946 56382 8970 56418
rect 8650 56366 8722 56382
rect 8774 56366 8846 56382
rect 8898 56366 8970 56382
rect 9022 56382 9032 56418
rect 9088 56418 9174 56438
rect 9230 56418 9316 56438
rect 9372 56418 9458 56438
rect 9514 56418 9600 56438
rect 9656 56418 9742 56438
rect 9798 56418 9884 56438
rect 9940 56418 10026 56438
rect 9088 56382 9094 56418
rect 9022 56366 9094 56382
rect 9146 56382 9174 56418
rect 9270 56382 9316 56418
rect 9394 56382 9458 56418
rect 9146 56366 9218 56382
rect 9270 56366 9342 56382
rect 9394 56366 9466 56382
rect 9518 56366 9590 56418
rect 9656 56382 9714 56418
rect 9798 56382 9838 56418
rect 9940 56382 9962 56418
rect 9642 56366 9714 56382
rect 9766 56366 9838 56382
rect 9890 56366 9962 56382
rect 10014 56382 10026 56418
rect 10082 56418 10168 56438
rect 10224 56418 10310 56438
rect 10366 56418 10452 56438
rect 10508 56418 10594 56438
rect 10650 56418 10736 56438
rect 10792 56418 10878 56438
rect 10934 56418 11020 56438
rect 10082 56382 10086 56418
rect 10014 56366 10086 56382
rect 10138 56382 10168 56418
rect 10262 56382 10310 56418
rect 10386 56382 10452 56418
rect 10138 56366 10210 56382
rect 10262 56366 10334 56382
rect 10386 56366 10458 56382
rect 10510 56366 10582 56418
rect 10650 56382 10706 56418
rect 10792 56382 10830 56418
rect 10934 56382 10954 56418
rect 10634 56366 10706 56382
rect 10758 56366 10830 56382
rect 10882 56366 10954 56382
rect 11006 56382 11020 56418
rect 11076 56418 11162 56438
rect 11218 56418 11304 56438
rect 11360 56418 11446 56438
rect 11502 56418 11588 56438
rect 11644 56418 11730 56438
rect 11786 56418 11872 56438
rect 11928 56418 12014 56438
rect 11076 56382 11078 56418
rect 11006 56366 11078 56382
rect 11130 56382 11162 56418
rect 11254 56382 11304 56418
rect 11378 56382 11446 56418
rect 11130 56366 11202 56382
rect 11254 56366 11326 56382
rect 11378 56366 11450 56382
rect 11502 56366 11574 56418
rect 11644 56382 11698 56418
rect 11786 56382 11822 56418
rect 11928 56382 11946 56418
rect 11626 56366 11698 56382
rect 11750 56366 11822 56382
rect 11874 56366 11946 56382
rect 11998 56382 12014 56418
rect 12070 56418 12156 56438
rect 12212 56418 12298 56438
rect 12354 56418 12440 56438
rect 12496 56418 12582 56438
rect 12638 56418 12724 56438
rect 12780 56418 12866 56438
rect 11998 56366 12070 56382
rect 12122 56382 12156 56418
rect 12246 56382 12298 56418
rect 12370 56382 12440 56418
rect 12496 56382 12566 56418
rect 12638 56382 12690 56418
rect 12780 56382 12814 56418
rect 12122 56366 12194 56382
rect 12246 56366 12318 56382
rect 12370 56366 12442 56382
rect 12494 56366 12566 56382
rect 12618 56366 12690 56382
rect 12742 56366 12814 56382
rect 12922 56418 13008 56438
rect 13064 56418 13150 56438
rect 13206 56418 13292 56438
rect 13348 56418 13434 56438
rect 13490 56418 13576 56438
rect 12922 56382 12938 56418
rect 12866 56366 12938 56382
rect 12990 56382 13008 56418
rect 13114 56382 13150 56418
rect 13238 56382 13292 56418
rect 12990 56366 13062 56382
rect 13114 56366 13186 56382
rect 13238 56366 13310 56382
rect 13362 56366 13434 56418
rect 13490 56382 13558 56418
rect 13632 56382 13642 56438
rect 13486 56366 13558 56382
rect 13610 56366 13642 56382
rect 2490 56296 13642 56366
rect 2490 56240 2500 56296
rect 2556 56294 2642 56296
rect 2698 56294 2784 56296
rect 2840 56294 2926 56296
rect 2982 56294 3068 56296
rect 3124 56294 3210 56296
rect 2574 56242 2642 56294
rect 2698 56242 2770 56294
rect 2840 56242 2894 56294
rect 2982 56242 3018 56294
rect 3124 56242 3142 56294
rect 3194 56242 3210 56294
rect 2556 56240 2642 56242
rect 2698 56240 2784 56242
rect 2840 56240 2926 56242
rect 2982 56240 3068 56242
rect 3124 56240 3210 56242
rect 3266 56294 3352 56296
rect 3408 56294 3494 56296
rect 3550 56294 3636 56296
rect 3692 56294 3778 56296
rect 3834 56294 3920 56296
rect 3976 56294 4062 56296
rect 3318 56242 3352 56294
rect 3442 56242 3494 56294
rect 3566 56242 3636 56294
rect 3692 56242 3762 56294
rect 3834 56242 3886 56294
rect 3976 56242 4010 56294
rect 3266 56240 3352 56242
rect 3408 56240 3494 56242
rect 3550 56240 3636 56242
rect 3692 56240 3778 56242
rect 3834 56240 3920 56242
rect 3976 56240 4062 56242
rect 4118 56294 4204 56296
rect 4260 56294 4346 56296
rect 4402 56294 4488 56296
rect 4544 56294 4630 56296
rect 4686 56294 4772 56296
rect 4828 56294 4914 56296
rect 4970 56294 5056 56296
rect 4118 56242 4134 56294
rect 4186 56242 4204 56294
rect 4310 56242 4346 56294
rect 4434 56242 4488 56294
rect 4558 56242 4630 56294
rect 4686 56242 4754 56294
rect 4828 56242 4878 56294
rect 4970 56242 5002 56294
rect 5054 56242 5056 56294
rect 4118 56240 4204 56242
rect 4260 56240 4346 56242
rect 4402 56240 4488 56242
rect 4544 56240 4630 56242
rect 4686 56240 4772 56242
rect 4828 56240 4914 56242
rect 4970 56240 5056 56242
rect 5112 56294 5198 56296
rect 5254 56294 5340 56296
rect 5396 56294 5482 56296
rect 5538 56294 5624 56296
rect 5680 56294 5766 56296
rect 5822 56294 5908 56296
rect 5964 56294 6050 56296
rect 5112 56242 5126 56294
rect 5178 56242 5198 56294
rect 5302 56242 5340 56294
rect 5426 56242 5482 56294
rect 5550 56242 5622 56294
rect 5680 56242 5746 56294
rect 5822 56242 5870 56294
rect 5964 56242 5994 56294
rect 6046 56242 6050 56294
rect 5112 56240 5198 56242
rect 5254 56240 5340 56242
rect 5396 56240 5482 56242
rect 5538 56240 5624 56242
rect 5680 56240 5766 56242
rect 5822 56240 5908 56242
rect 5964 56240 6050 56242
rect 6106 56294 6192 56296
rect 6248 56294 6334 56296
rect 6390 56294 6476 56296
rect 6532 56294 6618 56296
rect 6674 56294 6760 56296
rect 6816 56294 6902 56296
rect 6958 56294 7044 56296
rect 6106 56242 6118 56294
rect 6170 56242 6192 56294
rect 6294 56242 6334 56294
rect 6418 56242 6476 56294
rect 6542 56242 6614 56294
rect 6674 56242 6738 56294
rect 6816 56242 6862 56294
rect 6958 56242 6986 56294
rect 7038 56242 7044 56294
rect 6106 56240 6192 56242
rect 6248 56240 6334 56242
rect 6390 56240 6476 56242
rect 6532 56240 6618 56242
rect 6674 56240 6760 56242
rect 6816 56240 6902 56242
rect 6958 56240 7044 56242
rect 7100 56294 7186 56296
rect 7242 56294 7328 56296
rect 7384 56294 7470 56296
rect 7526 56294 7612 56296
rect 7668 56294 7754 56296
rect 7810 56294 7896 56296
rect 7952 56294 8038 56296
rect 7100 56242 7110 56294
rect 7162 56242 7186 56294
rect 7286 56242 7328 56294
rect 7410 56242 7470 56294
rect 7534 56242 7606 56294
rect 7668 56242 7730 56294
rect 7810 56242 7854 56294
rect 7952 56242 7978 56294
rect 8030 56242 8038 56294
rect 7100 56240 7186 56242
rect 7242 56240 7328 56242
rect 7384 56240 7470 56242
rect 7526 56240 7612 56242
rect 7668 56240 7754 56242
rect 7810 56240 7896 56242
rect 7952 56240 8038 56242
rect 8094 56294 8180 56296
rect 8236 56294 8322 56296
rect 8378 56294 8464 56296
rect 8520 56294 8606 56296
rect 8662 56294 8748 56296
rect 8804 56294 8890 56296
rect 8946 56294 9032 56296
rect 8094 56242 8102 56294
rect 8154 56242 8180 56294
rect 8278 56242 8322 56294
rect 8402 56242 8464 56294
rect 8526 56242 8598 56294
rect 8662 56242 8722 56294
rect 8804 56242 8846 56294
rect 8946 56242 8970 56294
rect 9022 56242 9032 56294
rect 8094 56240 8180 56242
rect 8236 56240 8322 56242
rect 8378 56240 8464 56242
rect 8520 56240 8606 56242
rect 8662 56240 8748 56242
rect 8804 56240 8890 56242
rect 8946 56240 9032 56242
rect 9088 56294 9174 56296
rect 9230 56294 9316 56296
rect 9372 56294 9458 56296
rect 9514 56294 9600 56296
rect 9656 56294 9742 56296
rect 9798 56294 9884 56296
rect 9940 56294 10026 56296
rect 9088 56242 9094 56294
rect 9146 56242 9174 56294
rect 9270 56242 9316 56294
rect 9394 56242 9458 56294
rect 9518 56242 9590 56294
rect 9656 56242 9714 56294
rect 9798 56242 9838 56294
rect 9940 56242 9962 56294
rect 10014 56242 10026 56294
rect 9088 56240 9174 56242
rect 9230 56240 9316 56242
rect 9372 56240 9458 56242
rect 9514 56240 9600 56242
rect 9656 56240 9742 56242
rect 9798 56240 9884 56242
rect 9940 56240 10026 56242
rect 10082 56294 10168 56296
rect 10224 56294 10310 56296
rect 10366 56294 10452 56296
rect 10508 56294 10594 56296
rect 10650 56294 10736 56296
rect 10792 56294 10878 56296
rect 10934 56294 11020 56296
rect 10082 56242 10086 56294
rect 10138 56242 10168 56294
rect 10262 56242 10310 56294
rect 10386 56242 10452 56294
rect 10510 56242 10582 56294
rect 10650 56242 10706 56294
rect 10792 56242 10830 56294
rect 10934 56242 10954 56294
rect 11006 56242 11020 56294
rect 10082 56240 10168 56242
rect 10224 56240 10310 56242
rect 10366 56240 10452 56242
rect 10508 56240 10594 56242
rect 10650 56240 10736 56242
rect 10792 56240 10878 56242
rect 10934 56240 11020 56242
rect 11076 56294 11162 56296
rect 11218 56294 11304 56296
rect 11360 56294 11446 56296
rect 11502 56294 11588 56296
rect 11644 56294 11730 56296
rect 11786 56294 11872 56296
rect 11928 56294 12014 56296
rect 11076 56242 11078 56294
rect 11130 56242 11162 56294
rect 11254 56242 11304 56294
rect 11378 56242 11446 56294
rect 11502 56242 11574 56294
rect 11644 56242 11698 56294
rect 11786 56242 11822 56294
rect 11928 56242 11946 56294
rect 11998 56242 12014 56294
rect 11076 56240 11162 56242
rect 11218 56240 11304 56242
rect 11360 56240 11446 56242
rect 11502 56240 11588 56242
rect 11644 56240 11730 56242
rect 11786 56240 11872 56242
rect 11928 56240 12014 56242
rect 12070 56294 12156 56296
rect 12212 56294 12298 56296
rect 12354 56294 12440 56296
rect 12496 56294 12582 56296
rect 12638 56294 12724 56296
rect 12780 56294 12866 56296
rect 12122 56242 12156 56294
rect 12246 56242 12298 56294
rect 12370 56242 12440 56294
rect 12496 56242 12566 56294
rect 12638 56242 12690 56294
rect 12780 56242 12814 56294
rect 12070 56240 12156 56242
rect 12212 56240 12298 56242
rect 12354 56240 12440 56242
rect 12496 56240 12582 56242
rect 12638 56240 12724 56242
rect 12780 56240 12866 56242
rect 12922 56294 13008 56296
rect 13064 56294 13150 56296
rect 13206 56294 13292 56296
rect 13348 56294 13434 56296
rect 13490 56294 13576 56296
rect 12922 56242 12938 56294
rect 12990 56242 13008 56294
rect 13114 56242 13150 56294
rect 13238 56242 13292 56294
rect 13362 56242 13434 56294
rect 13490 56242 13558 56294
rect 12922 56240 13008 56242
rect 13064 56240 13150 56242
rect 13206 56240 13292 56242
rect 13348 56240 13434 56242
rect 13490 56240 13576 56242
rect 13632 56240 13642 56296
rect 2490 56170 13642 56240
rect 2490 56154 2522 56170
rect 2574 56154 2646 56170
rect 2490 56098 2500 56154
rect 2574 56118 2642 56154
rect 2698 56118 2770 56170
rect 2822 56154 2894 56170
rect 2946 56154 3018 56170
rect 3070 56154 3142 56170
rect 2840 56118 2894 56154
rect 2982 56118 3018 56154
rect 3124 56118 3142 56154
rect 3194 56154 3266 56170
rect 3194 56118 3210 56154
rect 2556 56098 2642 56118
rect 2698 56098 2784 56118
rect 2840 56098 2926 56118
rect 2982 56098 3068 56118
rect 3124 56098 3210 56118
rect 3318 56154 3390 56170
rect 3442 56154 3514 56170
rect 3566 56154 3638 56170
rect 3690 56154 3762 56170
rect 3814 56154 3886 56170
rect 3938 56154 4010 56170
rect 3318 56118 3352 56154
rect 3442 56118 3494 56154
rect 3566 56118 3636 56154
rect 3692 56118 3762 56154
rect 3834 56118 3886 56154
rect 3976 56118 4010 56154
rect 4062 56154 4134 56170
rect 3266 56098 3352 56118
rect 3408 56098 3494 56118
rect 3550 56098 3636 56118
rect 3692 56098 3778 56118
rect 3834 56098 3920 56118
rect 3976 56098 4062 56118
rect 4118 56118 4134 56154
rect 4186 56154 4258 56170
rect 4310 56154 4382 56170
rect 4434 56154 4506 56170
rect 4186 56118 4204 56154
rect 4310 56118 4346 56154
rect 4434 56118 4488 56154
rect 4558 56118 4630 56170
rect 4682 56154 4754 56170
rect 4806 56154 4878 56170
rect 4930 56154 5002 56170
rect 4686 56118 4754 56154
rect 4828 56118 4878 56154
rect 4970 56118 5002 56154
rect 5054 56154 5126 56170
rect 5054 56118 5056 56154
rect 4118 56098 4204 56118
rect 4260 56098 4346 56118
rect 4402 56098 4488 56118
rect 4544 56098 4630 56118
rect 4686 56098 4772 56118
rect 4828 56098 4914 56118
rect 4970 56098 5056 56118
rect 5112 56118 5126 56154
rect 5178 56154 5250 56170
rect 5302 56154 5374 56170
rect 5426 56154 5498 56170
rect 5178 56118 5198 56154
rect 5302 56118 5340 56154
rect 5426 56118 5482 56154
rect 5550 56118 5622 56170
rect 5674 56154 5746 56170
rect 5798 56154 5870 56170
rect 5922 56154 5994 56170
rect 5680 56118 5746 56154
rect 5822 56118 5870 56154
rect 5964 56118 5994 56154
rect 6046 56154 6118 56170
rect 6046 56118 6050 56154
rect 5112 56098 5198 56118
rect 5254 56098 5340 56118
rect 5396 56098 5482 56118
rect 5538 56098 5624 56118
rect 5680 56098 5766 56118
rect 5822 56098 5908 56118
rect 5964 56098 6050 56118
rect 6106 56118 6118 56154
rect 6170 56154 6242 56170
rect 6294 56154 6366 56170
rect 6418 56154 6490 56170
rect 6170 56118 6192 56154
rect 6294 56118 6334 56154
rect 6418 56118 6476 56154
rect 6542 56118 6614 56170
rect 6666 56154 6738 56170
rect 6790 56154 6862 56170
rect 6914 56154 6986 56170
rect 6674 56118 6738 56154
rect 6816 56118 6862 56154
rect 6958 56118 6986 56154
rect 7038 56154 7110 56170
rect 7038 56118 7044 56154
rect 6106 56098 6192 56118
rect 6248 56098 6334 56118
rect 6390 56098 6476 56118
rect 6532 56098 6618 56118
rect 6674 56098 6760 56118
rect 6816 56098 6902 56118
rect 6958 56098 7044 56118
rect 7100 56118 7110 56154
rect 7162 56154 7234 56170
rect 7286 56154 7358 56170
rect 7410 56154 7482 56170
rect 7162 56118 7186 56154
rect 7286 56118 7328 56154
rect 7410 56118 7470 56154
rect 7534 56118 7606 56170
rect 7658 56154 7730 56170
rect 7782 56154 7854 56170
rect 7906 56154 7978 56170
rect 7668 56118 7730 56154
rect 7810 56118 7854 56154
rect 7952 56118 7978 56154
rect 8030 56154 8102 56170
rect 8030 56118 8038 56154
rect 7100 56098 7186 56118
rect 7242 56098 7328 56118
rect 7384 56098 7470 56118
rect 7526 56098 7612 56118
rect 7668 56098 7754 56118
rect 7810 56098 7896 56118
rect 7952 56098 8038 56118
rect 8094 56118 8102 56154
rect 8154 56154 8226 56170
rect 8278 56154 8350 56170
rect 8402 56154 8474 56170
rect 8154 56118 8180 56154
rect 8278 56118 8322 56154
rect 8402 56118 8464 56154
rect 8526 56118 8598 56170
rect 8650 56154 8722 56170
rect 8774 56154 8846 56170
rect 8898 56154 8970 56170
rect 8662 56118 8722 56154
rect 8804 56118 8846 56154
rect 8946 56118 8970 56154
rect 9022 56154 9094 56170
rect 9022 56118 9032 56154
rect 8094 56098 8180 56118
rect 8236 56098 8322 56118
rect 8378 56098 8464 56118
rect 8520 56098 8606 56118
rect 8662 56098 8748 56118
rect 8804 56098 8890 56118
rect 8946 56098 9032 56118
rect 9088 56118 9094 56154
rect 9146 56154 9218 56170
rect 9270 56154 9342 56170
rect 9394 56154 9466 56170
rect 9146 56118 9174 56154
rect 9270 56118 9316 56154
rect 9394 56118 9458 56154
rect 9518 56118 9590 56170
rect 9642 56154 9714 56170
rect 9766 56154 9838 56170
rect 9890 56154 9962 56170
rect 9656 56118 9714 56154
rect 9798 56118 9838 56154
rect 9940 56118 9962 56154
rect 10014 56154 10086 56170
rect 10014 56118 10026 56154
rect 9088 56098 9174 56118
rect 9230 56098 9316 56118
rect 9372 56098 9458 56118
rect 9514 56098 9600 56118
rect 9656 56098 9742 56118
rect 9798 56098 9884 56118
rect 9940 56098 10026 56118
rect 10082 56118 10086 56154
rect 10138 56154 10210 56170
rect 10262 56154 10334 56170
rect 10386 56154 10458 56170
rect 10138 56118 10168 56154
rect 10262 56118 10310 56154
rect 10386 56118 10452 56154
rect 10510 56118 10582 56170
rect 10634 56154 10706 56170
rect 10758 56154 10830 56170
rect 10882 56154 10954 56170
rect 10650 56118 10706 56154
rect 10792 56118 10830 56154
rect 10934 56118 10954 56154
rect 11006 56154 11078 56170
rect 11006 56118 11020 56154
rect 10082 56098 10168 56118
rect 10224 56098 10310 56118
rect 10366 56098 10452 56118
rect 10508 56098 10594 56118
rect 10650 56098 10736 56118
rect 10792 56098 10878 56118
rect 10934 56098 11020 56118
rect 11076 56118 11078 56154
rect 11130 56154 11202 56170
rect 11254 56154 11326 56170
rect 11378 56154 11450 56170
rect 11130 56118 11162 56154
rect 11254 56118 11304 56154
rect 11378 56118 11446 56154
rect 11502 56118 11574 56170
rect 11626 56154 11698 56170
rect 11750 56154 11822 56170
rect 11874 56154 11946 56170
rect 11644 56118 11698 56154
rect 11786 56118 11822 56154
rect 11928 56118 11946 56154
rect 11998 56154 12070 56170
rect 11998 56118 12014 56154
rect 11076 56098 11162 56118
rect 11218 56098 11304 56118
rect 11360 56098 11446 56118
rect 11502 56098 11588 56118
rect 11644 56098 11730 56118
rect 11786 56098 11872 56118
rect 11928 56098 12014 56118
rect 12122 56154 12194 56170
rect 12246 56154 12318 56170
rect 12370 56154 12442 56170
rect 12494 56154 12566 56170
rect 12618 56154 12690 56170
rect 12742 56154 12814 56170
rect 12122 56118 12156 56154
rect 12246 56118 12298 56154
rect 12370 56118 12440 56154
rect 12496 56118 12566 56154
rect 12638 56118 12690 56154
rect 12780 56118 12814 56154
rect 12866 56154 12938 56170
rect 12070 56098 12156 56118
rect 12212 56098 12298 56118
rect 12354 56098 12440 56118
rect 12496 56098 12582 56118
rect 12638 56098 12724 56118
rect 12780 56098 12866 56118
rect 12922 56118 12938 56154
rect 12990 56154 13062 56170
rect 13114 56154 13186 56170
rect 13238 56154 13310 56170
rect 12990 56118 13008 56154
rect 13114 56118 13150 56154
rect 13238 56118 13292 56154
rect 13362 56118 13434 56170
rect 13486 56154 13558 56170
rect 13610 56154 13642 56170
rect 13490 56118 13558 56154
rect 12922 56098 13008 56118
rect 13064 56098 13150 56118
rect 13206 56098 13292 56118
rect 13348 56098 13434 56118
rect 13490 56098 13576 56118
rect 13632 56098 13642 56154
rect 2490 56088 13642 56098
rect 3500 55849 13350 55925
rect 3500 55837 4096 55849
rect 3500 55785 3512 55837
rect 4084 55785 4096 55837
rect 3500 55773 4096 55785
rect 8030 55829 8106 55849
rect 4938 55758 5014 55770
rect 4938 55751 4950 55758
rect 5002 55751 5014 55758
rect 4750 55741 4826 55751
rect 2309 55711 2385 55741
rect 2309 55555 2321 55711
rect 2373 55555 2385 55711
rect 2309 54460 2385 55555
rect 4750 55685 4760 55741
rect 4816 55685 4826 55741
rect 4750 55599 4762 55685
rect 4814 55599 4826 55685
rect 4750 55543 4760 55599
rect 4816 55543 4826 55599
rect 2593 55463 4238 55475
rect 2593 55411 2605 55463
rect 2761 55411 4238 55463
rect 2593 55399 4238 55411
rect 4162 54692 4238 55399
rect 4750 55457 4762 55543
rect 4814 55457 4826 55543
rect 4750 55401 4760 55457
rect 4816 55401 4826 55457
rect 4750 55315 4762 55401
rect 4814 55315 4826 55401
rect 4750 55259 4760 55315
rect 4816 55259 4826 55315
rect 4750 55173 4762 55259
rect 4814 55173 4826 55259
rect 4750 55117 4760 55173
rect 4816 55117 4826 55173
rect 4750 55031 4762 55117
rect 4814 55031 4826 55117
rect 4750 54975 4760 55031
rect 4816 54975 4826 55031
rect 4750 54889 4762 54975
rect 4814 54889 4826 54975
rect 4938 55695 4948 55751
rect 5004 55695 5014 55751
rect 4938 55609 4950 55695
rect 5002 55609 5014 55695
rect 4938 55553 4948 55609
rect 5004 55553 5014 55609
rect 4938 55467 4950 55553
rect 5002 55467 5014 55553
rect 4938 55411 4948 55467
rect 5004 55411 5014 55467
rect 4938 55325 4950 55411
rect 5002 55325 5014 55411
rect 4938 55269 4948 55325
rect 5004 55269 5014 55325
rect 4938 55183 4950 55269
rect 5002 55183 5014 55269
rect 4938 55127 4948 55183
rect 5004 55127 5014 55183
rect 4938 55041 4950 55127
rect 5002 55041 5014 55127
rect 4938 54985 4948 55041
rect 5004 54985 5014 55041
rect 4938 54978 4950 54985
rect 5002 54978 5014 54985
rect 4938 54966 5014 54978
rect 5426 55767 5502 55779
rect 5426 55760 5438 55767
rect 5490 55760 5502 55767
rect 5426 55704 5436 55760
rect 5492 55704 5502 55760
rect 5426 55618 5438 55704
rect 5490 55618 5502 55704
rect 5426 55562 5436 55618
rect 5492 55562 5502 55618
rect 5426 55476 5438 55562
rect 5490 55476 5502 55562
rect 5426 55420 5436 55476
rect 5492 55420 5502 55476
rect 5426 55334 5438 55420
rect 5490 55334 5502 55420
rect 5426 55278 5436 55334
rect 5492 55278 5502 55334
rect 5426 55192 5438 55278
rect 5490 55192 5502 55278
rect 5426 55136 5436 55192
rect 5492 55136 5502 55192
rect 5426 55050 5438 55136
rect 5490 55050 5502 55136
rect 5426 54994 5436 55050
rect 5492 54994 5502 55050
rect 5426 54987 5438 54994
rect 5490 54987 5502 54994
rect 5426 54975 5502 54987
rect 5914 55767 5990 55779
rect 5914 55760 5926 55767
rect 5978 55760 5990 55767
rect 5914 55704 5924 55760
rect 5980 55704 5990 55760
rect 6278 55767 6354 55779
rect 6278 55760 6290 55767
rect 6342 55760 6354 55767
rect 5914 55618 5926 55704
rect 5978 55618 5990 55704
rect 5914 55562 5924 55618
rect 5980 55562 5990 55618
rect 5914 55476 5926 55562
rect 5978 55476 5990 55562
rect 5914 55420 5924 55476
rect 5980 55420 5990 55476
rect 5914 55334 5926 55420
rect 5978 55334 5990 55420
rect 5914 55278 5924 55334
rect 5980 55278 5990 55334
rect 5914 55192 5926 55278
rect 5978 55192 5990 55278
rect 5914 55136 5924 55192
rect 5980 55136 5990 55192
rect 5914 55050 5926 55136
rect 5978 55050 5990 55136
rect 5914 54994 5924 55050
rect 5980 54994 5990 55050
rect 5914 54987 5926 54994
rect 5978 54987 5990 54994
rect 5914 54975 5990 54987
rect 6096 55741 6172 55751
rect 6096 55685 6106 55741
rect 6162 55685 6172 55741
rect 6096 55599 6108 55685
rect 6160 55599 6172 55685
rect 6096 55543 6106 55599
rect 6162 55543 6172 55599
rect 6096 55457 6108 55543
rect 6160 55457 6172 55543
rect 6096 55401 6106 55457
rect 6162 55401 6172 55457
rect 6096 55315 6108 55401
rect 6160 55315 6172 55401
rect 6096 55259 6106 55315
rect 6162 55259 6172 55315
rect 6096 55173 6108 55259
rect 6160 55173 6172 55259
rect 6096 55117 6106 55173
rect 6162 55117 6172 55173
rect 6096 55031 6108 55117
rect 6160 55031 6172 55117
rect 6096 54975 6106 55031
rect 6162 54975 6172 55031
rect 6278 55704 6288 55760
rect 6344 55704 6354 55760
rect 6278 55618 6290 55704
rect 6342 55618 6354 55704
rect 6278 55562 6288 55618
rect 6344 55562 6354 55618
rect 6278 55476 6290 55562
rect 6342 55476 6354 55562
rect 6278 55420 6288 55476
rect 6344 55420 6354 55476
rect 6278 55334 6290 55420
rect 6342 55334 6354 55420
rect 6278 55278 6288 55334
rect 6344 55278 6354 55334
rect 6278 55192 6290 55278
rect 6342 55192 6354 55278
rect 6278 55136 6288 55192
rect 6344 55136 6354 55192
rect 6278 55050 6290 55136
rect 6342 55050 6354 55136
rect 6278 54994 6288 55050
rect 6344 54994 6354 55050
rect 6278 54987 6290 54994
rect 6342 54987 6354 54994
rect 6278 54975 6354 54987
rect 6766 55767 6842 55779
rect 6766 55760 6778 55767
rect 6830 55760 6842 55767
rect 6766 55704 6776 55760
rect 6832 55704 6842 55760
rect 6766 55618 6778 55704
rect 6830 55618 6842 55704
rect 6766 55562 6776 55618
rect 6832 55562 6842 55618
rect 6766 55476 6778 55562
rect 6830 55476 6842 55562
rect 6766 55420 6776 55476
rect 6832 55420 6842 55476
rect 6766 55334 6778 55420
rect 6830 55334 6842 55420
rect 6766 55278 6776 55334
rect 6832 55278 6842 55334
rect 6766 55192 6778 55278
rect 6830 55192 6842 55278
rect 6766 55136 6776 55192
rect 6832 55136 6842 55192
rect 6766 55050 6778 55136
rect 6830 55050 6842 55136
rect 6766 54994 6776 55050
rect 6832 54994 6842 55050
rect 6766 54987 6778 54994
rect 6830 54987 6842 54994
rect 6766 54975 6842 54987
rect 7254 55767 7330 55779
rect 7254 55760 7266 55767
rect 7318 55760 7330 55767
rect 7254 55704 7264 55760
rect 7320 55704 7330 55760
rect 7254 55618 7266 55704
rect 7318 55618 7330 55704
rect 7254 55562 7264 55618
rect 7320 55562 7330 55618
rect 7254 55476 7266 55562
rect 7318 55476 7330 55562
rect 7254 55420 7264 55476
rect 7320 55420 7330 55476
rect 7254 55334 7266 55420
rect 7318 55334 7330 55420
rect 7254 55278 7264 55334
rect 7320 55278 7330 55334
rect 7254 55192 7266 55278
rect 7318 55192 7330 55278
rect 7254 55136 7264 55192
rect 7320 55136 7330 55192
rect 7254 55050 7266 55136
rect 7318 55050 7330 55136
rect 7254 54994 7264 55050
rect 7320 54994 7330 55050
rect 7254 54987 7266 54994
rect 7318 54987 7330 54994
rect 7254 54975 7330 54987
rect 7442 55741 7518 55751
rect 7442 55685 7452 55741
rect 7508 55685 7518 55741
rect 7442 55599 7454 55685
rect 7506 55599 7518 55685
rect 7442 55543 7452 55599
rect 7508 55543 7518 55599
rect 7442 55457 7454 55543
rect 7506 55457 7518 55543
rect 7442 55401 7452 55457
rect 7508 55401 7518 55457
rect 7442 55315 7454 55401
rect 7506 55315 7518 55401
rect 7442 55259 7452 55315
rect 7508 55259 7518 55315
rect 7442 55173 7454 55259
rect 7506 55173 7518 55259
rect 7442 55117 7452 55173
rect 7508 55117 7518 55173
rect 7442 55031 7454 55117
rect 7506 55031 7518 55117
rect 7442 54975 7452 55031
rect 7508 54975 7518 55031
rect 4750 54833 4760 54889
rect 4816 54833 4826 54889
rect 4750 54823 4826 54833
rect 6096 54889 6108 54975
rect 6160 54889 6172 54975
rect 6096 54833 6106 54889
rect 6162 54833 6172 54889
rect 6096 54823 6172 54833
rect 7442 54889 7454 54975
rect 7506 54889 7518 54975
rect 7442 54833 7452 54889
rect 7508 54833 7518 54889
rect 7442 54823 7518 54833
rect 8030 54841 8042 55829
rect 8094 54841 8106 55829
rect 8030 54829 8106 54841
rect 8499 55829 8575 55849
rect 8499 54841 8511 55829
rect 8563 54841 8575 55829
rect 8499 54829 8575 54841
rect 8714 55829 8790 55849
rect 8714 54841 8726 55829
rect 8778 54841 8790 55829
rect 8714 54829 8790 54841
rect 8937 55829 9013 55849
rect 8937 54841 8949 55829
rect 9001 54841 9013 55829
rect 8937 54829 9013 54841
rect 9406 55829 9482 55849
rect 9406 54841 9418 55829
rect 9470 54841 9482 55829
rect 10182 55767 10258 55779
rect 10182 55760 10194 55767
rect 10246 55760 10258 55767
rect 9406 54829 9482 54841
rect 9994 55741 10070 55751
rect 9994 55685 10004 55741
rect 10060 55685 10070 55741
rect 9994 55599 10006 55685
rect 10058 55599 10070 55685
rect 9994 55543 10004 55599
rect 10060 55543 10070 55599
rect 9994 55457 10006 55543
rect 10058 55457 10070 55543
rect 9994 55401 10004 55457
rect 10060 55401 10070 55457
rect 9994 55315 10006 55401
rect 10058 55315 10070 55401
rect 9994 55259 10004 55315
rect 10060 55259 10070 55315
rect 9994 55173 10006 55259
rect 10058 55173 10070 55259
rect 9994 55117 10004 55173
rect 10060 55117 10070 55173
rect 9994 55031 10006 55117
rect 10058 55031 10070 55117
rect 9994 54975 10004 55031
rect 10060 54975 10070 55031
rect 10182 55704 10192 55760
rect 10248 55704 10258 55760
rect 10182 55618 10194 55704
rect 10246 55618 10258 55704
rect 10182 55562 10192 55618
rect 10248 55562 10258 55618
rect 10182 55476 10194 55562
rect 10246 55476 10258 55562
rect 10182 55420 10192 55476
rect 10248 55420 10258 55476
rect 10182 55334 10194 55420
rect 10246 55334 10258 55420
rect 10182 55278 10192 55334
rect 10248 55278 10258 55334
rect 10182 55192 10194 55278
rect 10246 55192 10258 55278
rect 10182 55136 10192 55192
rect 10248 55136 10258 55192
rect 10182 55050 10194 55136
rect 10246 55050 10258 55136
rect 10182 54994 10192 55050
rect 10248 54994 10258 55050
rect 10182 54987 10194 54994
rect 10246 54987 10258 54994
rect 10182 54975 10258 54987
rect 10670 55767 10746 55779
rect 10670 55760 10682 55767
rect 10734 55760 10746 55767
rect 10670 55704 10680 55760
rect 10736 55704 10746 55760
rect 10670 55618 10682 55704
rect 10734 55618 10746 55704
rect 10670 55562 10680 55618
rect 10736 55562 10746 55618
rect 10670 55476 10682 55562
rect 10734 55476 10746 55562
rect 10670 55420 10680 55476
rect 10736 55420 10746 55476
rect 10670 55334 10682 55420
rect 10734 55334 10746 55420
rect 10670 55278 10680 55334
rect 10736 55278 10746 55334
rect 10670 55192 10682 55278
rect 10734 55192 10746 55278
rect 10670 55136 10680 55192
rect 10736 55136 10746 55192
rect 10670 55050 10682 55136
rect 10734 55050 10746 55136
rect 10670 54994 10680 55050
rect 10736 54994 10746 55050
rect 10670 54987 10682 54994
rect 10734 54987 10746 54994
rect 10670 54975 10746 54987
rect 11158 55767 11234 55779
rect 11158 55760 11170 55767
rect 11222 55760 11234 55767
rect 11158 55704 11168 55760
rect 11224 55704 11234 55760
rect 11522 55767 11598 55779
rect 11522 55760 11534 55767
rect 11586 55760 11598 55767
rect 11158 55618 11170 55704
rect 11222 55618 11234 55704
rect 11158 55562 11168 55618
rect 11224 55562 11234 55618
rect 11158 55476 11170 55562
rect 11222 55476 11234 55562
rect 11158 55420 11168 55476
rect 11224 55420 11234 55476
rect 11158 55334 11170 55420
rect 11222 55334 11234 55420
rect 11158 55278 11168 55334
rect 11224 55278 11234 55334
rect 11158 55192 11170 55278
rect 11222 55192 11234 55278
rect 11158 55136 11168 55192
rect 11224 55136 11234 55192
rect 11158 55050 11170 55136
rect 11222 55050 11234 55136
rect 11158 54994 11168 55050
rect 11224 54994 11234 55050
rect 11158 54987 11170 54994
rect 11222 54987 11234 54994
rect 11158 54975 11234 54987
rect 11340 55741 11416 55751
rect 11340 55685 11350 55741
rect 11406 55685 11416 55741
rect 11340 55599 11352 55685
rect 11404 55599 11416 55685
rect 11340 55543 11350 55599
rect 11406 55543 11416 55599
rect 11340 55457 11352 55543
rect 11404 55457 11416 55543
rect 11340 55401 11350 55457
rect 11406 55401 11416 55457
rect 11340 55315 11352 55401
rect 11404 55315 11416 55401
rect 11340 55259 11350 55315
rect 11406 55259 11416 55315
rect 11340 55173 11352 55259
rect 11404 55173 11416 55259
rect 11340 55117 11350 55173
rect 11406 55117 11416 55173
rect 11340 55031 11352 55117
rect 11404 55031 11416 55117
rect 11340 54975 11350 55031
rect 11406 54975 11416 55031
rect 11522 55704 11532 55760
rect 11588 55704 11598 55760
rect 11522 55618 11534 55704
rect 11586 55618 11598 55704
rect 11522 55562 11532 55618
rect 11588 55562 11598 55618
rect 11522 55476 11534 55562
rect 11586 55476 11598 55562
rect 11522 55420 11532 55476
rect 11588 55420 11598 55476
rect 11522 55334 11534 55420
rect 11586 55334 11598 55420
rect 11522 55278 11532 55334
rect 11588 55278 11598 55334
rect 11522 55192 11534 55278
rect 11586 55192 11598 55278
rect 11522 55136 11532 55192
rect 11588 55136 11598 55192
rect 11522 55050 11534 55136
rect 11586 55050 11598 55136
rect 11522 54994 11532 55050
rect 11588 54994 11598 55050
rect 11522 54987 11534 54994
rect 11586 54987 11598 54994
rect 11522 54975 11598 54987
rect 12010 55767 12086 55779
rect 12010 55760 12022 55767
rect 12074 55760 12086 55767
rect 12010 55704 12020 55760
rect 12076 55704 12086 55760
rect 12010 55618 12022 55704
rect 12074 55618 12086 55704
rect 12010 55562 12020 55618
rect 12076 55562 12086 55618
rect 12010 55476 12022 55562
rect 12074 55476 12086 55562
rect 12010 55420 12020 55476
rect 12076 55420 12086 55476
rect 12010 55334 12022 55420
rect 12074 55334 12086 55420
rect 12010 55278 12020 55334
rect 12076 55278 12086 55334
rect 12010 55192 12022 55278
rect 12074 55192 12086 55278
rect 12010 55136 12020 55192
rect 12076 55136 12086 55192
rect 12010 55050 12022 55136
rect 12074 55050 12086 55136
rect 12010 54994 12020 55050
rect 12076 54994 12086 55050
rect 12010 54987 12022 54994
rect 12074 54987 12086 54994
rect 12010 54975 12086 54987
rect 12498 55767 12574 55779
rect 12498 55760 12510 55767
rect 12562 55760 12574 55767
rect 12498 55704 12508 55760
rect 12564 55704 12574 55760
rect 12498 55618 12510 55704
rect 12562 55618 12574 55704
rect 12498 55562 12508 55618
rect 12564 55562 12574 55618
rect 12498 55476 12510 55562
rect 12562 55476 12574 55562
rect 12498 55420 12508 55476
rect 12564 55420 12574 55476
rect 12498 55334 12510 55420
rect 12562 55334 12574 55420
rect 12498 55278 12508 55334
rect 12564 55278 12574 55334
rect 12498 55192 12510 55278
rect 12562 55192 12574 55278
rect 12498 55136 12508 55192
rect 12564 55136 12574 55192
rect 12498 55050 12510 55136
rect 12562 55050 12574 55136
rect 12498 54994 12508 55050
rect 12564 54994 12574 55050
rect 12498 54987 12510 54994
rect 12562 54987 12574 54994
rect 12498 54975 12574 54987
rect 12686 55741 12762 55751
rect 12686 55685 12696 55741
rect 12752 55685 12762 55741
rect 12686 55599 12698 55685
rect 12750 55599 12762 55685
rect 12686 55543 12696 55599
rect 12752 55543 12762 55599
rect 12686 55457 12698 55543
rect 12750 55457 12762 55543
rect 12686 55401 12696 55457
rect 12752 55401 12762 55457
rect 12686 55315 12698 55401
rect 12750 55315 12762 55401
rect 12686 55259 12696 55315
rect 12752 55259 12762 55315
rect 12686 55173 12698 55259
rect 12750 55173 12762 55259
rect 12686 55117 12696 55173
rect 12752 55117 12762 55173
rect 12686 55031 12698 55117
rect 12750 55031 12762 55117
rect 12686 54975 12696 55031
rect 12752 54975 12762 55031
rect 9994 54889 10006 54975
rect 10058 54889 10070 54975
rect 9994 54833 10004 54889
rect 10060 54833 10070 54889
rect 9994 54823 10070 54833
rect 11340 54889 11352 54975
rect 11404 54889 11416 54975
rect 11340 54833 11350 54889
rect 11406 54833 11416 54889
rect 11340 54823 11416 54833
rect 12686 54889 12698 54975
rect 12750 54889 12762 54975
rect 12686 54833 12696 54889
rect 12752 54833 12762 54889
rect 13274 55729 13350 55849
rect 13274 54845 13286 55729
rect 13338 54845 13350 55729
rect 13274 54833 13350 54845
rect 12686 54823 12762 54833
rect 4162 54616 13350 54692
rect 3470 54371 3546 54383
rect 2098 53590 2347 53666
rect 1886 53450 1962 53536
rect 1886 53394 1896 53450
rect 1952 53394 1962 53450
rect 1886 53308 1962 53394
rect 1886 53252 1896 53308
rect 1952 53252 1962 53308
rect 1886 53166 1962 53252
rect 1886 53110 1896 53166
rect 1952 53110 1962 53166
rect 1886 53024 1962 53110
rect 1886 52968 1896 53024
rect 1952 52968 1962 53024
rect 3470 53383 3482 54371
rect 3534 53383 3546 54371
rect 4162 54163 4238 54616
rect 6096 54267 6172 54279
rect 4162 53451 4174 54163
rect 3470 53019 3546 53383
rect 3769 53383 4174 53451
rect 4226 53383 4238 54163
rect 3769 53371 4238 53383
rect 4750 54163 4826 54175
rect 4750 54160 4762 54163
rect 4814 54160 4826 54163
rect 4750 54104 4760 54160
rect 4816 54104 4826 54160
rect 6096 54160 6108 54267
rect 6160 54160 6172 54267
rect 4750 54018 4762 54104
rect 4814 54018 4826 54104
rect 4750 53962 4760 54018
rect 4816 53962 4826 54018
rect 4750 53876 4762 53962
rect 4814 53876 4826 53962
rect 4750 53820 4760 53876
rect 4816 53820 4826 53876
rect 4750 53734 4762 53820
rect 4814 53734 4826 53820
rect 4750 53678 4760 53734
rect 4816 53678 4826 53734
rect 4750 53592 4762 53678
rect 4814 53592 4826 53678
rect 4750 53536 4760 53592
rect 4816 53536 4826 53592
rect 4750 53450 4762 53536
rect 4814 53450 4826 53536
rect 4750 53394 4760 53450
rect 4816 53394 4826 53450
rect 4750 53383 4762 53394
rect 4814 53383 4826 53394
rect 3769 53361 4163 53371
rect 3769 53019 3863 53361
rect 4750 53308 4826 53383
rect 4750 53252 4760 53308
rect 4816 53252 4826 53308
rect 4750 53242 4826 53252
rect 4938 54099 5014 54109
rect 4938 54043 4948 54099
rect 5004 54043 5014 54099
rect 4938 54002 5014 54043
rect 4938 53957 4950 54002
rect 5002 53957 5014 54002
rect 4938 53901 4948 53957
rect 5004 53901 5014 53957
rect 4938 53815 4950 53901
rect 5002 53815 5014 53901
rect 4938 53759 4948 53815
rect 5004 53759 5014 53815
rect 4938 53673 4950 53759
rect 5002 53673 5014 53759
rect 4938 53617 4948 53673
rect 5004 53617 5014 53673
rect 4938 53531 4950 53617
rect 5002 53531 5014 53617
rect 4938 53475 4948 53531
rect 5004 53475 5014 53531
rect 4938 53430 4950 53475
rect 5002 53430 5014 53475
rect 4938 53389 5014 53430
rect 4938 53333 4948 53389
rect 5004 53333 5014 53389
rect 1886 52882 1962 52968
rect 3366 53007 3546 53019
rect 3366 52955 3378 53007
rect 3534 52955 3546 53007
rect 3366 52943 3546 52955
rect 3683 53007 3863 53019
rect 3683 52955 3695 53007
rect 3851 52955 3863 53007
rect 3683 52943 3863 52955
rect 1886 52826 1896 52882
rect 1952 52826 1962 52882
rect 1886 52816 1962 52826
rect 4938 52691 5014 53333
rect 5426 54099 5502 54109
rect 5426 54043 5436 54099
rect 5492 54043 5502 54099
rect 5426 54002 5502 54043
rect 5426 53957 5438 54002
rect 5490 53957 5502 54002
rect 5426 53901 5436 53957
rect 5492 53901 5502 53957
rect 5426 53815 5438 53901
rect 5490 53815 5502 53901
rect 5426 53759 5436 53815
rect 5492 53759 5502 53815
rect 5426 53673 5438 53759
rect 5490 53673 5502 53759
rect 5426 53617 5436 53673
rect 5492 53617 5502 53673
rect 5426 53531 5438 53617
rect 5490 53531 5502 53617
rect 5426 53475 5436 53531
rect 5492 53475 5502 53531
rect 5426 53430 5438 53475
rect 5490 53430 5502 53475
rect 5426 53389 5502 53430
rect 5426 53333 5436 53389
rect 5492 53333 5502 53389
rect 5426 53323 5502 53333
rect 5914 54099 5990 54109
rect 5914 54043 5924 54099
rect 5980 54043 5990 54099
rect 5914 54002 5990 54043
rect 5914 53957 5926 54002
rect 5978 53957 5990 54002
rect 5914 53901 5924 53957
rect 5980 53901 5990 53957
rect 5914 53815 5926 53901
rect 5978 53815 5990 53901
rect 5914 53759 5924 53815
rect 5980 53759 5990 53815
rect 5914 53673 5926 53759
rect 5978 53673 5990 53759
rect 5914 53617 5924 53673
rect 5980 53617 5990 53673
rect 5914 53531 5926 53617
rect 5978 53531 5990 53617
rect 5914 53475 5924 53531
rect 5980 53475 5990 53531
rect 5914 53430 5926 53475
rect 5978 53430 5990 53475
rect 5914 53389 5990 53430
rect 5914 53333 5924 53389
rect 5980 53333 5990 53389
rect 5914 53323 5990 53333
rect 6096 54104 6106 54160
rect 6162 54104 6172 54160
rect 7442 54163 7518 54175
rect 7442 54160 7454 54163
rect 7506 54160 7518 54163
rect 6096 54018 6108 54104
rect 6160 54018 6172 54104
rect 6096 53962 6106 54018
rect 6162 53962 6172 54018
rect 6096 53876 6108 53962
rect 6160 53876 6172 53962
rect 6096 53820 6106 53876
rect 6162 53820 6172 53876
rect 6096 53734 6108 53820
rect 6160 53734 6172 53820
rect 6096 53678 6106 53734
rect 6162 53678 6172 53734
rect 6096 53592 6108 53678
rect 6160 53592 6172 53678
rect 6096 53536 6106 53592
rect 6162 53536 6172 53592
rect 6096 53450 6108 53536
rect 6160 53450 6172 53536
rect 6096 53394 6106 53450
rect 6162 53394 6172 53450
rect 6096 53383 6108 53394
rect 6160 53383 6172 53394
rect 6096 53308 6172 53383
rect 6278 54099 6354 54109
rect 6278 54043 6288 54099
rect 6344 54043 6354 54099
rect 6278 54002 6354 54043
rect 6278 53957 6290 54002
rect 6342 53957 6354 54002
rect 6278 53901 6288 53957
rect 6344 53901 6354 53957
rect 6278 53815 6290 53901
rect 6342 53815 6354 53901
rect 6278 53759 6288 53815
rect 6344 53759 6354 53815
rect 6278 53673 6290 53759
rect 6342 53673 6354 53759
rect 6278 53617 6288 53673
rect 6344 53617 6354 53673
rect 6278 53531 6290 53617
rect 6342 53531 6354 53617
rect 6278 53475 6288 53531
rect 6344 53475 6354 53531
rect 6278 53430 6290 53475
rect 6342 53430 6354 53475
rect 6278 53389 6354 53430
rect 6278 53333 6288 53389
rect 6344 53333 6354 53389
rect 6278 53323 6354 53333
rect 6766 54099 6842 54109
rect 6766 54043 6776 54099
rect 6832 54043 6842 54099
rect 6766 54002 6842 54043
rect 6766 53957 6778 54002
rect 6830 53957 6842 54002
rect 6766 53901 6776 53957
rect 6832 53901 6842 53957
rect 6766 53815 6778 53901
rect 6830 53815 6842 53901
rect 6766 53759 6776 53815
rect 6832 53759 6842 53815
rect 6766 53673 6778 53759
rect 6830 53673 6842 53759
rect 6766 53617 6776 53673
rect 6832 53617 6842 53673
rect 6766 53531 6778 53617
rect 6830 53531 6842 53617
rect 6766 53475 6776 53531
rect 6832 53475 6842 53531
rect 6766 53430 6778 53475
rect 6830 53430 6842 53475
rect 6766 53389 6842 53430
rect 6766 53333 6776 53389
rect 6832 53333 6842 53389
rect 6096 53252 6106 53308
rect 6162 53252 6172 53308
rect 6096 53242 6172 53252
rect 6766 52691 6842 53333
rect 7254 54099 7330 54109
rect 7254 54043 7264 54099
rect 7320 54043 7330 54099
rect 7254 54002 7330 54043
rect 7254 53957 7266 54002
rect 7318 53957 7330 54002
rect 7254 53901 7264 53957
rect 7320 53901 7330 53957
rect 7254 53815 7266 53901
rect 7318 53815 7330 53901
rect 7254 53759 7264 53815
rect 7320 53759 7330 53815
rect 7254 53673 7266 53759
rect 7318 53673 7330 53759
rect 7254 53617 7264 53673
rect 7320 53617 7330 53673
rect 7254 53531 7266 53617
rect 7318 53531 7330 53617
rect 7254 53475 7264 53531
rect 7320 53475 7330 53531
rect 7254 53430 7266 53475
rect 7318 53430 7330 53475
rect 7254 53389 7330 53430
rect 7254 53333 7264 53389
rect 7320 53333 7330 53389
rect 7254 52691 7330 53333
rect 7442 54104 7452 54160
rect 7508 54104 7518 54160
rect 7442 54018 7454 54104
rect 7506 54018 7518 54104
rect 7442 53962 7452 54018
rect 7508 53962 7518 54018
rect 7442 53876 7454 53962
rect 7506 53876 7518 53962
rect 7442 53820 7452 53876
rect 7508 53820 7518 53876
rect 7442 53734 7454 53820
rect 7506 53734 7518 53820
rect 7442 53678 7452 53734
rect 7508 53678 7518 53734
rect 7442 53592 7454 53678
rect 7506 53592 7518 53678
rect 7442 53536 7452 53592
rect 7508 53536 7518 53592
rect 7442 53450 7454 53536
rect 7506 53450 7518 53536
rect 7442 53394 7452 53450
rect 7508 53394 7518 53450
rect 7442 53383 7454 53394
rect 7506 53383 7518 53394
rect 7442 53308 7518 53383
rect 8030 54163 8106 54616
rect 8030 53383 8042 54163
rect 8094 53383 8106 54163
rect 8030 53371 8106 53383
rect 8718 54371 8794 54616
rect 8718 53383 8730 54371
rect 8782 53383 8794 54371
rect 11340 54267 11416 54279
rect 7442 53252 7452 53308
rect 7508 53252 7518 53308
rect 7442 53242 7518 53252
rect 8718 52839 8794 53383
rect 9149 54160 9549 54200
rect 9149 54104 9179 54160
rect 9235 54104 9321 54160
rect 9377 54104 9463 54160
rect 9519 54104 9549 54160
rect 9149 54018 9549 54104
rect 9149 53962 9179 54018
rect 9235 53962 9321 54018
rect 9377 53962 9463 54018
rect 9519 53962 9549 54018
rect 9149 53876 9549 53962
rect 9149 53820 9179 53876
rect 9235 53820 9321 53876
rect 9377 53820 9463 53876
rect 9519 53820 9549 53876
rect 9149 53734 9549 53820
rect 9149 53678 9179 53734
rect 9235 53678 9321 53734
rect 9377 53678 9463 53734
rect 9519 53678 9549 53734
rect 9149 53592 9549 53678
rect 9149 53536 9179 53592
rect 9235 53536 9321 53592
rect 9377 53536 9463 53592
rect 9519 53536 9549 53592
rect 9149 53450 9549 53536
rect 9149 53394 9179 53450
rect 9235 53394 9321 53450
rect 9377 53394 9463 53450
rect 9519 53394 9549 53450
rect 9149 53308 9549 53394
rect 9149 53252 9179 53308
rect 9235 53252 9321 53308
rect 9377 53252 9463 53308
rect 9519 53252 9549 53308
rect 9149 53166 9549 53252
rect 9994 54163 10070 54175
rect 9994 54160 10006 54163
rect 10058 54160 10070 54163
rect 9994 54104 10004 54160
rect 10060 54104 10070 54160
rect 11340 54160 11352 54267
rect 11404 54160 11416 54267
rect 9994 54018 10006 54104
rect 10058 54018 10070 54104
rect 9994 53962 10004 54018
rect 10060 53962 10070 54018
rect 9994 53876 10006 53962
rect 10058 53876 10070 53962
rect 9994 53820 10004 53876
rect 10060 53820 10070 53876
rect 9994 53734 10006 53820
rect 10058 53734 10070 53820
rect 9994 53678 10004 53734
rect 10060 53678 10070 53734
rect 9994 53592 10006 53678
rect 10058 53592 10070 53678
rect 9994 53536 10004 53592
rect 10060 53536 10070 53592
rect 9994 53450 10006 53536
rect 10058 53450 10070 53536
rect 9994 53394 10004 53450
rect 10060 53394 10070 53450
rect 9994 53383 10006 53394
rect 10058 53383 10070 53394
rect 9994 53308 10070 53383
rect 10182 54099 10258 54109
rect 10182 54043 10192 54099
rect 10248 54043 10258 54099
rect 10182 54002 10258 54043
rect 10182 53957 10194 54002
rect 10246 53957 10258 54002
rect 10182 53901 10192 53957
rect 10248 53901 10258 53957
rect 10182 53815 10194 53901
rect 10246 53815 10258 53901
rect 10182 53759 10192 53815
rect 10248 53759 10258 53815
rect 10182 53673 10194 53759
rect 10246 53673 10258 53759
rect 10182 53617 10192 53673
rect 10248 53617 10258 53673
rect 10182 53531 10194 53617
rect 10246 53531 10258 53617
rect 10182 53475 10192 53531
rect 10248 53475 10258 53531
rect 10182 53430 10194 53475
rect 10246 53430 10258 53475
rect 10182 53389 10258 53430
rect 10182 53333 10192 53389
rect 10248 53333 10258 53389
rect 10182 53323 10258 53333
rect 10670 54099 10746 54109
rect 10670 54043 10680 54099
rect 10736 54043 10746 54099
rect 10670 54002 10746 54043
rect 10670 53957 10682 54002
rect 10734 53957 10746 54002
rect 10670 53901 10680 53957
rect 10736 53901 10746 53957
rect 10670 53815 10682 53901
rect 10734 53815 10746 53901
rect 10670 53759 10680 53815
rect 10736 53759 10746 53815
rect 10670 53673 10682 53759
rect 10734 53673 10746 53759
rect 10670 53617 10680 53673
rect 10736 53617 10746 53673
rect 10670 53531 10682 53617
rect 10734 53531 10746 53617
rect 10670 53475 10680 53531
rect 10736 53475 10746 53531
rect 10670 53430 10682 53475
rect 10734 53430 10746 53475
rect 10670 53389 10746 53430
rect 10670 53333 10680 53389
rect 10736 53333 10746 53389
rect 10670 53323 10746 53333
rect 11158 54099 11234 54109
rect 11158 54043 11168 54099
rect 11224 54043 11234 54099
rect 11158 54002 11234 54043
rect 11158 53957 11170 54002
rect 11222 53957 11234 54002
rect 11158 53901 11168 53957
rect 11224 53901 11234 53957
rect 11158 53815 11170 53901
rect 11222 53815 11234 53901
rect 11158 53759 11168 53815
rect 11224 53759 11234 53815
rect 11158 53673 11170 53759
rect 11222 53673 11234 53759
rect 11158 53617 11168 53673
rect 11224 53617 11234 53673
rect 11158 53531 11170 53617
rect 11222 53531 11234 53617
rect 11158 53475 11168 53531
rect 11224 53475 11234 53531
rect 11158 53430 11170 53475
rect 11222 53430 11234 53475
rect 11158 53389 11234 53430
rect 11158 53333 11168 53389
rect 11224 53333 11234 53389
rect 11158 53323 11234 53333
rect 11340 54104 11350 54160
rect 11406 54104 11416 54160
rect 12686 54163 12762 54175
rect 12686 54160 12698 54163
rect 12750 54160 12762 54163
rect 11340 54018 11352 54104
rect 11404 54018 11416 54104
rect 11340 53962 11350 54018
rect 11406 53962 11416 54018
rect 11340 53876 11352 53962
rect 11404 53876 11416 53962
rect 11340 53820 11350 53876
rect 11406 53820 11416 53876
rect 11340 53734 11352 53820
rect 11404 53734 11416 53820
rect 11340 53678 11350 53734
rect 11406 53678 11416 53734
rect 11340 53592 11352 53678
rect 11404 53592 11416 53678
rect 11340 53536 11350 53592
rect 11406 53536 11416 53592
rect 11340 53450 11352 53536
rect 11404 53450 11416 53536
rect 11340 53394 11350 53450
rect 11406 53394 11416 53450
rect 11340 53383 11352 53394
rect 11404 53383 11416 53394
rect 9994 53252 10004 53308
rect 10060 53252 10070 53308
rect 9994 53242 10070 53252
rect 11340 53308 11416 53383
rect 11522 54099 11598 54109
rect 11522 54043 11532 54099
rect 11588 54043 11598 54099
rect 11522 54002 11598 54043
rect 11522 53957 11534 54002
rect 11586 53957 11598 54002
rect 11522 53901 11532 53957
rect 11588 53901 11598 53957
rect 11522 53815 11534 53901
rect 11586 53815 11598 53901
rect 11522 53759 11532 53815
rect 11588 53759 11598 53815
rect 11522 53673 11534 53759
rect 11586 53673 11598 53759
rect 11522 53617 11532 53673
rect 11588 53617 11598 53673
rect 11522 53531 11534 53617
rect 11586 53531 11598 53617
rect 11522 53475 11532 53531
rect 11588 53475 11598 53531
rect 11522 53430 11534 53475
rect 11586 53430 11598 53475
rect 11522 53389 11598 53430
rect 11522 53333 11532 53389
rect 11588 53333 11598 53389
rect 11522 53323 11598 53333
rect 12010 54099 12086 54109
rect 12010 54043 12020 54099
rect 12076 54043 12086 54099
rect 12010 54002 12086 54043
rect 12010 53957 12022 54002
rect 12074 53957 12086 54002
rect 12010 53901 12020 53957
rect 12076 53901 12086 53957
rect 12010 53815 12022 53901
rect 12074 53815 12086 53901
rect 12010 53759 12020 53815
rect 12076 53759 12086 53815
rect 12010 53673 12022 53759
rect 12074 53673 12086 53759
rect 12010 53617 12020 53673
rect 12076 53617 12086 53673
rect 12010 53531 12022 53617
rect 12074 53531 12086 53617
rect 12010 53475 12020 53531
rect 12076 53475 12086 53531
rect 12010 53430 12022 53475
rect 12074 53430 12086 53475
rect 12010 53389 12086 53430
rect 12010 53333 12020 53389
rect 12076 53333 12086 53389
rect 12010 53323 12086 53333
rect 12498 54099 12574 54109
rect 12498 54043 12508 54099
rect 12564 54043 12574 54099
rect 12498 54002 12574 54043
rect 12498 53957 12510 54002
rect 12562 53957 12574 54002
rect 12498 53901 12508 53957
rect 12564 53901 12574 53957
rect 12498 53815 12510 53901
rect 12562 53815 12574 53901
rect 12498 53759 12508 53815
rect 12564 53759 12574 53815
rect 12498 53673 12510 53759
rect 12562 53673 12574 53759
rect 12498 53617 12508 53673
rect 12564 53617 12574 53673
rect 12498 53531 12510 53617
rect 12562 53531 12574 53617
rect 12498 53475 12508 53531
rect 12564 53475 12574 53531
rect 12498 53430 12510 53475
rect 12562 53430 12574 53475
rect 12498 53389 12574 53430
rect 12498 53333 12508 53389
rect 12564 53333 12574 53389
rect 12498 53323 12574 53333
rect 12686 54104 12696 54160
rect 12752 54104 12762 54160
rect 12686 54018 12698 54104
rect 12750 54018 12762 54104
rect 12686 53962 12696 54018
rect 12752 53962 12762 54018
rect 12686 53876 12698 53962
rect 12750 53876 12762 53962
rect 12686 53820 12696 53876
rect 12752 53820 12762 53876
rect 12686 53734 12698 53820
rect 12750 53734 12762 53820
rect 12686 53678 12696 53734
rect 12752 53678 12762 53734
rect 12686 53592 12698 53678
rect 12750 53592 12762 53678
rect 12686 53536 12696 53592
rect 12752 53536 12762 53592
rect 12686 53450 12698 53536
rect 12750 53450 12762 53536
rect 12686 53394 12696 53450
rect 12752 53394 12762 53450
rect 12686 53383 12698 53394
rect 12750 53383 12762 53394
rect 11340 53252 11350 53308
rect 11406 53252 11416 53308
rect 11340 53242 11416 53252
rect 12686 53308 12762 53383
rect 13274 54163 13350 54616
rect 13274 53383 13286 54163
rect 13338 53383 13350 54163
rect 13274 53371 13350 53383
rect 12686 53252 12696 53308
rect 12752 53252 12762 53308
rect 12686 53242 12762 53252
rect 9149 53110 9179 53166
rect 9235 53110 9321 53166
rect 9377 53110 9463 53166
rect 9519 53110 9549 53166
rect 9149 53024 9549 53110
rect 9149 52968 9179 53024
rect 9235 52968 9321 53024
rect 9377 52968 9463 53024
rect 9519 52968 9549 53024
rect 9149 52882 9549 52968
rect 9149 52826 9179 52882
rect 9235 52826 9321 52882
rect 9377 52826 9463 52882
rect 9519 52826 9549 52882
rect 9149 52777 9549 52826
rect 4734 52679 5226 52691
rect 4734 52627 4746 52679
rect 5214 52627 5226 52679
rect 4734 52615 5226 52627
rect 6438 52679 6930 52691
rect 6438 52627 6450 52679
rect 6918 52627 6930 52679
rect 6438 52615 6930 52627
rect 7254 52679 7434 52691
rect 7254 52627 7266 52679
rect 7422 52627 7434 52679
rect 7254 52615 7434 52627
rect 9149 51265 9425 52777
rect 1852 50269 6816 50281
rect 1852 50217 1864 50269
rect 6804 50217 6816 50269
rect 1852 50205 6816 50217
rect 4594 49424 4994 50205
rect 4594 49372 4644 49424
rect 4696 49372 4768 49424
rect 4820 49372 4892 49424
rect 4944 49372 4994 49424
rect 4594 49300 4994 49372
rect 4594 49248 4644 49300
rect 4696 49248 4768 49300
rect 4820 49248 4892 49300
rect 4944 49248 4994 49300
rect 4594 49176 4994 49248
rect 4594 49124 4644 49176
rect 4696 49124 4768 49176
rect 4820 49124 4892 49176
rect 4944 49124 4994 49176
rect 4594 49052 4994 49124
rect 5513 49398 5913 50205
rect 5513 49138 5531 49398
rect 5895 49138 5913 49398
rect 5513 49080 5913 49138
rect 6416 49398 6816 50205
rect 7714 50269 8114 50281
rect 7714 50217 7732 50269
rect 8096 50217 8114 50269
rect 6416 49138 6434 49398
rect 6798 49138 6816 49398
rect 6416 49080 6816 49138
rect 4594 49000 4644 49052
rect 4696 49000 4768 49052
rect 4820 49000 4892 49052
rect 4944 49000 4994 49052
rect 4594 48928 4994 49000
rect 4594 48876 4644 48928
rect 4696 48876 4768 48928
rect 4820 48876 4892 48928
rect 4944 48876 4994 48928
rect 4594 48804 4994 48876
rect 4594 48752 4644 48804
rect 4696 48752 4768 48804
rect 4820 48752 4892 48804
rect 4944 48752 4994 48804
rect 4594 48680 4994 48752
rect 4594 48628 4644 48680
rect 4696 48628 4768 48680
rect 4820 48628 4892 48680
rect 4944 48628 4994 48680
rect 4594 48556 4994 48628
rect 4594 48504 4644 48556
rect 4696 48504 4768 48556
rect 4820 48504 4892 48556
rect 4944 48504 4994 48556
rect 4594 48432 4994 48504
rect 4594 48380 4644 48432
rect 4696 48380 4768 48432
rect 4820 48380 4892 48432
rect 4944 48380 4994 48432
rect 4594 48308 4994 48380
rect 4594 48256 4644 48308
rect 4696 48256 4768 48308
rect 4820 48256 4892 48308
rect 4944 48256 4994 48308
rect 4594 48184 4994 48256
rect 4594 48132 4644 48184
rect 4696 48132 4768 48184
rect 4820 48132 4892 48184
rect 4944 48132 4994 48184
rect 4594 48060 4994 48132
rect 4594 48008 4644 48060
rect 4696 48008 4768 48060
rect 4820 48008 4892 48060
rect 4944 48008 4994 48060
rect 4594 47936 4994 48008
rect 4594 47884 4644 47936
rect 4696 47884 4768 47936
rect 4820 47884 4892 47936
rect 4944 47884 4994 47936
rect 3608 47788 3684 47800
rect 3608 47760 3620 47788
rect 3672 47760 3684 47788
rect 3608 47704 3618 47760
rect 3674 47704 3684 47760
rect 3608 47618 3620 47704
rect 3672 47618 3684 47704
rect 3608 47562 3618 47618
rect 3674 47562 3684 47618
rect 3608 47476 3620 47562
rect 3672 47476 3684 47562
rect 3608 47420 3618 47476
rect 3674 47420 3684 47476
rect 3608 47334 3620 47420
rect 3672 47334 3684 47420
rect 3608 47278 3618 47334
rect 3674 47278 3684 47334
rect 3608 47192 3620 47278
rect 3672 47192 3684 47278
rect 3608 47136 3618 47192
rect 3674 47136 3684 47192
rect 3608 47050 3620 47136
rect 3672 47050 3684 47136
rect 3608 46994 3618 47050
rect 3674 46994 3684 47050
rect 3608 46908 3620 46994
rect 3672 46908 3684 46994
rect 3608 46852 3618 46908
rect 3674 46852 3684 46908
rect 3608 46766 3620 46852
rect 3672 46766 3684 46852
rect 3608 46710 3618 46766
rect 3674 46710 3684 46766
rect 3608 46696 3620 46710
rect 3672 46696 3684 46710
rect 3608 46684 3684 46696
rect 4594 46620 4994 47884
rect 3158 46504 4378 46520
rect 3158 46036 3197 46504
rect 3353 46036 4378 46504
rect 3158 46020 4378 46036
rect 7427 46020 7627 49561
rect 7714 49398 8114 50217
rect 7714 49138 7732 49398
rect 8096 49138 8114 49398
rect 7714 49080 8114 49138
rect 8416 50269 8816 50281
rect 8416 50217 8434 50269
rect 8798 50217 8816 50269
rect 8416 49398 8816 50217
rect 8416 49138 8434 49398
rect 8798 49138 8816 49398
rect 8416 49080 8816 49138
rect 9149 48662 9549 51265
rect 11574 49902 11762 49912
rect 11574 49846 11584 49902
rect 11640 49846 11696 49902
rect 11752 49846 11762 49902
rect 11574 49790 11762 49846
rect 11574 49734 11584 49790
rect 11640 49734 11696 49790
rect 11752 49734 11762 49790
rect 11574 49678 11762 49734
rect 11574 49622 11584 49678
rect 11640 49622 11696 49678
rect 11752 49622 11762 49678
rect 11574 49612 11762 49622
rect 10782 49360 10858 49372
rect 10782 49304 10792 49360
rect 10848 49304 10858 49360
rect 10782 49218 10794 49304
rect 10846 49218 10858 49304
rect 10782 49162 10792 49218
rect 10848 49162 10858 49218
rect 10782 49076 10794 49162
rect 10846 49076 10858 49162
rect 10782 49020 10792 49076
rect 10848 49020 10858 49076
rect 10782 48934 10794 49020
rect 10846 48934 10858 49020
rect 10782 48878 10792 48934
rect 10848 48878 10858 48934
rect 10782 48792 10794 48878
rect 10846 48792 10858 48878
rect 10782 48736 10792 48792
rect 10848 48736 10858 48792
rect 10782 48650 10794 48736
rect 10846 48650 10858 48736
rect 10782 48594 10792 48650
rect 10848 48594 10858 48650
rect 10782 48508 10794 48594
rect 10846 48508 10858 48594
rect 10782 48452 10792 48508
rect 10848 48452 10858 48508
rect 10782 48372 10794 48452
rect 10846 48372 10858 48452
rect 10782 48366 10858 48372
rect 10782 48310 10792 48366
rect 10848 48310 10858 48366
rect 10782 48300 10858 48310
rect 10424 48036 10642 48046
rect 9713 46200 9931 48031
rect 10424 47980 10434 48036
rect 10594 47980 10642 48036
rect 10424 47970 10642 47980
rect 10566 46330 10642 47970
rect 11589 47942 11742 49612
rect 11589 47786 11630 47942
rect 11682 47786 11742 47942
rect 11589 47774 11742 47786
rect 11001 47744 11077 47754
rect 11001 47688 11011 47744
rect 11067 47688 11077 47744
rect 11001 47602 11013 47688
rect 11065 47602 11077 47688
rect 11001 47546 11011 47602
rect 11067 47546 11077 47602
rect 11001 47460 11013 47546
rect 11065 47460 11077 47546
rect 11001 47404 11011 47460
rect 11067 47404 11077 47460
rect 11001 47318 11013 47404
rect 11065 47318 11077 47404
rect 11001 47262 11011 47318
rect 11067 47262 11077 47318
rect 11001 47176 11013 47262
rect 11065 47176 11077 47262
rect 11001 47120 11011 47176
rect 11067 47120 11077 47176
rect 11001 47110 11077 47120
rect 12260 46966 12660 46978
rect 12260 46914 12272 46966
rect 12324 46914 12380 46966
rect 12432 46914 12488 46966
rect 12540 46914 12596 46966
rect 12648 46914 12660 46966
rect 12260 46902 12660 46914
rect 10566 46254 10964 46330
rect 9713 44800 10470 46200
rect 10888 46170 10964 46254
rect 10888 46126 11093 46170
rect 10888 44822 10898 46126
rect 10954 44822 11027 46126
rect 11083 44822 11093 46126
rect 10888 44770 11093 44822
rect 3608 44560 3684 44570
rect 3608 44504 3618 44560
rect 3674 44504 3684 44560
rect 3608 44418 3620 44504
rect 3672 44418 3684 44504
rect 3608 44362 3618 44418
rect 3674 44362 3684 44418
rect 3608 44276 3620 44362
rect 3672 44276 3684 44362
rect 3608 44220 3618 44276
rect 3674 44220 3684 44276
rect 3608 44134 3620 44220
rect 3672 44134 3684 44220
rect 3608 44078 3618 44134
rect 3674 44078 3684 44134
rect 3608 43992 3620 44078
rect 3672 43992 3684 44078
rect 3608 43936 3618 43992
rect 3674 43936 3684 43992
rect 3608 43850 3620 43936
rect 3672 43850 3684 43936
rect 3608 43794 3618 43850
rect 3674 43794 3684 43850
rect 3608 43708 3620 43794
rect 3672 43708 3684 43794
rect 3608 43652 3618 43708
rect 3674 43652 3684 43708
rect 3608 43566 3620 43652
rect 3672 43566 3684 43652
rect 3608 43510 3618 43566
rect 3674 43510 3684 43566
rect 3608 43424 3620 43510
rect 3672 43424 3684 43510
rect 3608 43368 3618 43424
rect 3674 43368 3684 43424
rect 3608 43282 3620 43368
rect 3672 43282 3684 43368
rect 3608 43226 3618 43282
rect 3674 43226 3684 43282
rect 3608 43216 3684 43226
rect 3608 42960 3684 42970
rect 3608 42904 3618 42960
rect 3674 42904 3684 42960
rect 3608 42818 3620 42904
rect 3672 42818 3684 42904
rect 3608 42762 3618 42818
rect 3674 42762 3684 42818
rect 3608 42676 3620 42762
rect 3672 42676 3684 42762
rect 3608 42620 3618 42676
rect 3674 42620 3684 42676
rect 3608 42534 3620 42620
rect 3672 42534 3684 42620
rect 3608 42478 3618 42534
rect 3674 42478 3684 42534
rect 3608 42392 3620 42478
rect 3672 42392 3684 42478
rect 3608 42336 3618 42392
rect 3674 42336 3684 42392
rect 3608 42250 3620 42336
rect 3672 42250 3684 42336
rect 3608 42194 3618 42250
rect 3674 42194 3684 42250
rect 3608 42108 3620 42194
rect 3672 42108 3684 42194
rect 3608 42052 3618 42108
rect 3674 42052 3684 42108
rect 3608 41966 3620 42052
rect 3672 41966 3684 42052
rect 3608 41910 3618 41966
rect 3674 41910 3684 41966
rect 3608 41824 3620 41910
rect 3672 41824 3684 41910
rect 3608 41768 3618 41824
rect 3674 41768 3684 41824
rect 3608 41682 3620 41768
rect 3672 41682 3684 41768
rect 3608 41626 3618 41682
rect 3674 41626 3684 41682
rect 3608 41616 3684 41626
rect 1836 41072 3758 41082
rect 1836 41016 1846 41072
rect 1902 41070 1988 41072
rect 2044 41070 2130 41072
rect 2186 41070 2272 41072
rect 2328 41070 2414 41072
rect 2470 41070 2556 41072
rect 2612 41070 2698 41072
rect 2754 41070 2840 41072
rect 2896 41070 2982 41072
rect 3038 41070 3124 41072
rect 3180 41070 3266 41072
rect 3322 41070 3408 41072
rect 3464 41070 3550 41072
rect 3606 41070 3692 41072
rect 3668 41018 3692 41070
rect 1902 41016 1988 41018
rect 2044 41016 2130 41018
rect 2186 41016 2272 41018
rect 2328 41016 2414 41018
rect 2470 41016 2556 41018
rect 2612 41016 2698 41018
rect 2754 41016 2840 41018
rect 2896 41016 2982 41018
rect 3038 41016 3124 41018
rect 3180 41016 3266 41018
rect 3322 41016 3408 41018
rect 3464 41016 3550 41018
rect 3606 41016 3692 41018
rect 3748 41016 3758 41072
rect 1836 41006 3758 41016
rect 1913 40734 2093 40746
rect 1913 40682 1925 40734
rect 2081 40682 2093 40734
rect 1913 40670 2093 40682
rect 4837 40734 5017 40746
rect 4837 40682 4849 40734
rect 5005 40682 5017 40734
rect 4837 40670 5017 40682
rect 7053 40734 7233 40746
rect 7053 40682 7065 40734
rect 7221 40682 7233 40734
rect 7053 40670 7233 40682
rect 1596 40568 1776 40580
rect 1596 40516 1608 40568
rect 1764 40516 1776 40568
rect 1596 40504 1776 40516
rect 1184 39027 1260 40503
rect 1771 39788 1847 39800
rect 1771 39760 1783 39788
rect 1835 39760 1847 39788
rect 1771 39704 1781 39760
rect 1837 39704 1847 39760
rect 1771 39618 1783 39704
rect 1835 39618 1847 39704
rect 1771 39562 1781 39618
rect 1837 39562 1847 39618
rect 1771 39476 1783 39562
rect 1835 39476 1847 39562
rect 1771 39420 1781 39476
rect 1837 39420 1847 39476
rect 1771 39334 1783 39420
rect 1835 39334 1847 39420
rect 1771 39278 1781 39334
rect 1837 39278 1847 39334
rect 1771 39216 1783 39278
rect 1835 39216 1847 39278
rect 1771 39192 1847 39216
rect 1771 39136 1781 39192
rect 1837 39136 1847 39192
rect 1771 39126 1847 39136
rect 1913 39057 1989 40670
rect 2357 40316 4563 40326
rect 2357 40260 2367 40316
rect 2423 40314 2509 40316
rect 2565 40314 2651 40316
rect 2707 40314 2793 40316
rect 2849 40314 2935 40316
rect 2991 40314 3077 40316
rect 3133 40314 3219 40316
rect 3275 40314 3361 40316
rect 3417 40314 3503 40316
rect 3559 40314 3645 40316
rect 3701 40314 3787 40316
rect 3843 40314 3929 40316
rect 3985 40314 4071 40316
rect 4127 40314 4213 40316
rect 4269 40314 4355 40316
rect 4411 40314 4497 40316
rect 2423 40262 2445 40314
rect 4473 40262 4497 40314
rect 2423 40260 2509 40262
rect 2565 40260 2651 40262
rect 2707 40260 2793 40262
rect 2849 40260 2935 40262
rect 2991 40260 3077 40262
rect 3133 40260 3219 40262
rect 3275 40260 3361 40262
rect 3417 40260 3503 40262
rect 3559 40260 3645 40262
rect 3701 40260 3787 40262
rect 3843 40260 3929 40262
rect 3985 40260 4071 40262
rect 4127 40260 4213 40262
rect 4269 40260 4355 40262
rect 4411 40260 4497 40262
rect 4553 40260 4563 40316
rect 2357 40250 4563 40260
rect 4941 39057 5017 40670
rect 5566 40568 5746 40580
rect 5566 40516 5578 40568
rect 5734 40516 5746 40568
rect 5566 40504 5746 40516
rect 5083 39760 5159 39770
rect 5083 39704 5093 39760
rect 5149 39704 5159 39760
rect 5083 39618 5095 39704
rect 5147 39618 5159 39704
rect 5083 39562 5093 39618
rect 5149 39562 5159 39618
rect 5083 39476 5095 39562
rect 5147 39476 5159 39562
rect 5083 39420 5093 39476
rect 5149 39420 5159 39476
rect 5083 39334 5095 39420
rect 5147 39334 5159 39420
rect 5083 39278 5093 39334
rect 5149 39278 5159 39334
rect 5083 39192 5095 39278
rect 5147 39192 5159 39278
rect 5083 39136 5093 39192
rect 5149 39136 5159 39192
rect 5083 39126 5159 39136
rect 5670 39027 5746 40504
rect 6049 39758 6125 39770
rect 6049 39754 6061 39758
rect 6113 39754 6125 39758
rect 6049 39698 6059 39754
rect 6115 39698 6125 39754
rect 6049 39612 6061 39698
rect 6113 39612 6125 39698
rect 6049 39556 6059 39612
rect 6115 39556 6125 39612
rect 6049 39470 6061 39556
rect 6113 39470 6125 39556
rect 6049 39414 6059 39470
rect 6115 39414 6125 39470
rect 6049 39328 6061 39414
rect 6113 39328 6125 39414
rect 6049 39272 6059 39328
rect 6115 39272 6125 39328
rect 6049 39186 6061 39272
rect 6113 39186 6125 39272
rect 6049 39130 6059 39186
rect 6115 39130 6125 39186
rect 6049 39044 6061 39130
rect 6113 39044 6125 39130
rect 7015 39760 7091 39770
rect 7015 39704 7025 39760
rect 7081 39704 7091 39760
rect 7015 39618 7027 39704
rect 7079 39618 7091 39704
rect 7015 39562 7025 39618
rect 7081 39562 7091 39618
rect 7015 39476 7027 39562
rect 7079 39476 7091 39562
rect 7015 39420 7025 39476
rect 7081 39420 7091 39476
rect 7015 39334 7027 39420
rect 7079 39334 7091 39420
rect 7015 39278 7025 39334
rect 7081 39278 7091 39334
rect 7015 39192 7027 39278
rect 7079 39192 7091 39278
rect 7015 39136 7025 39192
rect 7081 39136 7091 39192
rect 7015 39126 7091 39136
rect 7157 39057 7233 40670
rect 6049 38988 6059 39044
rect 6115 38988 6125 39044
rect 6049 38902 6061 38988
rect 6113 38902 6125 38988
rect 6049 38846 6059 38902
rect 6115 38846 6125 38902
rect 6049 38770 6061 38846
rect 6113 38770 6125 38846
rect 6049 38760 6125 38770
rect 6049 38704 6059 38760
rect 6115 38704 6125 38760
rect 6049 38694 6125 38704
rect 32 38167 122 38200
rect 32 38111 56 38167
rect 112 38111 122 38167
rect 32 38025 58 38111
rect 110 38025 122 38111
rect 32 37969 56 38025
rect 112 37969 122 38025
rect 32 37883 58 37969
rect 110 37883 122 37969
rect 32 37827 56 37883
rect 112 37827 122 37883
rect 32 37741 58 37827
rect 110 37741 122 37827
rect 32 37685 56 37741
rect 112 37685 122 37741
rect 32 37599 58 37685
rect 110 37599 122 37685
rect 32 37543 56 37599
rect 112 37543 122 37599
rect 32 37457 58 37543
rect 110 37457 122 37543
rect 32 37401 56 37457
rect 112 37401 122 37457
rect 32 37315 58 37401
rect 110 37315 122 37401
rect 32 37259 56 37315
rect 112 37259 122 37315
rect 32 37173 58 37259
rect 110 37173 122 37259
rect 32 37117 56 37173
rect 112 37117 122 37173
rect 32 37031 58 37117
rect 110 37031 122 37117
rect 32 36975 56 37031
rect 112 36975 122 37031
rect 32 36889 58 36975
rect 110 36889 122 36975
rect 32 36833 56 36889
rect 112 36833 122 36889
rect 32 36800 122 36833
rect 704 38160 817 38512
rect 704 38104 734 38160
rect 790 38104 817 38160
rect 704 38018 817 38104
rect 704 37962 734 38018
rect 790 37962 817 38018
rect 704 37876 817 37962
rect 704 37820 734 37876
rect 790 37820 817 37876
rect 704 37734 817 37820
rect 704 37678 734 37734
rect 790 37678 817 37734
rect 704 37592 817 37678
rect 704 37536 734 37592
rect 790 37536 817 37592
rect 704 37524 817 37536
rect 869 38160 1104 38512
rect 869 38104 876 38160
rect 932 38104 1018 38160
rect 1074 38104 1104 38160
rect 869 38018 1104 38104
rect 869 37962 876 38018
rect 932 37962 1018 38018
rect 1074 37962 1104 38018
rect 869 37876 1104 37962
rect 3427 38512 3503 38524
rect 869 37820 876 37876
rect 932 37820 1018 37876
rect 1074 37820 1104 37876
rect 869 37734 1104 37820
rect 869 37678 876 37734
rect 932 37678 1018 37734
rect 1074 37678 1104 37734
rect 869 37592 1104 37678
rect 869 37536 876 37592
rect 932 37536 1018 37592
rect 1074 37536 1104 37592
rect 869 37524 1104 37536
rect 704 37450 1104 37524
rect 704 37394 734 37450
rect 790 37394 876 37450
rect 932 37394 1018 37450
rect 1074 37394 1104 37450
rect 704 37308 1104 37394
rect 704 37252 734 37308
rect 790 37252 876 37308
rect 932 37252 1018 37308
rect 1074 37252 1104 37308
rect 704 37166 1104 37252
rect 704 37110 734 37166
rect 790 37110 876 37166
rect 932 37110 1018 37166
rect 1074 37110 1104 37166
rect 704 37024 1104 37110
rect 704 36968 734 37024
rect 790 36968 876 37024
rect 932 36968 1018 37024
rect 1074 36968 1104 37024
rect 704 36882 1104 36968
rect 704 36826 734 36882
rect 790 36826 876 36882
rect 932 36826 1018 36882
rect 1074 36826 1104 36882
rect 704 36800 1104 36826
rect 2393 37939 2783 37951
rect 2393 37783 2719 37939
rect 2771 37783 2783 37939
rect 2393 37771 2783 37783
rect 3195 37939 3271 37951
rect 3195 37783 3207 37939
rect 3259 37783 3271 37939
rect 2393 36638 2469 37771
rect 2066 36626 2469 36638
rect 165 36548 383 36600
rect 165 36492 175 36548
rect 231 36492 317 36548
rect 373 36492 383 36548
rect 2066 36574 2088 36626
rect 2452 36574 2469 36626
rect 2066 36562 2469 36574
rect 165 36406 383 36492
rect 165 36350 175 36406
rect 231 36350 317 36406
rect 373 36350 383 36406
rect 165 36264 383 36350
rect 165 36208 175 36264
rect 231 36208 317 36264
rect 373 36208 383 36264
rect 1822 36490 2002 36502
rect 1822 36438 1834 36490
rect 1990 36438 2002 36490
rect 1822 36426 2002 36438
rect 165 36122 383 36208
rect 165 36066 175 36122
rect 231 36066 317 36122
rect 373 36066 383 36122
rect 165 35980 383 36066
rect 1310 36218 1490 36230
rect 1310 36166 1322 36218
rect 1478 36166 1490 36218
rect 1310 36154 1490 36166
rect 165 35924 175 35980
rect 231 35924 317 35980
rect 373 35924 383 35980
rect 165 35838 383 35924
rect 165 35782 175 35838
rect 231 35782 317 35838
rect 373 35782 383 35838
rect 165 35696 383 35782
rect 165 35640 175 35696
rect 231 35640 317 35696
rect 373 35640 383 35696
rect 165 35554 383 35640
rect 165 35498 175 35554
rect 231 35498 317 35554
rect 373 35498 383 35554
rect 165 35412 383 35498
rect 165 35356 175 35412
rect 231 35356 317 35412
rect 373 35356 383 35412
rect 165 35270 383 35356
rect 165 35214 175 35270
rect 231 35214 317 35270
rect 373 35214 383 35270
rect 165 35128 383 35214
rect 165 35072 175 35128
rect 231 35072 317 35128
rect 373 35072 383 35128
rect 165 34986 383 35072
rect 165 34930 175 34986
rect 231 34930 317 34986
rect 373 34930 383 34986
rect 165 34844 383 34930
rect 165 34788 175 34844
rect 231 34788 317 34844
rect 373 34788 383 34844
rect 165 34702 383 34788
rect 165 34646 175 34702
rect 231 34646 317 34702
rect 373 34646 383 34702
rect 165 34560 383 34646
rect 165 34504 175 34560
rect 231 34504 317 34560
rect 373 34504 383 34560
rect 165 34418 383 34504
rect 165 34362 175 34418
rect 231 34362 317 34418
rect 373 34362 383 34418
rect 165 34276 383 34362
rect 165 34220 175 34276
rect 231 34220 317 34276
rect 373 34220 383 34276
rect 165 34134 383 34220
rect 165 34078 175 34134
rect 231 34078 317 34134
rect 373 34078 383 34134
rect 165 33992 383 34078
rect 486 35987 562 35997
rect 486 35931 496 35987
rect 552 35931 562 35987
rect 486 35845 498 35931
rect 550 35845 562 35931
rect 486 35789 496 35845
rect 552 35789 562 35845
rect 486 35703 498 35789
rect 550 35703 562 35789
rect 486 35647 496 35703
rect 552 35647 562 35703
rect 486 35561 498 35647
rect 550 35561 562 35647
rect 486 35505 496 35561
rect 552 35505 562 35561
rect 486 35419 498 35505
rect 550 35419 562 35505
rect 486 35363 496 35419
rect 552 35363 562 35419
rect 486 35277 498 35363
rect 550 35277 562 35363
rect 486 35221 496 35277
rect 552 35221 562 35277
rect 486 35135 498 35221
rect 550 35135 562 35221
rect 486 35079 496 35135
rect 552 35079 562 35135
rect 486 34993 498 35079
rect 550 34993 562 35079
rect 486 34937 496 34993
rect 552 34937 562 34993
rect 486 34851 498 34937
rect 550 34851 562 34937
rect 486 34795 496 34851
rect 552 34795 562 34851
rect 486 34709 498 34795
rect 550 34709 562 34795
rect 486 34653 496 34709
rect 552 34653 562 34709
rect 486 34567 498 34653
rect 550 34567 562 34653
rect 486 34511 496 34567
rect 552 34511 562 34567
rect 486 34425 498 34511
rect 550 34425 562 34511
rect 724 35982 800 35992
rect 724 35926 734 35982
rect 790 35926 800 35982
rect 724 35840 736 35926
rect 788 35840 800 35926
rect 724 35784 734 35840
rect 790 35784 800 35840
rect 724 35698 736 35784
rect 788 35698 800 35784
rect 724 35642 734 35698
rect 790 35642 800 35698
rect 724 35556 736 35642
rect 788 35556 800 35642
rect 724 35500 734 35556
rect 790 35500 800 35556
rect 724 35414 736 35500
rect 788 35414 800 35500
rect 724 35358 734 35414
rect 790 35358 800 35414
rect 724 35272 736 35358
rect 788 35272 800 35358
rect 724 35216 734 35272
rect 790 35216 800 35272
rect 724 35130 736 35216
rect 788 35130 800 35216
rect 724 35074 734 35130
rect 790 35074 800 35130
rect 724 34988 736 35074
rect 788 34988 800 35074
rect 724 34932 734 34988
rect 790 34932 800 34988
rect 724 34846 736 34932
rect 788 34846 800 34932
rect 724 34790 734 34846
rect 790 34790 800 34846
rect 724 34704 736 34790
rect 788 34704 800 34790
rect 724 34648 734 34704
rect 790 34648 800 34704
rect 724 34562 736 34648
rect 788 34562 800 34648
rect 724 34506 734 34562
rect 790 34506 800 34562
rect 724 34496 800 34506
rect 486 34369 496 34425
rect 552 34369 562 34425
rect 486 34283 498 34369
rect 550 34283 562 34369
rect 486 34227 496 34283
rect 552 34227 562 34283
rect 486 34141 498 34227
rect 550 34141 562 34227
rect 486 34085 496 34141
rect 552 34085 562 34141
rect 486 34075 562 34085
rect 165 33936 175 33992
rect 231 33936 317 33992
rect 373 33936 383 33992
rect 165 33850 383 33936
rect 165 33794 175 33850
rect 231 33794 317 33850
rect 373 33794 383 33850
rect 165 33708 383 33794
rect 165 33652 175 33708
rect 231 33652 317 33708
rect 373 33652 383 33708
rect 165 28632 383 33652
rect 486 33851 562 33863
rect 486 33348 498 33851
rect 550 33348 562 33851
rect 486 33292 496 33348
rect 552 33292 562 33348
rect 486 33206 498 33292
rect 550 33206 562 33292
rect 486 33150 496 33206
rect 552 33150 562 33206
rect 486 33064 498 33150
rect 550 33064 562 33150
rect 486 33008 496 33064
rect 552 33008 562 33064
rect 486 32922 498 33008
rect 550 32922 562 33008
rect 486 32866 496 32922
rect 552 32866 562 32922
rect 1310 32888 1386 36154
rect 1822 34435 1898 36426
rect 1822 34279 1834 34435
rect 1886 34279 1898 34435
rect 1822 34267 1898 34279
rect 2066 34435 2142 36562
rect 3195 36502 3271 37783
rect 3091 36490 3271 36502
rect 3091 36438 3103 36490
rect 3259 36438 3271 36490
rect 3091 36426 3271 36438
rect 3427 37524 3439 38512
rect 3491 37524 3503 38512
rect 6049 38512 6125 38524
rect 6049 38160 6061 38512
rect 6113 38160 6125 38512
rect 6049 38104 6059 38160
rect 6115 38104 6125 38160
rect 6049 38018 6061 38104
rect 6113 38018 6125 38104
rect 6049 37962 6059 38018
rect 6115 37962 6125 38018
rect 2066 34279 2078 34435
rect 2130 34279 2142 34435
rect 2066 34267 2142 34279
rect 2482 36354 2662 36366
rect 2482 36302 2494 36354
rect 2650 36302 2662 36354
rect 2482 36290 2662 36302
rect 2482 34435 2558 36290
rect 3427 36230 3503 37524
rect 3659 37939 3735 37951
rect 3659 37783 3671 37939
rect 3723 37783 3735 37939
rect 3659 36502 3735 37783
rect 4147 37939 4537 37951
rect 4147 37783 4159 37939
rect 4211 37783 4537 37939
rect 4147 37771 4537 37783
rect 4461 36638 4537 37771
rect 6049 37876 6061 37962
rect 6113 37876 6125 37962
rect 6049 37820 6059 37876
rect 6115 37820 6125 37876
rect 6049 37734 6061 37820
rect 6113 37734 6125 37820
rect 6049 37678 6059 37734
rect 6115 37678 6125 37734
rect 6049 37592 6061 37678
rect 6113 37592 6125 37678
rect 6049 37536 6059 37592
rect 6115 37536 6125 37592
rect 6049 37524 6061 37536
rect 6113 37524 6125 37536
rect 6049 37450 6125 37524
rect 6049 37394 6059 37450
rect 6115 37394 6125 37450
rect 6049 37308 6125 37394
rect 6049 37252 6059 37308
rect 6115 37252 6125 37308
rect 6049 37166 6125 37252
rect 6049 37110 6059 37166
rect 6115 37110 6125 37166
rect 6049 37024 6125 37110
rect 6049 36968 6059 37024
rect 6115 36968 6125 37024
rect 6049 36882 6125 36968
rect 6049 36826 6059 36882
rect 6115 36826 6125 36882
rect 6049 36816 6125 36826
rect 4461 36626 4641 36638
rect 4461 36574 4473 36626
rect 4629 36574 4641 36626
rect 4461 36562 4641 36574
rect 5810 36626 5990 36638
rect 5810 36574 5822 36626
rect 5978 36574 5990 36626
rect 5810 36562 5990 36574
rect 3659 36490 3839 36502
rect 3659 36438 3671 36490
rect 3827 36438 3839 36490
rect 3659 36426 3839 36438
rect 5394 36354 5574 36366
rect 5394 36302 5406 36354
rect 5562 36302 5574 36354
rect 5394 36290 5574 36302
rect 3092 36154 3503 36230
rect 3092 35982 3168 36154
rect 3092 35926 3102 35982
rect 3158 35926 3168 35982
rect 3092 35840 3104 35926
rect 3156 35840 3168 35926
rect 3092 35784 3102 35840
rect 3158 35784 3168 35840
rect 3092 35698 3104 35784
rect 3156 35698 3168 35784
rect 3092 35642 3102 35698
rect 3158 35642 3168 35698
rect 3092 35556 3104 35642
rect 3156 35556 3168 35642
rect 3092 35500 3102 35556
rect 3158 35500 3168 35556
rect 3092 35414 3104 35500
rect 3156 35414 3168 35500
rect 3092 35358 3102 35414
rect 3158 35358 3168 35414
rect 3092 35272 3104 35358
rect 3156 35272 3168 35358
rect 3092 35216 3102 35272
rect 3158 35216 3168 35272
rect 3092 35130 3104 35216
rect 3156 35130 3168 35216
rect 3092 35074 3102 35130
rect 3158 35074 3168 35130
rect 3092 34988 3104 35074
rect 3156 34988 3168 35074
rect 3092 34932 3102 34988
rect 3158 34932 3168 34988
rect 3092 34846 3104 34932
rect 3156 34846 3168 34932
rect 3092 34790 3102 34846
rect 3158 34790 3168 34846
rect 3092 34704 3104 34790
rect 3156 34704 3168 34790
rect 3092 34648 3102 34704
rect 3158 34648 3168 34704
rect 3092 34562 3104 34648
rect 3156 34562 3168 34648
rect 3092 34506 3102 34562
rect 3158 34506 3168 34562
rect 3092 34496 3168 34506
rect 3386 36082 3566 36094
rect 3386 36030 3398 36082
rect 3554 36030 3566 36082
rect 3386 36018 3566 36030
rect 3990 36086 4066 36096
rect 3990 36030 4000 36086
rect 4056 36030 4066 36086
rect 2482 34279 2494 34435
rect 2546 34279 2558 34435
rect 2482 34267 2558 34279
rect 3386 34267 3462 36018
rect 3990 35946 4066 36030
rect 4490 36082 4670 36094
rect 4490 36030 4502 36082
rect 4658 36030 4670 36082
rect 4490 36018 4670 36030
rect 3990 35944 4002 35946
rect 4054 35944 4066 35946
rect 3990 35888 4000 35944
rect 4056 35888 4066 35944
rect 3990 35802 4002 35888
rect 4054 35802 4066 35888
rect 3990 35746 4000 35802
rect 4056 35746 4066 35802
rect 3990 35660 4002 35746
rect 4054 35660 4066 35746
rect 3990 35604 4000 35660
rect 4056 35604 4066 35660
rect 3990 35518 4002 35604
rect 4054 35518 4066 35604
rect 3990 35462 4000 35518
rect 4056 35462 4066 35518
rect 3990 35376 4002 35462
rect 4054 35376 4066 35462
rect 3990 35320 4000 35376
rect 4056 35320 4066 35376
rect 3990 35234 4002 35320
rect 4054 35234 4066 35320
rect 3990 35178 4000 35234
rect 4056 35178 4066 35234
rect 3990 35092 4002 35178
rect 4054 35092 4066 35178
rect 3990 35036 4000 35092
rect 4056 35036 4066 35092
rect 3990 34950 4002 35036
rect 4054 34950 4066 35036
rect 3990 34894 4000 34950
rect 4056 34894 4066 34950
rect 3990 34808 4002 34894
rect 4054 34808 4066 34894
rect 3990 34752 4000 34808
rect 4056 34752 4066 34808
rect 3990 34666 4002 34752
rect 4054 34666 4066 34752
rect 3990 34610 4000 34666
rect 4056 34610 4066 34666
rect 3990 34524 4002 34610
rect 4054 34524 4066 34610
rect 3990 34468 4000 34524
rect 4056 34468 4066 34524
rect 3990 34382 4002 34468
rect 4054 34382 4066 34468
rect 3990 34326 4000 34382
rect 4056 34326 4066 34382
rect 3990 34240 4002 34326
rect 4054 34240 4066 34326
rect 4594 34267 4670 36018
rect 4888 35982 4964 35992
rect 4888 35926 4898 35982
rect 4954 35926 4964 35982
rect 4888 35840 4900 35926
rect 4952 35840 4964 35926
rect 4888 35784 4898 35840
rect 4954 35784 4964 35840
rect 4888 35698 4900 35784
rect 4952 35698 4964 35784
rect 4888 35642 4898 35698
rect 4954 35642 4964 35698
rect 4888 35556 4900 35642
rect 4952 35556 4964 35642
rect 4888 35500 4898 35556
rect 4954 35500 4964 35556
rect 4888 35414 4900 35500
rect 4952 35414 4964 35500
rect 4888 35358 4898 35414
rect 4954 35358 4964 35414
rect 4888 35272 4900 35358
rect 4952 35272 4964 35358
rect 4888 35216 4898 35272
rect 4954 35216 4964 35272
rect 4888 35130 4900 35216
rect 4952 35130 4964 35216
rect 4888 35074 4898 35130
rect 4954 35074 4964 35130
rect 4888 34988 4900 35074
rect 4952 34988 4964 35074
rect 4888 34932 4898 34988
rect 4954 34932 4964 34988
rect 4888 34846 4900 34932
rect 4952 34846 4964 34932
rect 4888 34790 4898 34846
rect 4954 34790 4964 34846
rect 4888 34704 4900 34790
rect 4952 34704 4964 34790
rect 4888 34648 4898 34704
rect 4954 34648 4964 34704
rect 4888 34562 4900 34648
rect 4952 34562 4964 34648
rect 4888 34506 4898 34562
rect 4954 34506 4964 34562
rect 4888 34496 4964 34506
rect 5498 34435 5574 36290
rect 5498 34279 5510 34435
rect 5562 34279 5574 34435
rect 5498 34267 5574 34279
rect 5914 34435 5990 36562
rect 6054 36490 6234 36502
rect 6054 36438 6066 36490
rect 6222 36438 6234 36490
rect 6054 36426 6234 36438
rect 5914 34279 5926 34435
rect 5978 34279 5990 34435
rect 5914 34267 5990 34279
rect 6158 34435 6234 36426
rect 6566 36218 6746 36230
rect 6566 36166 6578 36218
rect 6734 36166 6746 36218
rect 6566 36154 6746 36166
rect 6158 34279 6170 34435
rect 6222 34279 6234 34435
rect 6158 34267 6234 34279
rect 3990 34184 4000 34240
rect 4056 34184 4066 34240
rect 3990 34098 4002 34184
rect 4054 34098 4066 34184
rect 3990 34042 4000 34098
rect 4056 34042 4066 34098
rect 3990 33956 4002 34042
rect 4054 33956 4066 34042
rect 3990 33900 4000 33956
rect 4056 33900 4066 33956
rect 3990 33814 4002 33900
rect 4054 33814 4066 33900
rect 3990 33758 4000 33814
rect 4056 33758 4066 33814
rect 3990 33672 4002 33758
rect 4054 33672 4066 33758
rect 3990 33616 4000 33672
rect 4056 33616 4066 33672
rect 3990 33294 4002 33616
rect 4054 33294 4066 33616
rect 3990 33282 4066 33294
rect 3990 32905 4066 32915
rect 486 32780 498 32866
rect 550 32780 562 32866
rect 486 32724 496 32780
rect 552 32724 562 32780
rect 486 32638 498 32724
rect 550 32638 562 32724
rect 3990 32849 4000 32905
rect 4056 32849 4066 32905
rect 6670 32888 6746 36154
rect 3990 32825 4066 32849
rect 3990 32763 4002 32825
rect 4054 32763 4066 32825
rect 3990 32707 4000 32763
rect 4056 32707 4066 32763
rect 486 32582 496 32638
rect 552 32582 562 32638
rect 486 32496 498 32582
rect 550 32496 562 32582
rect 486 32440 496 32496
rect 552 32440 562 32496
rect 486 32354 498 32440
rect 550 32354 562 32440
rect 486 32298 496 32354
rect 552 32298 562 32354
rect 486 32212 498 32298
rect 550 32212 562 32298
rect 486 32156 496 32212
rect 552 32156 562 32212
rect 486 32070 498 32156
rect 550 32070 562 32156
rect 486 32014 496 32070
rect 552 32014 562 32070
rect 486 31928 498 32014
rect 550 31928 562 32014
rect 486 31872 496 31928
rect 552 31872 562 31928
rect 486 31786 498 31872
rect 550 31786 562 31872
rect 486 31730 496 31786
rect 552 31730 562 31786
rect 486 31644 498 31730
rect 550 31644 562 31730
rect 486 31588 496 31644
rect 552 31588 562 31644
rect 486 31502 498 31588
rect 550 31502 562 31588
rect 486 31446 496 31502
rect 552 31446 562 31502
rect 486 31360 498 31446
rect 550 31360 562 31446
rect 486 31304 496 31360
rect 552 31304 562 31360
rect 486 31218 498 31304
rect 550 31218 562 31304
rect 486 31162 496 31218
rect 552 31162 562 31218
rect 486 31076 498 31162
rect 550 31076 562 31162
rect 486 31020 496 31076
rect 552 31020 562 31076
rect 486 30934 498 31020
rect 550 30934 562 31020
rect 486 30878 496 30934
rect 552 30878 562 30934
rect 486 30792 498 30878
rect 550 30792 562 30878
rect 486 30736 496 30792
rect 552 30736 562 30792
rect 486 30650 498 30736
rect 550 30650 562 30736
rect 486 30594 496 30650
rect 552 30594 562 30650
rect 486 30508 498 30594
rect 550 30508 562 30594
rect 486 30452 496 30508
rect 552 30452 562 30508
rect 486 30055 498 30452
rect 550 30055 562 30452
rect 968 32692 1044 32702
rect 968 32636 978 32692
rect 1034 32636 1044 32692
rect 968 32550 980 32636
rect 1032 32550 1044 32636
rect 968 32494 978 32550
rect 1034 32494 1044 32550
rect 968 32408 980 32494
rect 1032 32408 1044 32494
rect 968 32352 978 32408
rect 1034 32352 1044 32408
rect 968 32266 980 32352
rect 1032 32266 1044 32352
rect 968 32210 978 32266
rect 1034 32210 1044 32266
rect 968 32124 980 32210
rect 1032 32124 1044 32210
rect 968 32068 978 32124
rect 1034 32068 1044 32124
rect 968 31982 980 32068
rect 1032 31982 1044 32068
rect 968 31926 978 31982
rect 1034 31926 1044 31982
rect 968 31840 980 31926
rect 1032 31840 1044 31926
rect 968 31784 978 31840
rect 1034 31784 1044 31840
rect 968 31698 980 31784
rect 1032 31698 1044 31784
rect 968 31642 978 31698
rect 1034 31642 1044 31698
rect 968 31556 980 31642
rect 1032 31556 1044 31642
rect 968 31500 978 31556
rect 1034 31500 1044 31556
rect 968 31414 980 31500
rect 1032 31414 1044 31500
rect 968 31358 978 31414
rect 1034 31358 1044 31414
rect 968 31272 980 31358
rect 1032 31272 1044 31358
rect 968 31216 978 31272
rect 1034 31216 1044 31272
rect 968 31130 980 31216
rect 1032 31130 1044 31216
rect 968 31074 978 31130
rect 1034 31074 1044 31130
rect 968 30988 980 31074
rect 1032 30988 1044 31074
rect 968 30932 978 30988
rect 1034 30932 1044 30988
rect 968 30846 980 30932
rect 1032 30846 1044 30932
rect 968 30790 978 30846
rect 1034 30790 1044 30846
rect 968 30704 980 30790
rect 1032 30704 1044 30790
rect 968 30648 978 30704
rect 1034 30648 1044 30704
rect 2360 32692 2436 32702
rect 2360 32636 2370 32692
rect 2426 32636 2436 32692
rect 2360 32550 2372 32636
rect 2424 32550 2436 32636
rect 2360 32494 2370 32550
rect 2426 32494 2436 32550
rect 2360 32408 2372 32494
rect 2424 32408 2436 32494
rect 2360 32352 2370 32408
rect 2426 32352 2436 32408
rect 2360 32266 2372 32352
rect 2424 32266 2436 32352
rect 2360 32210 2370 32266
rect 2426 32210 2436 32266
rect 2360 32124 2372 32210
rect 2424 32124 2436 32210
rect 2360 32068 2370 32124
rect 2426 32068 2436 32124
rect 2360 31982 2372 32068
rect 2424 31982 2436 32068
rect 2360 31926 2370 31982
rect 2426 31926 2436 31982
rect 2360 31840 2372 31926
rect 2424 31840 2436 31926
rect 2360 31784 2370 31840
rect 2426 31784 2436 31840
rect 2360 31698 2372 31784
rect 2424 31698 2436 31784
rect 2360 31642 2370 31698
rect 2426 31642 2436 31698
rect 2360 31556 2372 31642
rect 2424 31556 2436 31642
rect 2360 31500 2370 31556
rect 2426 31500 2436 31556
rect 2360 31414 2372 31500
rect 2424 31414 2436 31500
rect 2360 31358 2370 31414
rect 2426 31358 2436 31414
rect 2360 31272 2372 31358
rect 2424 31272 2436 31358
rect 2360 31216 2370 31272
rect 2426 31216 2436 31272
rect 2360 31130 2372 31216
rect 2424 31130 2436 31216
rect 2360 31074 2370 31130
rect 2426 31074 2436 31130
rect 2360 30988 2372 31074
rect 2424 30988 2436 31074
rect 2360 30932 2370 30988
rect 2426 30932 2436 30988
rect 2360 30846 2372 30932
rect 2424 30846 2436 30932
rect 2360 30790 2370 30846
rect 2426 30790 2436 30846
rect 2360 30704 2372 30790
rect 2424 30704 2436 30790
rect 968 30562 980 30648
rect 1032 30562 1044 30648
rect 968 30506 978 30562
rect 1034 30506 1044 30562
rect 968 30454 980 30506
rect 1032 30454 1044 30506
rect 968 30442 1044 30454
rect 1444 30678 1544 30690
rect 1444 30314 1468 30678
rect 1520 30314 1544 30678
rect 1444 30201 1544 30314
rect 486 30043 562 30055
rect 1007 30101 1544 30201
rect 1688 30678 1788 30690
rect 1688 30314 1712 30678
rect 1764 30314 1788 30678
rect 2360 30648 2370 30704
rect 2426 30648 2436 30704
rect 2360 30562 2372 30648
rect 2424 30562 2436 30648
rect 2360 30506 2370 30562
rect 2426 30506 2436 30562
rect 2360 30454 2372 30506
rect 2424 30454 2436 30506
rect 2360 30442 2436 30454
rect 2776 32692 2852 32702
rect 2776 32636 2786 32692
rect 2842 32636 2852 32692
rect 2776 32550 2788 32636
rect 2840 32550 2852 32636
rect 2776 32494 2786 32550
rect 2842 32494 2852 32550
rect 2776 32408 2788 32494
rect 2840 32408 2852 32494
rect 2776 32352 2786 32408
rect 2842 32352 2852 32408
rect 2776 32266 2788 32352
rect 2840 32266 2852 32352
rect 2776 32210 2786 32266
rect 2842 32210 2852 32266
rect 2776 32124 2788 32210
rect 2840 32124 2852 32210
rect 2776 32068 2786 32124
rect 2842 32068 2852 32124
rect 2776 31982 2788 32068
rect 2840 31982 2852 32068
rect 2776 31926 2786 31982
rect 2842 31926 2852 31982
rect 2776 31840 2788 31926
rect 2840 31840 2852 31926
rect 2776 31784 2786 31840
rect 2842 31784 2852 31840
rect 2776 31698 2788 31784
rect 2840 31698 2852 31784
rect 2776 31642 2786 31698
rect 2842 31642 2852 31698
rect 2776 31556 2788 31642
rect 2840 31556 2852 31642
rect 2776 31500 2786 31556
rect 2842 31500 2852 31556
rect 2776 31414 2788 31500
rect 2840 31414 2852 31500
rect 2776 31358 2786 31414
rect 2842 31358 2852 31414
rect 2776 31272 2788 31358
rect 2840 31272 2852 31358
rect 2776 31216 2786 31272
rect 2842 31216 2852 31272
rect 2776 31130 2788 31216
rect 2840 31130 2852 31216
rect 2776 31074 2786 31130
rect 2842 31074 2852 31130
rect 2776 30988 2788 31074
rect 2840 30988 2852 31074
rect 3264 32693 3340 32703
rect 3264 32637 3274 32693
rect 3330 32637 3340 32693
rect 3264 32551 3276 32637
rect 3328 32551 3340 32637
rect 3264 32495 3274 32551
rect 3330 32495 3340 32551
rect 3264 32409 3276 32495
rect 3328 32409 3340 32495
rect 3264 32353 3274 32409
rect 3330 32353 3340 32409
rect 3264 32267 3276 32353
rect 3328 32267 3340 32353
rect 3264 32211 3274 32267
rect 3330 32211 3340 32267
rect 3264 32125 3276 32211
rect 3328 32125 3340 32211
rect 3264 32069 3274 32125
rect 3330 32069 3340 32125
rect 3264 31983 3276 32069
rect 3328 31983 3340 32069
rect 3264 31927 3274 31983
rect 3330 31927 3340 31983
rect 3264 31841 3276 31927
rect 3328 31841 3340 31927
rect 3264 31785 3274 31841
rect 3330 31785 3340 31841
rect 3264 31699 3276 31785
rect 3328 31699 3340 31785
rect 3264 31643 3274 31699
rect 3330 31643 3340 31699
rect 3264 31557 3276 31643
rect 3328 31557 3340 31643
rect 3264 31501 3274 31557
rect 3330 31501 3340 31557
rect 3264 31415 3276 31501
rect 3328 31415 3340 31501
rect 3264 31359 3274 31415
rect 3330 31359 3340 31415
rect 3264 31273 3276 31359
rect 3328 31273 3340 31359
rect 3264 31217 3274 31273
rect 3330 31217 3340 31273
rect 3264 31131 3276 31217
rect 3328 31131 3340 31217
rect 3264 31075 3274 31131
rect 3330 31075 3340 31131
rect 3264 31065 3340 31075
rect 3752 32642 3828 32652
rect 3752 32586 3762 32642
rect 3818 32586 3828 32642
rect 3752 32500 3764 32586
rect 3816 32500 3828 32586
rect 3752 32444 3762 32500
rect 3818 32444 3828 32500
rect 3752 32358 3764 32444
rect 3816 32358 3828 32444
rect 3752 32302 3762 32358
rect 3818 32302 3828 32358
rect 3752 32216 3764 32302
rect 3816 32216 3828 32302
rect 3752 32160 3762 32216
rect 3818 32160 3828 32216
rect 3752 32074 3764 32160
rect 3816 32074 3828 32160
rect 3752 32018 3762 32074
rect 3818 32018 3828 32074
rect 3752 31932 3764 32018
rect 3816 31932 3828 32018
rect 3752 31876 3762 31932
rect 3818 31876 3828 31932
rect 3752 31790 3764 31876
rect 3816 31790 3828 31876
rect 3752 31734 3762 31790
rect 3818 31734 3828 31790
rect 3752 31648 3764 31734
rect 3816 31648 3828 31734
rect 3752 31592 3762 31648
rect 3818 31592 3828 31648
rect 3752 31506 3764 31592
rect 3816 31506 3828 31592
rect 3752 31450 3762 31506
rect 3818 31450 3828 31506
rect 3752 31364 3764 31450
rect 3816 31364 3828 31450
rect 3752 31308 3762 31364
rect 3818 31308 3828 31364
rect 3752 31222 3764 31308
rect 3816 31222 3828 31308
rect 3752 31166 3762 31222
rect 3818 31166 3828 31222
rect 3752 31080 3764 31166
rect 3816 31080 3828 31166
rect 3752 31024 3762 31080
rect 3818 31024 3828 31080
rect 3752 31014 3828 31024
rect 3990 32621 4002 32707
rect 4054 32621 4066 32707
rect 4716 32693 4792 32703
rect 3990 32565 4000 32621
rect 4056 32565 4066 32621
rect 3990 32479 4002 32565
rect 4054 32479 4066 32565
rect 3990 32423 4000 32479
rect 4056 32423 4066 32479
rect 3990 32337 4002 32423
rect 4054 32337 4066 32423
rect 3990 32281 4000 32337
rect 4056 32281 4066 32337
rect 3990 32195 4002 32281
rect 4054 32195 4066 32281
rect 3990 32139 4000 32195
rect 4056 32139 4066 32195
rect 3990 32053 4002 32139
rect 4054 32053 4066 32139
rect 3990 31997 4000 32053
rect 4056 31997 4066 32053
rect 3990 31911 4002 31997
rect 4054 31911 4066 31997
rect 3990 31855 4000 31911
rect 4056 31855 4066 31911
rect 3990 31769 4002 31855
rect 4054 31769 4066 31855
rect 3990 31713 4000 31769
rect 4056 31713 4066 31769
rect 3990 31627 4002 31713
rect 4054 31627 4066 31713
rect 3990 31571 4000 31627
rect 4056 31571 4066 31627
rect 3990 31485 4002 31571
rect 4054 31485 4066 31571
rect 3990 31429 4000 31485
rect 4056 31429 4066 31485
rect 3990 31343 4002 31429
rect 4054 31343 4066 31429
rect 3990 31287 4000 31343
rect 4056 31287 4066 31343
rect 3990 31201 4002 31287
rect 4054 31201 4066 31287
rect 3990 31145 4000 31201
rect 4056 31145 4066 31201
rect 3990 31059 4002 31145
rect 4054 31059 4066 31145
rect 3990 31003 4000 31059
rect 4056 31003 4066 31059
rect 4228 32642 4304 32652
rect 4228 32586 4238 32642
rect 4294 32586 4304 32642
rect 4228 32500 4240 32586
rect 4292 32500 4304 32586
rect 4228 32444 4238 32500
rect 4294 32444 4304 32500
rect 4228 32358 4240 32444
rect 4292 32358 4304 32444
rect 4228 32302 4238 32358
rect 4294 32302 4304 32358
rect 4228 32216 4240 32302
rect 4292 32216 4304 32302
rect 4228 32160 4238 32216
rect 4294 32160 4304 32216
rect 4228 32074 4240 32160
rect 4292 32074 4304 32160
rect 4228 32018 4238 32074
rect 4294 32018 4304 32074
rect 4228 31932 4240 32018
rect 4292 31932 4304 32018
rect 4228 31876 4238 31932
rect 4294 31876 4304 31932
rect 4228 31790 4240 31876
rect 4292 31790 4304 31876
rect 4228 31734 4238 31790
rect 4294 31734 4304 31790
rect 4228 31648 4240 31734
rect 4292 31648 4304 31734
rect 4228 31592 4238 31648
rect 4294 31592 4304 31648
rect 4228 31506 4240 31592
rect 4292 31506 4304 31592
rect 4228 31450 4238 31506
rect 4294 31450 4304 31506
rect 4228 31364 4240 31450
rect 4292 31364 4304 31450
rect 4228 31308 4238 31364
rect 4294 31308 4304 31364
rect 4228 31222 4240 31308
rect 4292 31222 4304 31308
rect 4228 31166 4238 31222
rect 4294 31166 4304 31222
rect 4228 31080 4240 31166
rect 4292 31080 4304 31166
rect 4228 31024 4238 31080
rect 4294 31024 4304 31080
rect 4716 32637 4726 32693
rect 4782 32637 4792 32693
rect 4716 32551 4728 32637
rect 4780 32551 4792 32637
rect 4716 32495 4726 32551
rect 4782 32495 4792 32551
rect 4716 32409 4728 32495
rect 4780 32409 4792 32495
rect 4716 32353 4726 32409
rect 4782 32353 4792 32409
rect 4716 32267 4728 32353
rect 4780 32267 4792 32353
rect 4716 32211 4726 32267
rect 4782 32211 4792 32267
rect 4716 32125 4728 32211
rect 4780 32125 4792 32211
rect 4716 32069 4726 32125
rect 4782 32069 4792 32125
rect 4716 31983 4728 32069
rect 4780 31983 4792 32069
rect 4716 31927 4726 31983
rect 4782 31927 4792 31983
rect 4716 31841 4728 31927
rect 4780 31841 4792 31927
rect 4716 31785 4726 31841
rect 4782 31785 4792 31841
rect 4716 31699 4728 31785
rect 4780 31699 4792 31785
rect 4716 31643 4726 31699
rect 4782 31643 4792 31699
rect 4716 31557 4728 31643
rect 4780 31557 4792 31643
rect 4716 31501 4726 31557
rect 4782 31501 4792 31557
rect 4716 31415 4728 31501
rect 4780 31415 4792 31501
rect 4716 31359 4726 31415
rect 4782 31359 4792 31415
rect 4716 31273 4728 31359
rect 4780 31273 4792 31359
rect 4716 31217 4726 31273
rect 4782 31217 4792 31273
rect 4716 31131 4728 31217
rect 4780 31131 4792 31217
rect 4716 31075 4726 31131
rect 4782 31075 4792 31131
rect 4716 31065 4792 31075
rect 5204 32693 5280 32703
rect 5204 32637 5214 32693
rect 5270 32637 5280 32693
rect 5204 32551 5216 32637
rect 5268 32551 5280 32637
rect 5204 32495 5214 32551
rect 5270 32495 5280 32551
rect 5204 32409 5216 32495
rect 5268 32409 5280 32495
rect 5204 32353 5214 32409
rect 5270 32353 5280 32409
rect 5204 32267 5216 32353
rect 5268 32267 5280 32353
rect 5204 32211 5214 32267
rect 5270 32211 5280 32267
rect 5204 32125 5216 32211
rect 5268 32125 5280 32211
rect 5204 32069 5214 32125
rect 5270 32069 5280 32125
rect 5204 31983 5216 32069
rect 5268 31983 5280 32069
rect 5204 31927 5214 31983
rect 5270 31927 5280 31983
rect 5204 31841 5216 31927
rect 5268 31841 5280 31927
rect 5204 31785 5214 31841
rect 5270 31785 5280 31841
rect 5204 31699 5216 31785
rect 5268 31699 5280 31785
rect 5204 31643 5214 31699
rect 5270 31643 5280 31699
rect 5204 31557 5216 31643
rect 5268 31557 5280 31643
rect 5204 31501 5214 31557
rect 5270 31501 5280 31557
rect 5204 31415 5216 31501
rect 5268 31415 5280 31501
rect 5204 31359 5214 31415
rect 5270 31359 5280 31415
rect 5204 31273 5216 31359
rect 5268 31273 5280 31359
rect 5204 31217 5214 31273
rect 5270 31217 5280 31273
rect 5204 31131 5216 31217
rect 5268 31131 5280 31217
rect 5204 31075 5214 31131
rect 5270 31075 5280 31131
rect 5204 31065 5280 31075
rect 5620 32693 5696 32703
rect 5620 32637 5630 32693
rect 5686 32637 5696 32693
rect 5620 32551 5632 32637
rect 5684 32551 5696 32637
rect 5620 32495 5630 32551
rect 5686 32495 5696 32551
rect 5620 32409 5632 32495
rect 5684 32409 5696 32495
rect 5620 32353 5630 32409
rect 5686 32353 5696 32409
rect 5620 32267 5632 32353
rect 5684 32267 5696 32353
rect 5620 32211 5630 32267
rect 5686 32211 5696 32267
rect 5620 32125 5632 32211
rect 5684 32125 5696 32211
rect 5620 32069 5630 32125
rect 5686 32069 5696 32125
rect 5620 31983 5632 32069
rect 5684 31983 5696 32069
rect 5620 31927 5630 31983
rect 5686 31927 5696 31983
rect 5620 31841 5632 31927
rect 5684 31841 5696 31927
rect 5620 31785 5630 31841
rect 5686 31785 5696 31841
rect 5620 31699 5632 31785
rect 5684 31699 5696 31785
rect 5620 31643 5630 31699
rect 5686 31643 5696 31699
rect 5620 31557 5632 31643
rect 5684 31557 5696 31643
rect 5620 31501 5630 31557
rect 5686 31501 5696 31557
rect 5620 31415 5632 31501
rect 5684 31415 5696 31501
rect 5620 31359 5630 31415
rect 5686 31359 5696 31415
rect 5620 31273 5632 31359
rect 5684 31273 5696 31359
rect 5620 31217 5630 31273
rect 5686 31217 5696 31273
rect 5620 31131 5632 31217
rect 5684 31131 5696 31217
rect 5620 31075 5630 31131
rect 5686 31075 5696 31131
rect 5620 31065 5696 31075
rect 7012 32692 7088 32702
rect 7012 32636 7022 32692
rect 7078 32636 7088 32692
rect 7012 32550 7024 32636
rect 7076 32550 7088 32636
rect 7012 32494 7022 32550
rect 7078 32494 7088 32550
rect 7012 32408 7024 32494
rect 7076 32408 7088 32494
rect 7012 32352 7022 32408
rect 7078 32352 7088 32408
rect 7012 32266 7024 32352
rect 7076 32266 7088 32352
rect 7012 32210 7022 32266
rect 7078 32210 7088 32266
rect 7012 32124 7024 32210
rect 7076 32124 7088 32210
rect 7012 32068 7022 32124
rect 7078 32068 7088 32124
rect 7012 31982 7024 32068
rect 7076 31982 7088 32068
rect 7012 31926 7022 31982
rect 7078 31926 7088 31982
rect 7012 31840 7024 31926
rect 7076 31840 7088 31926
rect 7012 31784 7022 31840
rect 7078 31784 7088 31840
rect 7012 31698 7024 31784
rect 7076 31698 7088 31784
rect 7012 31642 7022 31698
rect 7078 31642 7088 31698
rect 7012 31556 7024 31642
rect 7076 31556 7088 31642
rect 7012 31500 7022 31556
rect 7078 31500 7088 31556
rect 7012 31414 7024 31500
rect 7076 31414 7088 31500
rect 7012 31358 7022 31414
rect 7078 31358 7088 31414
rect 7012 31272 7024 31358
rect 7076 31272 7088 31358
rect 7012 31216 7022 31272
rect 7078 31216 7088 31272
rect 7012 31130 7024 31216
rect 7076 31130 7088 31216
rect 7012 31074 7022 31130
rect 7078 31074 7088 31130
rect 4228 31014 4304 31024
rect 3990 30993 4066 31003
rect 2776 30932 2786 30988
rect 2842 30932 2852 30988
rect 2776 30846 2788 30932
rect 2840 30846 2852 30932
rect 7012 30988 7024 31074
rect 7076 30988 7088 31074
rect 7012 30932 7022 30988
rect 7078 30932 7088 30988
rect 2776 30790 2786 30846
rect 2842 30790 2852 30846
rect 2776 30704 2788 30790
rect 2840 30704 2852 30790
rect 2776 30648 2786 30704
rect 2842 30648 2852 30704
rect 2776 30562 2788 30648
rect 2840 30562 2852 30648
rect 2776 30506 2786 30562
rect 2842 30506 2852 30562
rect 2776 30454 2788 30506
rect 2840 30454 2852 30506
rect 3020 30858 4243 30870
rect 3020 30494 3032 30858
rect 3084 30770 4243 30858
rect 3084 30494 3096 30770
rect 3020 30482 3096 30494
rect 3496 30678 3596 30690
rect 2776 30442 2852 30454
rect 165 28567 586 28632
rect 165 28511 175 28567
rect 231 28511 317 28567
rect 373 28511 586 28567
rect 165 28425 586 28511
rect 165 28369 175 28425
rect 231 28369 317 28425
rect 373 28369 586 28425
rect 1007 28401 1107 30101
rect 1688 30021 1788 30314
rect 3496 30314 3520 30678
rect 3572 30314 3596 30678
rect 1985 30109 3339 30119
rect 1985 30053 1995 30109
rect 2051 30107 2137 30109
rect 2193 30107 2279 30109
rect 2335 30107 2421 30109
rect 2477 30107 2563 30109
rect 2619 30107 2705 30109
rect 2761 30107 2847 30109
rect 2903 30107 2989 30109
rect 3045 30107 3131 30109
rect 3187 30107 3273 30109
rect 2051 30053 2137 30055
rect 2193 30053 2279 30055
rect 2335 30053 2421 30055
rect 2477 30053 2563 30055
rect 2619 30053 2705 30055
rect 2761 30053 2847 30055
rect 2903 30053 2989 30055
rect 3045 30053 3131 30055
rect 3187 30053 3273 30055
rect 3329 30053 3339 30109
rect 1985 30043 3339 30053
rect 1187 29921 1788 30021
rect 1187 28401 1287 29921
rect 1367 29817 1547 29829
rect 1367 29765 1379 29817
rect 1535 29765 1547 29817
rect 1367 29753 1547 29765
rect 1367 28401 1467 29753
rect 1547 29637 1727 29649
rect 1547 29585 1559 29637
rect 1715 29585 1727 29637
rect 1547 29573 1727 29585
rect 1547 28401 1655 29573
rect 3496 29442 3596 30314
rect 4143 29469 4243 30770
rect 4472 30858 6002 30870
rect 4472 30494 4484 30858
rect 4536 30770 6002 30858
rect 4536 30494 4548 30770
rect 4472 30482 4548 30494
rect 4948 30678 5048 30690
rect 3496 29430 3676 29442
rect 3496 29378 3508 29430
rect 3664 29378 3676 29430
rect 3496 29366 3676 29378
rect 4143 29313 4167 29469
rect 4219 29313 4243 29469
rect 4143 29301 4243 29313
rect 4948 30314 4972 30678
rect 5024 30314 5048 30678
rect 4948 29469 5048 30314
rect 4948 29313 4972 29469
rect 5024 29313 5048 29469
rect 4948 29301 5048 29313
rect 5902 29469 6002 30770
rect 7012 30846 7024 30932
rect 7076 30846 7088 30932
rect 7012 30790 7022 30846
rect 7078 30790 7088 30846
rect 7012 30704 7024 30790
rect 7076 30704 7088 30790
rect 6512 30678 6612 30690
rect 6512 30314 6536 30678
rect 6588 30314 6612 30678
rect 6512 29829 6612 30314
rect 6432 29817 6612 29829
rect 6432 29765 6444 29817
rect 6600 29765 6612 29817
rect 6432 29753 6612 29765
rect 6756 30678 6856 30690
rect 6756 30314 6780 30678
rect 6832 30314 6856 30678
rect 7012 30648 7022 30704
rect 7078 30648 7088 30704
rect 7012 30562 7024 30648
rect 7076 30562 7088 30648
rect 7012 30506 7022 30562
rect 7078 30506 7088 30562
rect 7012 30454 7024 30506
rect 7076 30454 7088 30506
rect 7012 30442 7088 30454
rect 6756 29649 6856 30314
rect 6676 29637 6856 29649
rect 6676 29585 6688 29637
rect 6844 29585 6856 29637
rect 6676 29573 6856 29585
rect 5902 29313 5926 29469
rect 5978 29313 6002 29469
rect 5902 29301 6002 29313
rect 165 28283 586 28369
rect 165 28227 175 28283
rect 231 28227 317 28283
rect 373 28227 586 28283
rect 165 28141 586 28227
rect 165 28085 175 28141
rect 231 28085 317 28141
rect 373 28085 586 28141
rect 165 27999 586 28085
rect 7332 28015 7732 41648
rect 11017 40972 11093 44770
rect 12406 44053 12624 44065
rect 12406 44001 12434 44053
rect 12590 44001 12624 44053
rect 11426 41815 11658 41827
rect 11426 41659 11583 41815
rect 11635 41659 11658 41815
rect 11426 41647 11658 41659
rect 11017 40816 11029 40972
rect 11081 40816 11093 40972
rect 11017 40804 11093 40816
rect 11200 41163 11362 41175
rect 11200 41007 11298 41163
rect 11350 41007 11362 41163
rect 11200 40995 11362 41007
rect 11426 41080 11502 41647
rect 11571 41341 12060 41353
rect 11571 41185 11583 41341
rect 11635 41185 12060 41341
rect 11571 41173 12060 41185
rect 11426 41004 11596 41080
rect 10888 40734 11068 40746
rect 10888 40682 10900 40734
rect 11056 40682 11068 40734
rect 10888 40670 11068 40682
rect 10644 40462 10824 40474
rect 10644 40410 10656 40462
rect 10812 40410 10824 40462
rect 10644 40398 10824 40410
rect 7888 40316 9767 40326
rect 7888 40314 7997 40316
rect 8053 40314 8139 40316
rect 8195 40314 8281 40316
rect 8337 40314 8423 40316
rect 8479 40314 8565 40316
rect 8621 40314 8707 40316
rect 8763 40314 8849 40316
rect 8905 40314 8991 40316
rect 9047 40314 9133 40316
rect 9189 40314 9275 40316
rect 9331 40314 9417 40316
rect 9473 40314 9559 40316
rect 9615 40314 9701 40316
rect 7888 40262 7900 40314
rect 7888 40260 7997 40262
rect 8053 40260 8139 40262
rect 8195 40260 8281 40262
rect 8337 40260 8423 40262
rect 8479 40260 8565 40262
rect 8621 40260 8707 40262
rect 8763 40260 8849 40262
rect 8905 40260 8991 40262
rect 9047 40260 9133 40262
rect 9189 40260 9275 40262
rect 9331 40260 9417 40262
rect 9473 40260 9559 40262
rect 9615 40260 9701 40262
rect 9757 40260 9767 40316
rect 7888 40250 9767 40260
rect 10327 39788 10403 39800
rect 10327 39760 10339 39788
rect 10391 39760 10403 39788
rect 10327 39704 10337 39760
rect 10393 39704 10403 39760
rect 10327 39618 10339 39704
rect 10391 39618 10403 39704
rect 10327 39562 10337 39618
rect 10393 39562 10403 39618
rect 10327 39476 10339 39562
rect 10391 39476 10403 39562
rect 10327 39420 10337 39476
rect 10393 39420 10403 39476
rect 10327 39334 10339 39420
rect 10391 39334 10403 39420
rect 10327 39278 10337 39334
rect 10393 39278 10403 39334
rect 10327 39192 10339 39278
rect 10391 39192 10403 39278
rect 10327 39136 10337 39192
rect 10393 39136 10403 39192
rect 10327 39050 10339 39136
rect 10391 39050 10403 39136
rect 10327 38994 10337 39050
rect 10393 38994 10403 39050
rect 10327 38908 10339 38994
rect 10391 38908 10403 38994
rect 10327 38852 10337 38908
rect 10393 38852 10403 38908
rect 10644 39046 10720 40398
rect 10644 38890 10656 39046
rect 10708 38890 10720 39046
rect 10644 38878 10720 38890
rect 10888 39046 10964 40670
rect 10888 38890 10900 39046
rect 10952 38890 10964 39046
rect 10888 38878 10964 38890
rect 11200 39788 11276 40995
rect 11520 40610 11596 41004
rect 11416 40598 11596 40610
rect 11416 40546 11428 40598
rect 11584 40546 11596 40598
rect 11416 40534 11596 40546
rect 11200 39760 11212 39788
rect 11264 39760 11276 39788
rect 11200 39704 11210 39760
rect 11266 39704 11276 39760
rect 11200 39618 11212 39704
rect 11264 39618 11276 39704
rect 11200 39562 11210 39618
rect 11266 39562 11276 39618
rect 11200 39476 11212 39562
rect 11264 39476 11276 39562
rect 11200 39420 11210 39476
rect 11266 39420 11276 39476
rect 11200 39334 11212 39420
rect 11264 39334 11276 39420
rect 11200 39278 11210 39334
rect 11266 39278 11276 39334
rect 11200 39192 11212 39278
rect 11264 39192 11276 39278
rect 11200 39136 11210 39192
rect 11266 39136 11276 39192
rect 11200 39050 11212 39136
rect 11264 39050 11276 39136
rect 11200 38994 11210 39050
rect 11266 38994 11276 39050
rect 11200 38908 11212 38994
rect 11264 38908 11276 38994
rect 10327 38800 10339 38852
rect 10391 38800 10403 38852
rect 10327 38766 10403 38800
rect 10327 38710 10337 38766
rect 10393 38710 10403 38766
rect 10327 38700 10403 38710
rect 11200 38852 11210 38908
rect 11266 38852 11276 38908
rect 11200 38800 11212 38852
rect 11264 38800 11276 38852
rect 11200 38766 11276 38800
rect 11200 38710 11210 38766
rect 11266 38710 11276 38766
rect 11200 38700 11276 38710
rect 8293 38688 8369 38700
rect 8293 38532 8305 38688
rect 8357 38532 8369 38688
rect 8293 36774 8369 38532
rect 11520 38685 11596 40534
rect 11520 38529 11532 38685
rect 11584 38529 11596 38685
rect 8671 38512 8747 38524
rect 11520 38517 11596 38529
rect 11690 40883 11890 40910
rect 11690 40831 11714 40883
rect 11870 40831 11890 40883
rect 8439 37939 8515 37951
rect 8439 37783 8451 37939
rect 8503 37783 8515 37939
rect 8439 37002 8515 37783
rect 8439 36846 8451 37002
rect 8503 36846 8515 37002
rect 8439 36834 8515 36846
rect 8671 37524 8683 38512
rect 8735 37524 8747 38512
rect 8895 37939 9566 37951
rect 8895 37783 8907 37939
rect 8959 37783 9566 37939
rect 8895 37771 9566 37783
rect 8293 36762 8473 36774
rect 8293 36710 8305 36762
rect 8461 36710 8473 36762
rect 8293 36698 8473 36710
rect 8318 36218 8498 36230
rect 8318 36166 8330 36218
rect 8486 36166 8498 36218
rect 8318 36154 8498 36166
rect 8318 32888 8394 36154
rect 8671 35982 8747 37524
rect 8970 36626 9150 36638
rect 8970 36574 8982 36626
rect 9138 36574 9150 36626
rect 8970 36562 9150 36574
rect 8671 35958 8681 35982
rect 8567 35946 8681 35958
rect 8567 35894 8579 35946
rect 8737 35926 8747 35982
rect 8735 35894 8747 35926
rect 8567 35882 8747 35894
rect 8671 35840 8747 35882
rect 8671 35784 8681 35840
rect 8737 35784 8747 35840
rect 8671 35698 8747 35784
rect 8671 35642 8681 35698
rect 8737 35642 8747 35698
rect 8671 35556 8747 35642
rect 8671 35500 8681 35556
rect 8737 35500 8747 35556
rect 8671 35414 8747 35500
rect 8671 35358 8681 35414
rect 8737 35358 8747 35414
rect 8671 35272 8747 35358
rect 8671 35216 8681 35272
rect 8737 35216 8747 35272
rect 8671 35130 8747 35216
rect 8671 35074 8681 35130
rect 8737 35074 8747 35130
rect 8671 34988 8747 35074
rect 8671 34932 8681 34988
rect 8737 34932 8747 34988
rect 8671 34846 8747 34932
rect 8671 34790 8681 34846
rect 8737 34790 8747 34846
rect 8671 34704 8747 34790
rect 8671 34648 8681 34704
rect 8737 34648 8747 34704
rect 8671 34562 8747 34648
rect 8671 34506 8681 34562
rect 8737 34506 8747 34562
rect 8671 34496 8747 34506
rect 8830 36490 9010 36502
rect 8830 36438 8842 36490
rect 8998 36438 9010 36490
rect 8830 36426 9010 36438
rect 8830 34435 8906 36426
rect 8830 34279 8842 34435
rect 8894 34279 8906 34435
rect 8830 34267 8906 34279
rect 9074 34435 9150 36562
rect 9074 34279 9086 34435
rect 9138 34279 9150 34435
rect 9074 34267 9150 34279
rect 9490 36366 9566 37771
rect 11690 37712 11890 40831
rect 11984 40474 12060 41173
rect 11984 40462 12164 40474
rect 11984 40410 11996 40462
rect 12152 40410 12164 40462
rect 11984 40398 12164 40410
rect 12406 38160 12624 44001
rect 13096 42968 13608 42996
rect 13096 42912 13191 42968
rect 13247 42912 13303 42968
rect 13359 42912 13415 42968
rect 13471 42912 13608 42968
rect 13096 42868 13608 42912
rect 13096 42712 13108 42868
rect 13160 42856 13544 42868
rect 13160 42800 13191 42856
rect 13247 42800 13303 42856
rect 13359 42800 13415 42856
rect 13471 42800 13544 42856
rect 13160 42744 13544 42800
rect 13160 42712 13191 42744
rect 13096 42688 13191 42712
rect 13247 42688 13303 42744
rect 13359 42688 13415 42744
rect 13471 42712 13544 42744
rect 13596 42712 13608 42868
rect 13471 42688 13608 42712
rect 13096 42632 13608 42688
rect 13096 42576 13191 42632
rect 13247 42576 13303 42632
rect 13359 42576 13415 42632
rect 13471 42576 13608 42632
rect 13096 42520 13608 42576
rect 13096 42464 13191 42520
rect 13247 42464 13303 42520
rect 13359 42464 13415 42520
rect 13471 42464 13608 42520
rect 13096 42408 13608 42464
rect 13096 42352 13191 42408
rect 13247 42352 13303 42408
rect 13359 42352 13415 42408
rect 13471 42352 13608 42408
rect 13096 42296 13608 42352
rect 13096 42240 13191 42296
rect 13247 42240 13303 42296
rect 13359 42240 13415 42296
rect 13471 42240 13608 42296
rect 13096 42184 13608 42240
rect 13096 42128 13191 42184
rect 13247 42128 13303 42184
rect 13359 42128 13415 42184
rect 13471 42128 13608 42184
rect 13096 42072 13608 42128
rect 13096 42016 13191 42072
rect 13247 42016 13303 42072
rect 13359 42016 13415 42072
rect 13471 42016 13608 42072
rect 13096 41960 13608 42016
rect 13096 41941 13191 41960
rect 13096 41785 13108 41941
rect 13160 41904 13191 41941
rect 13247 41904 13303 41960
rect 13359 41904 13415 41960
rect 13471 41941 13608 41960
rect 13471 41904 13544 41941
rect 13160 41848 13544 41904
rect 13160 41792 13191 41848
rect 13247 41792 13303 41848
rect 13359 41792 13415 41848
rect 13471 41792 13544 41848
rect 13160 41785 13544 41792
rect 13596 41785 13608 41941
rect 13096 41773 13608 41785
rect 13766 40610 13842 57263
rect 13662 40598 13842 40610
rect 13662 40546 13674 40598
rect 13830 40546 13842 40598
rect 13662 40534 13842 40546
rect 13912 40474 13988 57263
rect 14058 40838 14134 57263
rect 14204 51352 14280 57600
rect 14380 56715 14780 56747
rect 14380 56559 14392 56715
rect 14548 56559 14780 56715
rect 14380 55767 14780 56559
rect 14380 55711 14410 55767
rect 14466 55711 14552 55767
rect 14608 55711 14694 55767
rect 14750 55711 14780 55767
rect 14380 55625 14780 55711
rect 14380 55569 14410 55625
rect 14466 55569 14552 55625
rect 14608 55569 14694 55625
rect 14750 55569 14780 55625
rect 14380 55483 14780 55569
rect 14380 55427 14410 55483
rect 14466 55427 14552 55483
rect 14608 55427 14694 55483
rect 14750 55427 14780 55483
rect 14380 55341 14780 55427
rect 14380 55285 14410 55341
rect 14466 55285 14552 55341
rect 14608 55285 14694 55341
rect 14750 55285 14780 55341
rect 14380 55199 14780 55285
rect 14380 55143 14410 55199
rect 14466 55143 14552 55199
rect 14608 55143 14694 55199
rect 14750 55143 14780 55199
rect 14380 55057 14780 55143
rect 14380 55001 14410 55057
rect 14466 55001 14552 55057
rect 14608 55001 14694 55057
rect 14750 55001 14780 55057
rect 14380 54915 14780 55001
rect 14380 54859 14410 54915
rect 14466 54859 14552 54915
rect 14608 54859 14694 54915
rect 14750 54859 14780 54915
rect 14380 54773 14780 54859
rect 14380 54717 14410 54773
rect 14466 54717 14552 54773
rect 14608 54717 14694 54773
rect 14750 54717 14780 54773
rect 14380 54631 14780 54717
rect 14380 54575 14410 54631
rect 14466 54575 14552 54631
rect 14608 54575 14694 54631
rect 14750 54575 14780 54631
rect 14380 54489 14780 54575
rect 14380 54433 14410 54489
rect 14466 54433 14552 54489
rect 14608 54433 14694 54489
rect 14750 54433 14780 54489
rect 14204 45993 14280 49606
rect 14204 45837 14216 45993
rect 14268 45837 14280 45993
rect 14204 45825 14280 45837
rect 14380 49304 14780 54433
rect 14942 52491 15032 52600
rect 14942 52489 14954 52491
rect 15006 52489 15032 52491
rect 14942 52433 14952 52489
rect 15008 52433 15032 52489
rect 14942 52347 14954 52433
rect 15006 52347 15032 52433
rect 14942 52291 14952 52347
rect 15008 52291 15032 52347
rect 14942 52205 14954 52291
rect 15006 52205 15032 52291
rect 14942 52149 14952 52205
rect 15008 52149 15032 52205
rect 14942 52063 14954 52149
rect 15006 52063 15032 52149
rect 14942 52007 14952 52063
rect 15008 52007 15032 52063
rect 14942 51921 14954 52007
rect 15006 51921 15032 52007
rect 14942 51865 14952 51921
rect 15008 51865 15032 51921
rect 14942 51779 14954 51865
rect 15006 51779 15032 51865
rect 14942 51723 14952 51779
rect 15008 51723 15032 51779
rect 14942 51637 14954 51723
rect 15006 51637 15032 51723
rect 14942 51581 14952 51637
rect 15008 51581 15032 51637
rect 14942 51495 14954 51581
rect 15006 51495 15032 51581
rect 14942 51439 14952 51495
rect 15008 51439 15032 51495
rect 14942 51353 14954 51439
rect 15006 51353 15032 51439
rect 14942 51297 14952 51353
rect 15008 51297 15032 51353
rect 14942 51295 14954 51297
rect 15006 51295 15032 51297
rect 14942 51200 15032 51295
rect 14380 49252 14392 49304
rect 14444 49252 14500 49304
rect 14552 49252 14780 49304
rect 14380 49196 14780 49252
rect 14380 49144 14392 49196
rect 14444 49144 14500 49196
rect 14552 49144 14780 49196
rect 14380 49088 14780 49144
rect 14380 49036 14392 49088
rect 14444 49036 14500 49088
rect 14552 49036 14780 49088
rect 14380 48980 14780 49036
rect 14380 48928 14392 48980
rect 14444 48928 14500 48980
rect 14552 48928 14780 48980
rect 14380 48872 14780 48928
rect 14380 48820 14392 48872
rect 14444 48820 14500 48872
rect 14552 48820 14780 48872
rect 14380 48336 14780 48820
rect 14380 48284 14392 48336
rect 14444 48284 14500 48336
rect 14552 48284 14780 48336
rect 14380 48228 14780 48284
rect 14380 48176 14392 48228
rect 14444 48176 14500 48228
rect 14552 48176 14780 48228
rect 14380 48120 14780 48176
rect 14380 48068 14392 48120
rect 14444 48068 14500 48120
rect 14552 48068 14780 48120
rect 14380 48012 14780 48068
rect 14380 47960 14392 48012
rect 14444 47960 14500 48012
rect 14552 47960 14780 48012
rect 14380 47904 14780 47960
rect 14380 47852 14392 47904
rect 14444 47852 14500 47904
rect 14552 47852 14780 47904
rect 14380 47760 14780 47852
rect 14380 47704 14410 47760
rect 14466 47704 14552 47760
rect 14608 47704 14694 47760
rect 14750 47704 14780 47760
rect 14380 47618 14780 47704
rect 14380 47562 14410 47618
rect 14466 47562 14552 47618
rect 14608 47562 14694 47618
rect 14750 47562 14780 47618
rect 14380 47476 14780 47562
rect 14380 47420 14410 47476
rect 14466 47420 14552 47476
rect 14608 47420 14694 47476
rect 14750 47420 14780 47476
rect 14380 47334 14780 47420
rect 14380 47278 14410 47334
rect 14466 47278 14552 47334
rect 14608 47278 14694 47334
rect 14750 47278 14780 47334
rect 14380 47192 14780 47278
rect 14380 47136 14410 47192
rect 14466 47136 14552 47192
rect 14608 47136 14694 47192
rect 14750 47136 14780 47192
rect 14380 47050 14780 47136
rect 14380 46994 14410 47050
rect 14466 46994 14552 47050
rect 14608 46994 14694 47050
rect 14750 46994 14780 47050
rect 14380 46908 14780 46994
rect 14380 46852 14410 46908
rect 14466 46852 14552 46908
rect 14608 46852 14694 46908
rect 14750 46852 14780 46908
rect 14380 46766 14780 46852
rect 14380 46710 14410 46766
rect 14466 46710 14552 46766
rect 14608 46710 14694 46766
rect 14750 46710 14780 46766
rect 14380 46624 14780 46710
rect 14380 46568 14410 46624
rect 14466 46568 14552 46624
rect 14608 46568 14694 46624
rect 14750 46568 14780 46624
rect 14380 46482 14780 46568
rect 14380 46426 14410 46482
rect 14466 46426 14552 46482
rect 14608 46426 14694 46482
rect 14750 46426 14780 46482
rect 14058 40682 14070 40838
rect 14122 40682 14134 40838
rect 14058 40670 14134 40682
rect 14380 41360 14780 46426
rect 14380 41304 14410 41360
rect 14466 41304 14552 41360
rect 14608 41304 14694 41360
rect 14750 41304 14780 41360
rect 14380 41218 14780 41304
rect 14380 41162 14410 41218
rect 14466 41162 14552 41218
rect 14608 41162 14694 41218
rect 14750 41162 14780 41218
rect 14380 41076 14780 41162
rect 14380 41020 14410 41076
rect 14466 41020 14552 41076
rect 14608 41020 14694 41076
rect 14750 41020 14780 41076
rect 14380 40934 14780 41020
rect 14380 40878 14410 40934
rect 14466 40878 14552 40934
rect 14608 40878 14694 40934
rect 14750 40878 14780 40934
rect 14380 40792 14780 40878
rect 14380 40736 14410 40792
rect 14466 40736 14552 40792
rect 14608 40736 14694 40792
rect 14750 40736 14780 40792
rect 13808 40462 13988 40474
rect 13808 40410 13820 40462
rect 13976 40410 13988 40462
rect 13808 40398 13988 40410
rect 14380 40650 14780 40736
rect 14380 40594 14410 40650
rect 14466 40594 14552 40650
rect 14608 40594 14694 40650
rect 14750 40594 14780 40650
rect 14380 40508 14780 40594
rect 14380 40452 14410 40508
rect 14466 40452 14552 40508
rect 14608 40452 14694 40508
rect 14750 40452 14780 40508
rect 14380 40366 14780 40452
rect 12748 40316 13818 40326
rect 12748 40260 12758 40316
rect 12814 40314 12900 40316
rect 12956 40314 13042 40316
rect 13098 40314 13184 40316
rect 13240 40314 13326 40316
rect 13382 40314 13468 40316
rect 13524 40314 13610 40316
rect 13666 40314 13752 40316
rect 12814 40260 12900 40262
rect 12956 40260 13042 40262
rect 13098 40260 13184 40262
rect 13240 40260 13326 40262
rect 13382 40260 13468 40262
rect 13524 40260 13610 40262
rect 13666 40260 13752 40262
rect 13808 40260 13818 40316
rect 12748 40250 13818 40260
rect 14380 40310 14410 40366
rect 14466 40310 14552 40366
rect 14608 40310 14694 40366
rect 14750 40310 14780 40366
rect 14380 40224 14780 40310
rect 14380 40168 14410 40224
rect 14466 40168 14552 40224
rect 14608 40168 14694 40224
rect 14750 40168 14780 40224
rect 14380 40082 14780 40168
rect 14380 40026 14410 40082
rect 14466 40026 14552 40082
rect 14608 40026 14694 40082
rect 14750 40026 14780 40082
rect 13303 38675 13754 38687
rect 13303 38519 13315 38675
rect 13367 38519 13754 38675
rect 13303 38507 13754 38519
rect 12406 38104 12416 38160
rect 12472 38104 12558 38160
rect 12614 38104 12624 38160
rect 12406 38018 12624 38104
rect 12406 37962 12416 38018
rect 12472 37962 12558 38018
rect 12614 37962 12624 38018
rect 12406 37876 12624 37962
rect 12406 37820 12416 37876
rect 12472 37820 12558 37876
rect 12614 37820 12624 37876
rect 12406 37734 12624 37820
rect 10331 37570 11551 37580
rect 10331 37568 10435 37570
rect 10491 37568 10577 37570
rect 10633 37568 10719 37570
rect 10775 37568 10861 37570
rect 10917 37568 11003 37570
rect 11059 37568 11145 37570
rect 11201 37568 11287 37570
rect 11343 37568 11429 37570
rect 11485 37568 11551 37570
rect 10331 37516 10343 37568
rect 11539 37516 11551 37568
rect 10331 37514 10435 37516
rect 10491 37514 10577 37516
rect 10633 37514 10719 37516
rect 10775 37514 10861 37516
rect 10917 37514 11003 37516
rect 11059 37514 11145 37516
rect 11201 37514 11287 37516
rect 11343 37514 11429 37516
rect 11485 37514 11551 37516
rect 10331 37504 11551 37514
rect 11690 37512 12090 37712
rect 9490 36354 9670 36366
rect 9490 36302 9502 36354
rect 9658 36302 9670 36354
rect 9490 36290 9670 36302
rect 9490 34435 9566 36290
rect 10394 36082 10574 36094
rect 10394 36030 10406 36082
rect 10562 36030 10574 36082
rect 10394 36018 10574 36030
rect 10998 36086 11074 36096
rect 10998 36030 11008 36086
rect 11064 36030 11074 36086
rect 10100 35982 10176 35992
rect 10100 35926 10110 35982
rect 10166 35926 10176 35982
rect 10100 35840 10112 35926
rect 10164 35840 10176 35926
rect 10100 35784 10110 35840
rect 10166 35784 10176 35840
rect 10100 35698 10112 35784
rect 10164 35698 10176 35784
rect 10100 35642 10110 35698
rect 10166 35642 10176 35698
rect 10100 35556 10112 35642
rect 10164 35556 10176 35642
rect 10100 35500 10110 35556
rect 10166 35500 10176 35556
rect 10100 35414 10112 35500
rect 10164 35414 10176 35500
rect 10100 35358 10110 35414
rect 10166 35358 10176 35414
rect 10100 35272 10112 35358
rect 10164 35272 10176 35358
rect 10100 35216 10110 35272
rect 10166 35216 10176 35272
rect 10100 35130 10112 35216
rect 10164 35130 10176 35216
rect 10100 35074 10110 35130
rect 10166 35074 10176 35130
rect 10100 34988 10112 35074
rect 10164 34988 10176 35074
rect 10100 34932 10110 34988
rect 10166 34932 10176 34988
rect 10100 34846 10112 34932
rect 10164 34846 10176 34932
rect 10100 34790 10110 34846
rect 10166 34790 10176 34846
rect 10100 34704 10112 34790
rect 10164 34704 10176 34790
rect 10100 34648 10110 34704
rect 10166 34648 10176 34704
rect 10100 34562 10112 34648
rect 10164 34562 10176 34648
rect 10100 34506 10110 34562
rect 10166 34506 10176 34562
rect 10100 34496 10176 34506
rect 9490 34279 9502 34435
rect 9554 34279 9566 34435
rect 9490 34267 9566 34279
rect 10394 34267 10470 36018
rect 10998 35946 11074 36030
rect 11498 36082 11678 36094
rect 11498 36030 11510 36082
rect 11666 36030 11678 36082
rect 11498 36018 11678 36030
rect 10998 35944 11010 35946
rect 11062 35944 11074 35946
rect 10998 35888 11008 35944
rect 11064 35888 11074 35944
rect 10998 35802 11010 35888
rect 11062 35802 11074 35888
rect 10998 35746 11008 35802
rect 11064 35746 11074 35802
rect 10998 35660 11010 35746
rect 11062 35660 11074 35746
rect 10998 35604 11008 35660
rect 11064 35604 11074 35660
rect 10998 35518 11010 35604
rect 11062 35518 11074 35604
rect 10998 35462 11008 35518
rect 11064 35462 11074 35518
rect 10998 35376 11010 35462
rect 11062 35376 11074 35462
rect 10998 35320 11008 35376
rect 11064 35320 11074 35376
rect 10998 35234 11010 35320
rect 11062 35234 11074 35320
rect 10998 35178 11008 35234
rect 11064 35178 11074 35234
rect 10998 35092 11010 35178
rect 11062 35092 11074 35178
rect 10998 35036 11008 35092
rect 11064 35036 11074 35092
rect 10998 34950 11010 35036
rect 11062 34950 11074 35036
rect 10998 34894 11008 34950
rect 11064 34894 11074 34950
rect 10998 34808 11010 34894
rect 11062 34808 11074 34894
rect 10998 34752 11008 34808
rect 11064 34752 11074 34808
rect 10998 34666 11010 34752
rect 11062 34666 11074 34752
rect 10998 34610 11008 34666
rect 11064 34610 11074 34666
rect 10998 34524 11010 34610
rect 11062 34524 11074 34610
rect 10998 34468 11008 34524
rect 11064 34468 11074 34524
rect 10998 34382 11010 34468
rect 11062 34382 11074 34468
rect 10998 34326 11008 34382
rect 11064 34326 11074 34382
rect 10998 34240 11010 34326
rect 11062 34240 11074 34326
rect 11602 34267 11678 36018
rect 11890 35982 12090 37512
rect 12406 37678 12416 37734
rect 12472 37678 12558 37734
rect 12614 37678 12624 37734
rect 12406 37592 12624 37678
rect 12406 37536 12416 37592
rect 12472 37536 12558 37592
rect 12614 37536 12624 37592
rect 12406 37450 12624 37536
rect 12406 37394 12416 37450
rect 12472 37394 12558 37450
rect 12614 37394 12624 37450
rect 12406 37308 12624 37394
rect 12406 37252 12416 37308
rect 12472 37252 12558 37308
rect 12614 37252 12624 37308
rect 12406 37166 12624 37252
rect 12406 37110 12416 37166
rect 12472 37110 12558 37166
rect 12614 37110 12624 37166
rect 12406 37024 12624 37110
rect 12406 36968 12416 37024
rect 12472 36968 12558 37024
rect 12614 36968 12624 37024
rect 12406 36882 12624 36968
rect 13439 38023 13515 38035
rect 13439 37867 13451 38023
rect 13503 37867 13515 38023
rect 12406 36826 12416 36882
rect 12472 36826 12558 36882
rect 12614 36826 12624 36882
rect 13062 36898 13242 36910
rect 13062 36846 13074 36898
rect 13230 36846 13242 36898
rect 13062 36834 13242 36846
rect 12406 36800 12624 36826
rect 12922 36762 13102 36774
rect 12922 36710 12934 36762
rect 13090 36710 13102 36762
rect 12922 36698 13102 36710
rect 11890 35926 11906 35982
rect 11962 35926 12090 35982
rect 11890 35840 11908 35926
rect 11960 35840 12090 35926
rect 11890 35784 11906 35840
rect 11962 35784 12090 35840
rect 11890 35698 11908 35784
rect 11960 35698 12090 35784
rect 11890 35642 11906 35698
rect 11962 35642 12090 35698
rect 11890 35556 11908 35642
rect 11960 35556 12090 35642
rect 11890 35500 11906 35556
rect 11962 35500 12090 35556
rect 11890 35414 11908 35500
rect 11960 35414 12090 35500
rect 11890 35358 11906 35414
rect 11962 35358 12090 35414
rect 11890 35272 11908 35358
rect 11960 35272 12090 35358
rect 11890 35216 11906 35272
rect 11962 35216 12090 35272
rect 11890 35130 11908 35216
rect 11960 35130 12090 35216
rect 11890 35074 11906 35130
rect 11962 35074 12090 35130
rect 11890 34988 11908 35074
rect 11960 34988 12090 35074
rect 11890 34932 11906 34988
rect 11962 34932 12090 34988
rect 11890 34846 11908 34932
rect 11960 34846 12090 34932
rect 11890 34790 11906 34846
rect 11962 34790 12090 34846
rect 11890 34704 11908 34790
rect 11960 34704 12090 34790
rect 11890 34648 11906 34704
rect 11962 34648 12090 34704
rect 11890 34562 11908 34648
rect 11960 34562 12090 34648
rect 11890 34506 11906 34562
rect 11962 34506 12090 34562
rect 11890 34499 12090 34506
rect 12506 36354 12686 36366
rect 12506 36302 12518 36354
rect 12674 36302 12686 36354
rect 12506 36290 12686 36302
rect 11896 34496 11972 34499
rect 12506 34435 12582 36290
rect 12506 34279 12518 34435
rect 12570 34279 12582 34435
rect 12506 34267 12582 34279
rect 12922 34435 12998 36698
rect 12922 34279 12934 34435
rect 12986 34279 12998 34435
rect 12922 34267 12998 34279
rect 13166 34435 13242 36834
rect 13439 36094 13515 37867
rect 13678 36230 13754 38507
rect 13574 36218 13754 36230
rect 13574 36166 13586 36218
rect 13742 36166 13754 36218
rect 13574 36154 13754 36166
rect 13335 36082 13515 36094
rect 13335 36030 13347 36082
rect 13503 36030 13515 36082
rect 13335 36018 13515 36030
rect 13166 34279 13178 34435
rect 13230 34279 13242 34435
rect 13166 34267 13242 34279
rect 10998 34184 11008 34240
rect 11064 34184 11074 34240
rect 10998 34098 11010 34184
rect 11062 34098 11074 34184
rect 10998 34042 11008 34098
rect 11064 34042 11074 34098
rect 10998 33956 11010 34042
rect 11062 33956 11074 34042
rect 10998 33900 11008 33956
rect 11064 33900 11074 33956
rect 10998 33814 11010 33900
rect 11062 33814 11074 33900
rect 10998 33758 11008 33814
rect 11064 33758 11074 33814
rect 10998 33672 11010 33758
rect 11062 33672 11074 33758
rect 10998 33616 11008 33672
rect 11064 33616 11074 33672
rect 10998 33294 11010 33616
rect 11062 33294 11074 33616
rect 10998 33282 11074 33294
rect 10998 32905 11074 32915
rect 10998 32849 11008 32905
rect 11064 32849 11074 32905
rect 13678 32888 13754 36154
rect 14380 33851 14780 40026
rect 14942 38160 15032 38200
rect 14942 38104 14952 38160
rect 15008 38104 15032 38160
rect 14942 38018 14954 38104
rect 15006 38018 15032 38104
rect 14942 37962 14952 38018
rect 15008 37962 15032 38018
rect 14942 37876 14954 37962
rect 15006 37876 15032 37962
rect 14942 37820 14952 37876
rect 15008 37820 15032 37876
rect 14942 37734 14954 37820
rect 15006 37734 15032 37820
rect 14942 37678 14952 37734
rect 15008 37678 15032 37734
rect 14942 37592 14954 37678
rect 15006 37592 15032 37678
rect 14942 37536 14952 37592
rect 15008 37536 15032 37592
rect 14942 37450 14954 37536
rect 15006 37450 15032 37536
rect 14942 37394 14952 37450
rect 15008 37394 15032 37450
rect 14942 37308 14954 37394
rect 15006 37308 15032 37394
rect 14942 37252 14952 37308
rect 15008 37252 15032 37308
rect 14942 37166 14954 37252
rect 15006 37166 15032 37252
rect 14942 37110 14952 37166
rect 15008 37110 15032 37166
rect 14942 37024 14954 37110
rect 15006 37024 15032 37110
rect 14942 36968 14952 37024
rect 15008 36968 15032 37024
rect 14942 36882 14954 36968
rect 15006 36882 15032 36968
rect 14942 36826 14952 36882
rect 15008 36826 15032 36882
rect 14942 36800 15032 36826
rect 14380 33348 14514 33851
rect 14566 33348 14780 33851
rect 14380 33292 14410 33348
rect 14466 33292 14514 33348
rect 14608 33292 14694 33348
rect 14750 33292 14780 33348
rect 14380 33206 14514 33292
rect 14566 33206 14780 33292
rect 14380 33150 14410 33206
rect 14466 33150 14514 33206
rect 14608 33150 14694 33206
rect 14750 33150 14780 33206
rect 14380 33064 14514 33150
rect 14566 33064 14780 33150
rect 14380 33008 14410 33064
rect 14466 33008 14514 33064
rect 14608 33008 14694 33064
rect 14750 33008 14780 33064
rect 14380 32922 14514 33008
rect 14566 32922 14780 33008
rect 10998 32825 11074 32849
rect 10998 32763 11010 32825
rect 11062 32763 11074 32825
rect 10998 32707 11008 32763
rect 11064 32707 11074 32763
rect 7976 32692 8052 32702
rect 7976 32636 7986 32692
rect 8042 32636 8052 32692
rect 7976 32550 7988 32636
rect 8040 32550 8052 32636
rect 7976 32494 7986 32550
rect 8042 32494 8052 32550
rect 7976 32408 7988 32494
rect 8040 32408 8052 32494
rect 7976 32352 7986 32408
rect 8042 32352 8052 32408
rect 7976 32266 7988 32352
rect 8040 32266 8052 32352
rect 7976 32210 7986 32266
rect 8042 32210 8052 32266
rect 7976 32124 7988 32210
rect 8040 32124 8052 32210
rect 7976 32068 7986 32124
rect 8042 32068 8052 32124
rect 7976 31982 7988 32068
rect 8040 31982 8052 32068
rect 7976 31926 7986 31982
rect 8042 31926 8052 31982
rect 7976 31840 7988 31926
rect 8040 31840 8052 31926
rect 7976 31784 7986 31840
rect 8042 31784 8052 31840
rect 7976 31698 7988 31784
rect 8040 31698 8052 31784
rect 7976 31642 7986 31698
rect 8042 31642 8052 31698
rect 7976 31556 7988 31642
rect 8040 31556 8052 31642
rect 7976 31500 7986 31556
rect 8042 31500 8052 31556
rect 7976 31414 7988 31500
rect 8040 31414 8052 31500
rect 7976 31358 7986 31414
rect 8042 31358 8052 31414
rect 7976 31272 7988 31358
rect 8040 31272 8052 31358
rect 7976 31216 7986 31272
rect 8042 31216 8052 31272
rect 7976 31130 7988 31216
rect 8040 31130 8052 31216
rect 7976 31074 7986 31130
rect 8042 31074 8052 31130
rect 7976 30988 7988 31074
rect 8040 30988 8052 31074
rect 9368 32693 9444 32703
rect 9368 32637 9378 32693
rect 9434 32637 9444 32693
rect 9368 32551 9380 32637
rect 9432 32551 9444 32637
rect 9368 32495 9378 32551
rect 9434 32495 9444 32551
rect 9368 32409 9380 32495
rect 9432 32409 9444 32495
rect 9368 32353 9378 32409
rect 9434 32353 9444 32409
rect 9368 32267 9380 32353
rect 9432 32267 9444 32353
rect 9368 32211 9378 32267
rect 9434 32211 9444 32267
rect 9368 32125 9380 32211
rect 9432 32125 9444 32211
rect 9368 32069 9378 32125
rect 9434 32069 9444 32125
rect 9368 31983 9380 32069
rect 9432 31983 9444 32069
rect 9368 31927 9378 31983
rect 9434 31927 9444 31983
rect 9368 31841 9380 31927
rect 9432 31841 9444 31927
rect 9368 31785 9378 31841
rect 9434 31785 9444 31841
rect 9368 31699 9380 31785
rect 9432 31699 9444 31785
rect 9368 31643 9378 31699
rect 9434 31643 9444 31699
rect 9368 31557 9380 31643
rect 9432 31557 9444 31643
rect 9368 31501 9378 31557
rect 9434 31501 9444 31557
rect 9368 31415 9380 31501
rect 9432 31415 9444 31501
rect 9368 31359 9378 31415
rect 9434 31359 9444 31415
rect 9368 31273 9380 31359
rect 9432 31273 9444 31359
rect 9368 31217 9378 31273
rect 9434 31217 9444 31273
rect 9368 31131 9380 31217
rect 9432 31131 9444 31217
rect 9368 31075 9378 31131
rect 9434 31075 9444 31131
rect 9368 31065 9444 31075
rect 9784 32693 9860 32703
rect 9784 32637 9794 32693
rect 9850 32637 9860 32693
rect 9784 32551 9796 32637
rect 9848 32551 9860 32637
rect 9784 32495 9794 32551
rect 9850 32495 9860 32551
rect 9784 32409 9796 32495
rect 9848 32409 9860 32495
rect 9784 32353 9794 32409
rect 9850 32353 9860 32409
rect 9784 32267 9796 32353
rect 9848 32267 9860 32353
rect 9784 32211 9794 32267
rect 9850 32211 9860 32267
rect 9784 32125 9796 32211
rect 9848 32125 9860 32211
rect 9784 32069 9794 32125
rect 9850 32069 9860 32125
rect 9784 31983 9796 32069
rect 9848 31983 9860 32069
rect 9784 31927 9794 31983
rect 9850 31927 9860 31983
rect 9784 31841 9796 31927
rect 9848 31841 9860 31927
rect 9784 31785 9794 31841
rect 9850 31785 9860 31841
rect 9784 31699 9796 31785
rect 9848 31699 9860 31785
rect 9784 31643 9794 31699
rect 9850 31643 9860 31699
rect 9784 31557 9796 31643
rect 9848 31557 9860 31643
rect 9784 31501 9794 31557
rect 9850 31501 9860 31557
rect 9784 31415 9796 31501
rect 9848 31415 9860 31501
rect 9784 31359 9794 31415
rect 9850 31359 9860 31415
rect 9784 31273 9796 31359
rect 9848 31273 9860 31359
rect 9784 31217 9794 31273
rect 9850 31217 9860 31273
rect 9784 31131 9796 31217
rect 9848 31131 9860 31217
rect 9784 31075 9794 31131
rect 9850 31075 9860 31131
rect 9784 31065 9860 31075
rect 10272 32693 10348 32703
rect 10272 32637 10282 32693
rect 10338 32637 10348 32693
rect 10272 32551 10284 32637
rect 10336 32551 10348 32637
rect 10272 32495 10282 32551
rect 10338 32495 10348 32551
rect 10272 32409 10284 32495
rect 10336 32409 10348 32495
rect 10272 32353 10282 32409
rect 10338 32353 10348 32409
rect 10272 32267 10284 32353
rect 10336 32267 10348 32353
rect 10272 32211 10282 32267
rect 10338 32211 10348 32267
rect 10272 32125 10284 32211
rect 10336 32125 10348 32211
rect 10272 32069 10282 32125
rect 10338 32069 10348 32125
rect 10272 31983 10284 32069
rect 10336 31983 10348 32069
rect 10272 31927 10282 31983
rect 10338 31927 10348 31983
rect 10272 31841 10284 31927
rect 10336 31841 10348 31927
rect 10272 31785 10282 31841
rect 10338 31785 10348 31841
rect 10272 31699 10284 31785
rect 10336 31699 10348 31785
rect 10272 31643 10282 31699
rect 10338 31643 10348 31699
rect 10272 31557 10284 31643
rect 10336 31557 10348 31643
rect 10272 31501 10282 31557
rect 10338 31501 10348 31557
rect 10272 31415 10284 31501
rect 10336 31415 10348 31501
rect 10272 31359 10282 31415
rect 10338 31359 10348 31415
rect 10272 31273 10284 31359
rect 10336 31273 10348 31359
rect 10272 31217 10282 31273
rect 10338 31217 10348 31273
rect 10272 31131 10284 31217
rect 10336 31131 10348 31217
rect 10272 31075 10282 31131
rect 10338 31075 10348 31131
rect 10272 31065 10348 31075
rect 10760 32642 10836 32652
rect 10760 32586 10770 32642
rect 10826 32586 10836 32642
rect 10760 32500 10772 32586
rect 10824 32500 10836 32586
rect 10760 32444 10770 32500
rect 10826 32444 10836 32500
rect 10760 32358 10772 32444
rect 10824 32358 10836 32444
rect 10760 32302 10770 32358
rect 10826 32302 10836 32358
rect 10760 32216 10772 32302
rect 10824 32216 10836 32302
rect 10760 32160 10770 32216
rect 10826 32160 10836 32216
rect 10760 32074 10772 32160
rect 10824 32074 10836 32160
rect 10760 32018 10770 32074
rect 10826 32018 10836 32074
rect 10760 31932 10772 32018
rect 10824 31932 10836 32018
rect 10760 31876 10770 31932
rect 10826 31876 10836 31932
rect 10760 31790 10772 31876
rect 10824 31790 10836 31876
rect 10760 31734 10770 31790
rect 10826 31734 10836 31790
rect 10760 31648 10772 31734
rect 10824 31648 10836 31734
rect 10760 31592 10770 31648
rect 10826 31592 10836 31648
rect 10760 31506 10772 31592
rect 10824 31506 10836 31592
rect 10760 31450 10770 31506
rect 10826 31450 10836 31506
rect 10760 31364 10772 31450
rect 10824 31364 10836 31450
rect 10760 31308 10770 31364
rect 10826 31308 10836 31364
rect 10760 31222 10772 31308
rect 10824 31222 10836 31308
rect 10760 31166 10770 31222
rect 10826 31166 10836 31222
rect 10760 31080 10772 31166
rect 10824 31080 10836 31166
rect 10760 31024 10770 31080
rect 10826 31024 10836 31080
rect 10760 31014 10836 31024
rect 10998 32621 11010 32707
rect 11062 32621 11074 32707
rect 14380 32866 14410 32922
rect 14466 32866 14514 32922
rect 14608 32866 14694 32922
rect 14750 32866 14780 32922
rect 14380 32780 14514 32866
rect 14566 32780 14780 32866
rect 14380 32724 14410 32780
rect 14466 32724 14514 32780
rect 14608 32724 14694 32780
rect 14750 32724 14780 32780
rect 11724 32693 11800 32703
rect 10998 32565 11008 32621
rect 11064 32565 11074 32621
rect 10998 32479 11010 32565
rect 11062 32479 11074 32565
rect 10998 32423 11008 32479
rect 11064 32423 11074 32479
rect 10998 32337 11010 32423
rect 11062 32337 11074 32423
rect 10998 32281 11008 32337
rect 11064 32281 11074 32337
rect 10998 32195 11010 32281
rect 11062 32195 11074 32281
rect 10998 32139 11008 32195
rect 11064 32139 11074 32195
rect 10998 32053 11010 32139
rect 11062 32053 11074 32139
rect 10998 31997 11008 32053
rect 11064 31997 11074 32053
rect 10998 31911 11010 31997
rect 11062 31911 11074 31997
rect 10998 31855 11008 31911
rect 11064 31855 11074 31911
rect 10998 31769 11010 31855
rect 11062 31769 11074 31855
rect 10998 31713 11008 31769
rect 11064 31713 11074 31769
rect 10998 31627 11010 31713
rect 11062 31627 11074 31713
rect 10998 31571 11008 31627
rect 11064 31571 11074 31627
rect 10998 31485 11010 31571
rect 11062 31485 11074 31571
rect 10998 31429 11008 31485
rect 11064 31429 11074 31485
rect 10998 31343 11010 31429
rect 11062 31343 11074 31429
rect 10998 31287 11008 31343
rect 11064 31287 11074 31343
rect 10998 31201 11010 31287
rect 11062 31201 11074 31287
rect 10998 31145 11008 31201
rect 11064 31145 11074 31201
rect 10998 31059 11010 31145
rect 11062 31059 11074 31145
rect 10998 31003 11008 31059
rect 11064 31003 11074 31059
rect 11236 32642 11312 32652
rect 11236 32586 11246 32642
rect 11302 32586 11312 32642
rect 11236 32500 11248 32586
rect 11300 32500 11312 32586
rect 11236 32444 11246 32500
rect 11302 32444 11312 32500
rect 11236 32358 11248 32444
rect 11300 32358 11312 32444
rect 11236 32302 11246 32358
rect 11302 32302 11312 32358
rect 11236 32216 11248 32302
rect 11300 32216 11312 32302
rect 11236 32160 11246 32216
rect 11302 32160 11312 32216
rect 11236 32074 11248 32160
rect 11300 32074 11312 32160
rect 11236 32018 11246 32074
rect 11302 32018 11312 32074
rect 11236 31932 11248 32018
rect 11300 31932 11312 32018
rect 11236 31876 11246 31932
rect 11302 31876 11312 31932
rect 11236 31790 11248 31876
rect 11300 31790 11312 31876
rect 11236 31734 11246 31790
rect 11302 31734 11312 31790
rect 11236 31648 11248 31734
rect 11300 31648 11312 31734
rect 11236 31592 11246 31648
rect 11302 31592 11312 31648
rect 11236 31506 11248 31592
rect 11300 31506 11312 31592
rect 11236 31450 11246 31506
rect 11302 31450 11312 31506
rect 11236 31364 11248 31450
rect 11300 31364 11312 31450
rect 11236 31308 11246 31364
rect 11302 31308 11312 31364
rect 11236 31222 11248 31308
rect 11300 31222 11312 31308
rect 11236 31166 11246 31222
rect 11302 31166 11312 31222
rect 11236 31080 11248 31166
rect 11300 31080 11312 31166
rect 11236 31024 11246 31080
rect 11302 31024 11312 31080
rect 11724 32637 11734 32693
rect 11790 32637 11800 32693
rect 11724 32551 11736 32637
rect 11788 32551 11800 32637
rect 11724 32495 11734 32551
rect 11790 32495 11800 32551
rect 11724 32409 11736 32495
rect 11788 32409 11800 32495
rect 11724 32353 11734 32409
rect 11790 32353 11800 32409
rect 11724 32267 11736 32353
rect 11788 32267 11800 32353
rect 11724 32211 11734 32267
rect 11790 32211 11800 32267
rect 11724 32125 11736 32211
rect 11788 32125 11800 32211
rect 11724 32069 11734 32125
rect 11790 32069 11800 32125
rect 11724 31983 11736 32069
rect 11788 31983 11800 32069
rect 11724 31927 11734 31983
rect 11790 31927 11800 31983
rect 11724 31841 11736 31927
rect 11788 31841 11800 31927
rect 11724 31785 11734 31841
rect 11790 31785 11800 31841
rect 11724 31699 11736 31785
rect 11788 31699 11800 31785
rect 11724 31643 11734 31699
rect 11790 31643 11800 31699
rect 11724 31557 11736 31643
rect 11788 31557 11800 31643
rect 11724 31501 11734 31557
rect 11790 31501 11800 31557
rect 11724 31415 11736 31501
rect 11788 31415 11800 31501
rect 11724 31359 11734 31415
rect 11790 31359 11800 31415
rect 11724 31273 11736 31359
rect 11788 31273 11800 31359
rect 11724 31217 11734 31273
rect 11790 31217 11800 31273
rect 11724 31131 11736 31217
rect 11788 31131 11800 31217
rect 11724 31075 11734 31131
rect 11790 31075 11800 31131
rect 11724 31065 11800 31075
rect 12212 32692 12288 32702
rect 12212 32636 12222 32692
rect 12278 32636 12288 32692
rect 12212 32550 12224 32636
rect 12276 32550 12288 32636
rect 12212 32494 12222 32550
rect 12278 32494 12288 32550
rect 12212 32408 12224 32494
rect 12276 32408 12288 32494
rect 12212 32352 12222 32408
rect 12278 32352 12288 32408
rect 12212 32266 12224 32352
rect 12276 32266 12288 32352
rect 12212 32210 12222 32266
rect 12278 32210 12288 32266
rect 12212 32124 12224 32210
rect 12276 32124 12288 32210
rect 12212 32068 12222 32124
rect 12278 32068 12288 32124
rect 12212 31982 12224 32068
rect 12276 31982 12288 32068
rect 12212 31926 12222 31982
rect 12278 31926 12288 31982
rect 12212 31840 12224 31926
rect 12276 31840 12288 31926
rect 12212 31784 12222 31840
rect 12278 31784 12288 31840
rect 12212 31698 12224 31784
rect 12276 31698 12288 31784
rect 12212 31642 12222 31698
rect 12278 31642 12288 31698
rect 12212 31556 12224 31642
rect 12276 31556 12288 31642
rect 12212 31500 12222 31556
rect 12278 31500 12288 31556
rect 12212 31414 12224 31500
rect 12276 31414 12288 31500
rect 12212 31358 12222 31414
rect 12278 31358 12288 31414
rect 12212 31272 12224 31358
rect 12276 31272 12288 31358
rect 12212 31216 12222 31272
rect 12278 31216 12288 31272
rect 12212 31130 12224 31216
rect 12276 31130 12288 31216
rect 12212 31074 12222 31130
rect 12278 31074 12288 31130
rect 11236 31014 11312 31024
rect 10998 30993 11074 31003
rect 7976 30932 7986 30988
rect 8042 30932 8052 30988
rect 7976 30846 7988 30932
rect 8040 30846 8052 30932
rect 12212 30988 12224 31074
rect 12276 30988 12288 31074
rect 12212 30932 12222 30988
rect 12278 30932 12288 30988
rect 7976 30790 7986 30846
rect 8042 30790 8052 30846
rect 7976 30704 7988 30790
rect 8040 30704 8052 30790
rect 7976 30648 7986 30704
rect 8042 30648 8052 30704
rect 9062 30858 10592 30870
rect 9062 30770 10528 30858
rect 7976 30562 7988 30648
rect 8040 30562 8052 30648
rect 7976 30506 7986 30562
rect 8042 30506 8052 30562
rect 7976 30454 7988 30506
rect 8040 30454 8052 30506
rect 7976 30442 8052 30454
rect 8452 30678 8552 30690
rect 8452 30314 8476 30678
rect 8528 30314 8552 30678
rect 8452 29649 8552 30314
rect 8696 30678 8796 30690
rect 8696 30314 8720 30678
rect 8772 30314 8796 30678
rect 8696 29829 8796 30314
rect 8696 29817 8876 29829
rect 8696 29765 8708 29817
rect 8864 29765 8876 29817
rect 8696 29753 8876 29765
rect 8452 29637 8632 29649
rect 8452 29585 8464 29637
rect 8620 29585 8632 29637
rect 8452 29573 8632 29585
rect 9062 29469 9162 30770
rect 9062 29313 9088 29469
rect 9140 29313 9162 29469
rect 9062 29301 9162 29313
rect 10016 30678 10116 30690
rect 10016 30314 10040 30678
rect 10092 30314 10116 30678
rect 10516 30494 10528 30770
rect 10580 30494 10592 30858
rect 10516 30482 10592 30494
rect 10821 30858 12044 30870
rect 10821 30770 11980 30858
rect 10016 29469 10116 30314
rect 10016 29313 10042 29469
rect 10094 29313 10116 29469
rect 10016 29301 10116 29313
rect 10821 29469 10921 30770
rect 10821 29313 10847 29469
rect 10899 29313 10921 29469
rect 11468 30678 11568 30690
rect 11468 30314 11492 30678
rect 11544 30314 11568 30678
rect 11968 30494 11980 30770
rect 12032 30494 12044 30858
rect 11968 30482 12044 30494
rect 12212 30846 12224 30932
rect 12276 30846 12288 30932
rect 12212 30790 12222 30846
rect 12278 30790 12288 30846
rect 12212 30704 12224 30790
rect 12276 30704 12288 30790
rect 12212 30648 12222 30704
rect 12278 30648 12288 30704
rect 12212 30562 12224 30648
rect 12276 30562 12288 30648
rect 12212 30506 12222 30562
rect 12278 30506 12288 30562
rect 12212 30454 12224 30506
rect 12276 30454 12288 30506
rect 12212 30442 12288 30454
rect 12628 32692 12704 32702
rect 12628 32636 12638 32692
rect 12694 32636 12704 32692
rect 12628 32550 12640 32636
rect 12692 32550 12704 32636
rect 12628 32494 12638 32550
rect 12694 32494 12704 32550
rect 12628 32408 12640 32494
rect 12692 32408 12704 32494
rect 12628 32352 12638 32408
rect 12694 32352 12704 32408
rect 12628 32266 12640 32352
rect 12692 32266 12704 32352
rect 12628 32210 12638 32266
rect 12694 32210 12704 32266
rect 12628 32124 12640 32210
rect 12692 32124 12704 32210
rect 12628 32068 12638 32124
rect 12694 32068 12704 32124
rect 12628 31982 12640 32068
rect 12692 31982 12704 32068
rect 12628 31926 12638 31982
rect 12694 31926 12704 31982
rect 12628 31840 12640 31926
rect 12692 31840 12704 31926
rect 12628 31784 12638 31840
rect 12694 31784 12704 31840
rect 12628 31698 12640 31784
rect 12692 31698 12704 31784
rect 12628 31642 12638 31698
rect 12694 31642 12704 31698
rect 12628 31556 12640 31642
rect 12692 31556 12704 31642
rect 12628 31500 12638 31556
rect 12694 31500 12704 31556
rect 12628 31414 12640 31500
rect 12692 31414 12704 31500
rect 12628 31358 12638 31414
rect 12694 31358 12704 31414
rect 12628 31272 12640 31358
rect 12692 31272 12704 31358
rect 12628 31216 12638 31272
rect 12694 31216 12704 31272
rect 12628 31130 12640 31216
rect 12692 31130 12704 31216
rect 12628 31074 12638 31130
rect 12694 31074 12704 31130
rect 12628 30988 12640 31074
rect 12692 30988 12704 31074
rect 12628 30932 12638 30988
rect 12694 30932 12704 30988
rect 12628 30846 12640 30932
rect 12692 30846 12704 30932
rect 12628 30790 12638 30846
rect 12694 30790 12704 30846
rect 12628 30704 12640 30790
rect 12692 30704 12704 30790
rect 12628 30648 12638 30704
rect 12694 30648 12704 30704
rect 14020 32692 14096 32702
rect 14020 32636 14030 32692
rect 14086 32636 14096 32692
rect 14020 32550 14032 32636
rect 14084 32550 14096 32636
rect 14020 32494 14030 32550
rect 14086 32494 14096 32550
rect 14020 32408 14032 32494
rect 14084 32408 14096 32494
rect 14020 32352 14030 32408
rect 14086 32352 14096 32408
rect 14020 32266 14032 32352
rect 14084 32266 14096 32352
rect 14020 32210 14030 32266
rect 14086 32210 14096 32266
rect 14020 32124 14032 32210
rect 14084 32124 14096 32210
rect 14020 32068 14030 32124
rect 14086 32068 14096 32124
rect 14020 31982 14032 32068
rect 14084 31982 14096 32068
rect 14020 31926 14030 31982
rect 14086 31926 14096 31982
rect 14020 31840 14032 31926
rect 14084 31840 14096 31926
rect 14020 31784 14030 31840
rect 14086 31784 14096 31840
rect 14020 31698 14032 31784
rect 14084 31698 14096 31784
rect 14020 31642 14030 31698
rect 14086 31642 14096 31698
rect 14020 31556 14032 31642
rect 14084 31556 14096 31642
rect 14020 31500 14030 31556
rect 14086 31500 14096 31556
rect 14020 31414 14032 31500
rect 14084 31414 14096 31500
rect 14020 31358 14030 31414
rect 14086 31358 14096 31414
rect 14020 31272 14032 31358
rect 14084 31272 14096 31358
rect 14020 31216 14030 31272
rect 14086 31216 14096 31272
rect 14020 31130 14032 31216
rect 14084 31130 14096 31216
rect 14020 31074 14030 31130
rect 14086 31074 14096 31130
rect 14020 30988 14032 31074
rect 14084 30988 14096 31074
rect 14020 30932 14030 30988
rect 14086 30932 14096 30988
rect 14020 30846 14032 30932
rect 14084 30846 14096 30932
rect 14020 30790 14030 30846
rect 14086 30790 14096 30846
rect 14020 30704 14032 30790
rect 14084 30704 14096 30790
rect 12628 30562 12640 30648
rect 12692 30562 12704 30648
rect 12628 30506 12638 30562
rect 12694 30506 12704 30562
rect 12628 30454 12640 30506
rect 12692 30454 12704 30506
rect 12628 30442 12704 30454
rect 13520 30678 13620 30690
rect 11468 29442 11568 30314
rect 13520 30314 13544 30678
rect 13596 30314 13620 30678
rect 11922 30109 13276 30119
rect 11922 30053 11932 30109
rect 11988 30107 12074 30109
rect 12130 30107 12216 30109
rect 12272 30107 12358 30109
rect 12414 30107 12500 30109
rect 12556 30107 12642 30109
rect 12698 30107 12784 30109
rect 12840 30107 12926 30109
rect 12982 30107 13068 30109
rect 13124 30107 13210 30109
rect 11988 30053 12074 30055
rect 12130 30053 12216 30055
rect 12272 30053 12358 30055
rect 12414 30053 12500 30055
rect 12556 30053 12642 30055
rect 12698 30053 12784 30055
rect 12840 30053 12926 30055
rect 12982 30053 13068 30055
rect 13124 30053 13210 30055
rect 13266 30053 13276 30109
rect 11922 30043 13276 30053
rect 13520 30021 13620 30314
rect 13764 30678 13864 30690
rect 13764 30314 13788 30678
rect 13840 30314 13864 30678
rect 14020 30648 14030 30704
rect 14086 30648 14096 30704
rect 14020 30562 14032 30648
rect 14084 30562 14096 30648
rect 14020 30506 14030 30562
rect 14086 30506 14096 30562
rect 14020 30454 14032 30506
rect 14084 30454 14096 30506
rect 14020 30442 14096 30454
rect 14380 32638 14514 32724
rect 14566 32638 14780 32724
rect 14380 32582 14410 32638
rect 14466 32582 14514 32638
rect 14608 32582 14694 32638
rect 14750 32582 14780 32638
rect 14380 32496 14514 32582
rect 14566 32496 14780 32582
rect 14380 32440 14410 32496
rect 14466 32440 14514 32496
rect 14608 32440 14694 32496
rect 14750 32440 14780 32496
rect 14380 32354 14514 32440
rect 14566 32354 14780 32440
rect 14380 32298 14410 32354
rect 14466 32298 14514 32354
rect 14608 32298 14694 32354
rect 14750 32298 14780 32354
rect 14380 32212 14514 32298
rect 14566 32212 14780 32298
rect 14380 32156 14410 32212
rect 14466 32156 14514 32212
rect 14608 32156 14694 32212
rect 14750 32156 14780 32212
rect 14380 32070 14514 32156
rect 14566 32070 14780 32156
rect 14380 32014 14410 32070
rect 14466 32014 14514 32070
rect 14608 32014 14694 32070
rect 14750 32014 14780 32070
rect 14380 31928 14514 32014
rect 14566 31928 14780 32014
rect 14380 31872 14410 31928
rect 14466 31872 14514 31928
rect 14608 31872 14694 31928
rect 14750 31872 14780 31928
rect 14380 31786 14514 31872
rect 14566 31786 14780 31872
rect 14380 31730 14410 31786
rect 14466 31730 14514 31786
rect 14608 31730 14694 31786
rect 14750 31730 14780 31786
rect 14380 31644 14514 31730
rect 14566 31644 14780 31730
rect 14380 31588 14410 31644
rect 14466 31588 14514 31644
rect 14608 31588 14694 31644
rect 14750 31588 14780 31644
rect 14380 31502 14514 31588
rect 14566 31502 14780 31588
rect 14380 31446 14410 31502
rect 14466 31446 14514 31502
rect 14608 31446 14694 31502
rect 14750 31446 14780 31502
rect 14380 31360 14514 31446
rect 14566 31360 14780 31446
rect 14380 31304 14410 31360
rect 14466 31304 14514 31360
rect 14608 31304 14694 31360
rect 14750 31304 14780 31360
rect 14380 31218 14514 31304
rect 14566 31218 14780 31304
rect 14380 31162 14410 31218
rect 14466 31162 14514 31218
rect 14608 31162 14694 31218
rect 14750 31162 14780 31218
rect 14380 31076 14514 31162
rect 14566 31076 14780 31162
rect 14380 31020 14410 31076
rect 14466 31020 14514 31076
rect 14608 31020 14694 31076
rect 14750 31020 14780 31076
rect 14380 30934 14514 31020
rect 14566 30934 14780 31020
rect 14380 30878 14410 30934
rect 14466 30878 14514 30934
rect 14608 30878 14694 30934
rect 14750 30878 14780 30934
rect 14380 30792 14514 30878
rect 14566 30792 14780 30878
rect 14380 30736 14410 30792
rect 14466 30736 14514 30792
rect 14608 30736 14694 30792
rect 14750 30736 14780 30792
rect 14380 30650 14514 30736
rect 14566 30650 14780 30736
rect 14380 30594 14410 30650
rect 14466 30594 14514 30650
rect 14608 30594 14694 30650
rect 14750 30594 14780 30650
rect 14380 30508 14514 30594
rect 14566 30508 14780 30594
rect 14380 30452 14410 30508
rect 14466 30452 14514 30508
rect 14608 30452 14694 30508
rect 14750 30452 14780 30508
rect 13764 30201 13864 30314
rect 13764 30101 14059 30201
rect 13520 29921 13879 30021
rect 13519 29817 13699 29829
rect 13519 29765 13531 29817
rect 13687 29765 13699 29817
rect 13519 29753 13699 29765
rect 13339 29637 13519 29649
rect 13339 29585 13351 29637
rect 13507 29585 13519 29637
rect 13339 29573 13519 29585
rect 11390 29430 11570 29442
rect 11390 29378 11402 29430
rect 11558 29378 11570 29430
rect 11390 29366 11570 29378
rect 10821 29301 10921 29313
rect 13411 28401 13519 29573
rect 13599 28401 13699 29753
rect 13779 28401 13879 29921
rect 13959 28401 14059 30101
rect 14380 30167 14514 30452
rect 14566 30167 14780 30452
rect 14380 30111 14410 30167
rect 14466 30111 14514 30167
rect 14608 30111 14694 30167
rect 14750 30111 14780 30167
rect 14380 30055 14514 30111
rect 14566 30055 14780 30111
rect 14380 30025 14780 30055
rect 14380 29969 14410 30025
rect 14466 29969 14552 30025
rect 14608 29969 14694 30025
rect 14750 29969 14780 30025
rect 14380 29883 14780 29969
rect 14380 29827 14410 29883
rect 14466 29827 14552 29883
rect 14608 29827 14694 29883
rect 14750 29827 14780 29883
rect 14380 29741 14780 29827
rect 14380 29685 14410 29741
rect 14466 29685 14552 29741
rect 14608 29685 14694 29741
rect 14750 29685 14780 29741
rect 14380 29599 14780 29685
rect 14380 29543 14410 29599
rect 14466 29543 14552 29599
rect 14608 29543 14694 29599
rect 14750 29543 14780 29599
rect 14380 29457 14780 29543
rect 14380 29401 14410 29457
rect 14466 29401 14552 29457
rect 14608 29401 14694 29457
rect 14750 29401 14780 29457
rect 14380 29315 14780 29401
rect 14380 29259 14410 29315
rect 14466 29259 14552 29315
rect 14608 29259 14694 29315
rect 14750 29259 14780 29315
rect 14380 29173 14780 29259
rect 14380 29117 14410 29173
rect 14466 29117 14552 29173
rect 14608 29117 14694 29173
rect 14750 29117 14780 29173
rect 14380 29031 14780 29117
rect 14380 28975 14410 29031
rect 14466 28975 14552 29031
rect 14608 28975 14694 29031
rect 14750 28975 14780 29031
rect 14380 28889 14780 28975
rect 14380 28833 14410 28889
rect 14466 28833 14552 28889
rect 14608 28833 14694 28889
rect 14750 28833 14780 28889
rect 165 27943 175 27999
rect 231 27943 317 27999
rect 373 27943 586 27999
rect 165 27857 586 27943
rect 165 27801 175 27857
rect 231 27801 317 27857
rect 373 27801 586 27857
rect 165 27715 586 27801
rect 165 27659 175 27715
rect 231 27659 317 27715
rect 373 27659 586 27715
rect 165 27573 586 27659
rect 165 27517 175 27573
rect 231 27517 317 27573
rect 373 27517 586 27573
rect 165 27431 586 27517
rect 165 27375 175 27431
rect 231 27375 317 27431
rect 373 27375 586 27431
rect 165 27289 586 27375
rect 165 27233 175 27289
rect 231 27233 317 27289
rect 373 27233 586 27289
rect 165 27223 586 27233
rect 165 14114 383 27223
rect 14380 26948 14780 28833
rect 14380 26892 14410 26948
rect 14466 26892 14552 26948
rect 14608 26892 14694 26948
rect 14750 26892 14780 26948
rect 14380 26806 14780 26892
rect 14380 26750 14410 26806
rect 14466 26750 14552 26806
rect 14608 26750 14694 26806
rect 14750 26750 14780 26806
rect 14380 26664 14780 26750
rect 14380 26608 14410 26664
rect 14466 26608 14552 26664
rect 14608 26608 14694 26664
rect 14750 26608 14780 26664
rect 14380 26522 14780 26608
rect 14380 26466 14410 26522
rect 14466 26466 14552 26522
rect 14608 26466 14694 26522
rect 14750 26466 14780 26522
rect 14380 26380 14780 26466
rect 14380 26324 14410 26380
rect 14466 26324 14552 26380
rect 14608 26324 14694 26380
rect 14750 26324 14780 26380
rect 14380 26238 14780 26324
rect 14380 26182 14410 26238
rect 14466 26182 14552 26238
rect 14608 26182 14694 26238
rect 14750 26182 14780 26238
rect 14380 26096 14780 26182
rect 14380 26040 14410 26096
rect 14466 26040 14552 26096
rect 14608 26040 14694 26096
rect 14750 26040 14780 26096
rect 14380 25954 14780 26040
rect 14380 25898 14410 25954
rect 14466 25898 14552 25954
rect 14608 25898 14694 25954
rect 14750 25898 14780 25954
rect 14380 25812 14780 25898
rect 14380 25756 14410 25812
rect 14466 25756 14552 25812
rect 14608 25756 14694 25812
rect 14750 25756 14780 25812
rect 14380 25670 14780 25756
rect 14380 25614 14410 25670
rect 14466 25614 14552 25670
rect 14608 25614 14694 25670
rect 14750 25614 14780 25670
rect 14380 25528 14780 25614
rect 14380 25472 14410 25528
rect 14466 25472 14552 25528
rect 14608 25472 14694 25528
rect 14750 25472 14780 25528
rect 14380 25386 14780 25472
rect 14380 25330 14410 25386
rect 14466 25330 14552 25386
rect 14608 25330 14694 25386
rect 14750 25330 14780 25386
rect 14380 25244 14780 25330
rect 14380 25188 14410 25244
rect 14466 25188 14552 25244
rect 14608 25188 14694 25244
rect 14750 25188 14780 25244
rect 14380 25102 14780 25188
rect 14380 25046 14410 25102
rect 14466 25046 14552 25102
rect 14608 25046 14694 25102
rect 14750 25046 14780 25102
rect 14380 24960 14780 25046
rect 14380 24904 14410 24960
rect 14466 24904 14552 24960
rect 14608 24904 14694 24960
rect 14750 24904 14780 24960
rect 14380 24818 14780 24904
rect 14380 24762 14410 24818
rect 14466 24762 14552 24818
rect 14608 24762 14694 24818
rect 14750 24762 14780 24818
rect 14380 24676 14780 24762
rect 14380 24620 14410 24676
rect 14466 24620 14552 24676
rect 14608 24620 14694 24676
rect 14750 24620 14780 24676
rect 14380 24534 14780 24620
rect 14380 24478 14410 24534
rect 14466 24478 14552 24534
rect 14608 24478 14694 24534
rect 14750 24478 14780 24534
rect 14380 24392 14780 24478
rect 14380 24336 14410 24392
rect 14466 24336 14552 24392
rect 14608 24336 14694 24392
rect 14750 24336 14780 24392
rect 14380 24250 14780 24336
rect 14380 24194 14410 24250
rect 14466 24194 14552 24250
rect 14608 24194 14694 24250
rect 14750 24194 14780 24250
rect 14380 24108 14780 24194
rect 14380 24052 14410 24108
rect 14466 24052 14552 24108
rect 14608 24052 14694 24108
rect 14750 24052 14780 24108
rect 14380 23748 14780 24052
rect 14380 23692 14410 23748
rect 14466 23692 14552 23748
rect 14608 23692 14694 23748
rect 14750 23692 14780 23748
rect 14380 23606 14780 23692
rect 14380 23550 14410 23606
rect 14466 23550 14552 23606
rect 14608 23550 14694 23606
rect 14750 23550 14780 23606
rect 14380 23464 14780 23550
rect 14380 23408 14410 23464
rect 14466 23408 14552 23464
rect 14608 23408 14694 23464
rect 14750 23408 14780 23464
rect 14380 23322 14780 23408
rect 14380 23266 14410 23322
rect 14466 23266 14552 23322
rect 14608 23266 14694 23322
rect 14750 23266 14780 23322
rect 14380 23180 14780 23266
rect 14380 23124 14410 23180
rect 14466 23124 14552 23180
rect 14608 23124 14694 23180
rect 14750 23124 14780 23180
rect 14380 23038 14780 23124
rect 14380 22982 14410 23038
rect 14466 22982 14552 23038
rect 14608 22982 14694 23038
rect 14750 22982 14780 23038
rect 14380 22896 14780 22982
rect 14380 22840 14410 22896
rect 14466 22840 14552 22896
rect 14608 22840 14694 22896
rect 14750 22840 14780 22896
rect 14380 22754 14780 22840
rect 14380 22698 14410 22754
rect 14466 22698 14552 22754
rect 14608 22698 14694 22754
rect 14750 22698 14780 22754
rect 14380 22612 14780 22698
rect 14380 22556 14410 22612
rect 14466 22556 14552 22612
rect 14608 22556 14694 22612
rect 14750 22556 14780 22612
rect 14380 22470 14780 22556
rect 14380 22414 14410 22470
rect 14466 22414 14552 22470
rect 14608 22414 14694 22470
rect 14750 22414 14780 22470
rect 14380 22328 14780 22414
rect 14380 22272 14410 22328
rect 14466 22272 14552 22328
rect 14608 22272 14694 22328
rect 14750 22272 14780 22328
rect 14380 22186 14780 22272
rect 14380 22130 14410 22186
rect 14466 22130 14552 22186
rect 14608 22130 14694 22186
rect 14750 22130 14780 22186
rect 14380 22044 14780 22130
rect 14380 21988 14410 22044
rect 14466 21988 14552 22044
rect 14608 21988 14694 22044
rect 14750 21988 14780 22044
rect 14380 21902 14780 21988
rect 14380 21846 14410 21902
rect 14466 21846 14552 21902
rect 14608 21846 14694 21902
rect 14750 21846 14780 21902
rect 14380 21760 14780 21846
rect 14380 21704 14410 21760
rect 14466 21704 14552 21760
rect 14608 21704 14694 21760
rect 14750 21704 14780 21760
rect 14380 21618 14780 21704
rect 14380 21562 14410 21618
rect 14466 21562 14552 21618
rect 14608 21562 14694 21618
rect 14750 21562 14780 21618
rect 14380 21476 14780 21562
rect 14380 21420 14410 21476
rect 14466 21420 14552 21476
rect 14608 21420 14694 21476
rect 14750 21420 14780 21476
rect 14380 21334 14780 21420
rect 14380 21278 14410 21334
rect 14466 21278 14552 21334
rect 14608 21278 14694 21334
rect 14750 21278 14780 21334
rect 14380 21192 14780 21278
rect 14380 21136 14410 21192
rect 14466 21136 14552 21192
rect 14608 21136 14694 21192
rect 14750 21136 14780 21192
rect 14380 21050 14780 21136
rect 14380 20994 14410 21050
rect 14466 20994 14552 21050
rect 14608 20994 14694 21050
rect 14750 20994 14780 21050
rect 14380 20908 14780 20994
rect 14380 20852 14410 20908
rect 14466 20852 14552 20908
rect 14608 20852 14694 20908
rect 14750 20852 14780 20908
rect 14380 20548 14780 20852
rect 14380 20492 14410 20548
rect 14466 20492 14552 20548
rect 14608 20492 14694 20548
rect 14750 20492 14780 20548
rect 14380 20406 14780 20492
rect 14380 20350 14410 20406
rect 14466 20350 14552 20406
rect 14608 20350 14694 20406
rect 14750 20350 14780 20406
rect 14380 20264 14780 20350
rect 14380 20208 14410 20264
rect 14466 20208 14552 20264
rect 14608 20208 14694 20264
rect 14750 20208 14780 20264
rect 14380 20122 14780 20208
rect 14380 20066 14410 20122
rect 14466 20066 14552 20122
rect 14608 20066 14694 20122
rect 14750 20066 14780 20122
rect 14380 19980 14780 20066
rect 14380 19924 14410 19980
rect 14466 19924 14552 19980
rect 14608 19924 14694 19980
rect 14750 19924 14780 19980
rect 14380 19838 14780 19924
rect 14380 19782 14410 19838
rect 14466 19782 14552 19838
rect 14608 19782 14694 19838
rect 14750 19782 14780 19838
rect 14380 19696 14780 19782
rect 14380 19640 14410 19696
rect 14466 19640 14552 19696
rect 14608 19640 14694 19696
rect 14750 19640 14780 19696
rect 14380 19554 14780 19640
rect 14380 19498 14410 19554
rect 14466 19498 14552 19554
rect 14608 19498 14694 19554
rect 14750 19498 14780 19554
rect 14380 19412 14780 19498
rect 14380 19356 14410 19412
rect 14466 19356 14552 19412
rect 14608 19356 14694 19412
rect 14750 19356 14780 19412
rect 14380 19270 14780 19356
rect 14380 19214 14410 19270
rect 14466 19214 14552 19270
rect 14608 19214 14694 19270
rect 14750 19214 14780 19270
rect 14380 19128 14780 19214
rect 14380 19072 14410 19128
rect 14466 19072 14552 19128
rect 14608 19072 14694 19128
rect 14750 19072 14780 19128
rect 14380 18986 14780 19072
rect 14380 18930 14410 18986
rect 14466 18930 14552 18986
rect 14608 18930 14694 18986
rect 14750 18930 14780 18986
rect 14380 18844 14780 18930
rect 14380 18788 14410 18844
rect 14466 18788 14552 18844
rect 14608 18788 14694 18844
rect 14750 18788 14780 18844
rect 14380 18702 14780 18788
rect 14380 18646 14410 18702
rect 14466 18646 14552 18702
rect 14608 18646 14694 18702
rect 14750 18646 14780 18702
rect 14380 18560 14780 18646
rect 14380 18504 14410 18560
rect 14466 18504 14552 18560
rect 14608 18504 14694 18560
rect 14750 18504 14780 18560
rect 14380 18418 14780 18504
rect 14380 18362 14410 18418
rect 14466 18362 14552 18418
rect 14608 18362 14694 18418
rect 14750 18362 14780 18418
rect 14380 18276 14780 18362
rect 14380 18220 14410 18276
rect 14466 18220 14552 18276
rect 14608 18220 14694 18276
rect 14750 18220 14780 18276
rect 14380 18134 14780 18220
rect 14380 18078 14410 18134
rect 14466 18078 14552 18134
rect 14608 18078 14694 18134
rect 14750 18078 14780 18134
rect 14380 17992 14780 18078
rect 14380 17936 14410 17992
rect 14466 17936 14552 17992
rect 14608 17936 14694 17992
rect 14750 17936 14780 17992
rect 14380 17850 14780 17936
rect 14380 17794 14410 17850
rect 14466 17794 14552 17850
rect 14608 17794 14694 17850
rect 14750 17794 14780 17850
rect 14380 17708 14780 17794
rect 14380 17652 14410 17708
rect 14466 17652 14552 17708
rect 14608 17652 14694 17708
rect 14750 17652 14780 17708
rect 14380 17400 14780 17652
rect 14380 17348 14834 17400
rect 14380 17292 14410 17348
rect 14466 17292 14552 17348
rect 14608 17292 14694 17348
rect 14750 17292 14834 17348
rect 14380 17206 14834 17292
rect 14380 17150 14410 17206
rect 14466 17150 14552 17206
rect 14608 17150 14694 17206
rect 14750 17150 14834 17206
rect 14380 17064 14834 17150
rect 14380 17008 14410 17064
rect 14466 17008 14552 17064
rect 14608 17008 14694 17064
rect 14750 17008 14834 17064
rect 14380 16922 14834 17008
rect 14380 16866 14410 16922
rect 14466 16866 14552 16922
rect 14608 16866 14694 16922
rect 14750 16866 14834 16922
rect 14380 16780 14834 16866
rect 14380 16724 14410 16780
rect 14466 16724 14552 16780
rect 14608 16724 14694 16780
rect 14750 16724 14834 16780
rect 14380 16638 14834 16724
rect 14380 16582 14410 16638
rect 14466 16582 14552 16638
rect 14608 16582 14694 16638
rect 14750 16582 14834 16638
rect 14380 16496 14834 16582
rect 14380 16440 14410 16496
rect 14466 16440 14552 16496
rect 14608 16440 14694 16496
rect 14750 16440 14834 16496
rect 14380 16354 14834 16440
rect 14380 16298 14410 16354
rect 14466 16298 14552 16354
rect 14608 16298 14694 16354
rect 14750 16298 14834 16354
rect 14380 16212 14834 16298
rect 14380 16156 14410 16212
rect 14466 16156 14552 16212
rect 14608 16156 14694 16212
rect 14750 16156 14834 16212
rect 14380 16070 14834 16156
rect 14380 16014 14410 16070
rect 14466 16014 14552 16070
rect 14608 16014 14694 16070
rect 14750 16014 14834 16070
rect 14380 15928 14834 16014
rect 14380 15872 14410 15928
rect 14466 15872 14552 15928
rect 14608 15872 14694 15928
rect 14750 15872 14834 15928
rect 14380 15786 14834 15872
rect 14380 15730 14410 15786
rect 14466 15730 14552 15786
rect 14608 15730 14694 15786
rect 14750 15730 14834 15786
rect 14380 15644 14834 15730
rect 14380 15588 14410 15644
rect 14466 15588 14552 15644
rect 14608 15588 14694 15644
rect 14750 15588 14834 15644
rect 14380 15502 14834 15588
rect 14380 15446 14410 15502
rect 14466 15446 14552 15502
rect 14608 15446 14694 15502
rect 14750 15446 14834 15502
rect 14380 15360 14834 15446
rect 14380 15304 14410 15360
rect 14466 15304 14552 15360
rect 14608 15304 14694 15360
rect 14750 15304 14834 15360
rect 14380 15218 14834 15304
rect 14380 15162 14410 15218
rect 14466 15162 14552 15218
rect 14608 15162 14694 15218
rect 14750 15162 14834 15218
rect 14380 15076 14834 15162
rect 14380 15020 14410 15076
rect 14466 15020 14552 15076
rect 14608 15020 14694 15076
rect 14750 15020 14834 15076
rect 14380 14934 14834 15020
rect 14380 14878 14410 14934
rect 14466 14878 14552 14934
rect 14608 14878 14694 14934
rect 14750 14878 14834 14934
rect 14380 14792 14834 14878
rect 14380 14736 14410 14792
rect 14466 14736 14552 14792
rect 14608 14736 14694 14792
rect 14750 14736 14834 14792
rect 14380 14650 14834 14736
rect 14380 14594 14410 14650
rect 14466 14594 14552 14650
rect 14608 14594 14694 14650
rect 14750 14594 14834 14650
rect 14380 14508 14834 14594
rect 14380 14452 14410 14508
rect 14466 14452 14552 14508
rect 14608 14452 14694 14508
rect 14750 14452 14834 14508
rect 14380 14400 14834 14452
rect 165 12894 870 14114
rect 165 10948 383 12894
rect 14634 12293 14834 14400
rect 14169 11223 14834 12293
rect 165 10892 175 10948
rect 231 10892 317 10948
rect 373 10892 383 10948
rect 165 10806 383 10892
rect 165 10750 175 10806
rect 231 10750 317 10806
rect 373 10750 383 10806
rect 165 10664 383 10750
rect 165 10608 175 10664
rect 231 10608 317 10664
rect 373 10608 383 10664
rect 165 10522 383 10608
rect 165 10466 175 10522
rect 231 10466 317 10522
rect 373 10466 383 10522
rect 165 10380 383 10466
rect 165 10324 175 10380
rect 231 10324 317 10380
rect 373 10324 383 10380
rect 165 10238 383 10324
rect 165 10182 175 10238
rect 231 10182 317 10238
rect 373 10182 383 10238
rect 165 10096 383 10182
rect 165 10040 175 10096
rect 231 10040 317 10096
rect 373 10040 383 10096
rect 165 9954 383 10040
rect 165 9898 175 9954
rect 231 9898 317 9954
rect 373 9898 383 9954
rect 165 9812 383 9898
rect 165 9756 175 9812
rect 231 9756 317 9812
rect 373 9756 383 9812
rect 165 9670 383 9756
rect 165 9614 175 9670
rect 231 9614 317 9670
rect 373 9614 383 9670
rect 165 9528 383 9614
rect 165 9472 175 9528
rect 231 9472 317 9528
rect 373 9472 383 9528
rect 165 9386 383 9472
rect 165 9330 175 9386
rect 231 9330 317 9386
rect 373 9330 383 9386
rect 165 9244 383 9330
rect 165 9188 175 9244
rect 231 9188 317 9244
rect 373 9188 383 9244
rect 165 9102 383 9188
rect 165 9046 175 9102
rect 231 9046 317 9102
rect 373 9046 383 9102
rect 165 8960 383 9046
rect 165 8904 175 8960
rect 231 8904 317 8960
rect 373 8904 383 8960
rect 165 8818 383 8904
rect 165 8762 175 8818
rect 231 8762 317 8818
rect 373 8762 383 8818
rect 165 8676 383 8762
rect 165 8620 175 8676
rect 231 8620 317 8676
rect 373 8620 383 8676
rect 165 8534 383 8620
rect 165 8478 175 8534
rect 231 8478 317 8534
rect 373 8478 383 8534
rect 165 8392 383 8478
rect 165 8336 175 8392
rect 231 8336 317 8392
rect 373 8336 383 8392
rect 165 8250 383 8336
rect 165 8194 175 8250
rect 231 8194 317 8250
rect 373 8194 383 8250
rect 165 8108 383 8194
rect 165 8052 175 8108
rect 231 8052 317 8108
rect 373 8052 383 8108
rect 165 7748 383 8052
rect 165 7692 175 7748
rect 231 7692 317 7748
rect 373 7692 383 7748
rect 165 7606 383 7692
rect 165 7550 175 7606
rect 231 7550 317 7606
rect 373 7550 383 7606
rect 165 7464 383 7550
rect 165 7408 175 7464
rect 231 7408 317 7464
rect 373 7408 383 7464
rect 165 7322 383 7408
rect 165 7266 175 7322
rect 231 7266 317 7322
rect 373 7266 383 7322
rect 165 7180 383 7266
rect 165 7124 175 7180
rect 231 7124 317 7180
rect 373 7124 383 7180
rect 165 7038 383 7124
rect 165 6982 175 7038
rect 231 6982 317 7038
rect 373 6982 383 7038
rect 165 6896 383 6982
rect 165 6840 175 6896
rect 231 6840 317 6896
rect 373 6840 383 6896
rect 165 6754 383 6840
rect 165 6698 175 6754
rect 231 6698 317 6754
rect 373 6698 383 6754
rect 165 6612 383 6698
rect 165 6556 175 6612
rect 231 6556 317 6612
rect 373 6556 383 6612
rect 165 6470 383 6556
rect 165 6414 175 6470
rect 231 6414 317 6470
rect 373 6414 383 6470
rect 165 6328 383 6414
rect 165 6272 175 6328
rect 231 6272 317 6328
rect 373 6272 383 6328
rect 165 6186 383 6272
rect 165 6130 175 6186
rect 231 6130 317 6186
rect 373 6130 383 6186
rect 165 6044 383 6130
rect 165 5988 175 6044
rect 231 5988 317 6044
rect 373 5988 383 6044
rect 165 5902 383 5988
rect 165 5846 175 5902
rect 231 5846 317 5902
rect 373 5846 383 5902
rect 165 5760 383 5846
rect 165 5704 175 5760
rect 231 5704 317 5760
rect 373 5704 383 5760
rect 165 5618 383 5704
rect 165 5562 175 5618
rect 231 5562 317 5618
rect 373 5562 383 5618
rect 165 5476 383 5562
rect 165 5420 175 5476
rect 231 5420 317 5476
rect 373 5420 383 5476
rect 165 5334 383 5420
rect 165 5278 175 5334
rect 231 5278 317 5334
rect 373 5278 383 5334
rect 165 5192 383 5278
rect 165 5136 175 5192
rect 231 5136 317 5192
rect 373 5136 383 5192
rect 165 5050 383 5136
rect 165 4994 175 5050
rect 231 4994 317 5050
rect 373 4994 383 5050
rect 165 4908 383 4994
rect 165 4852 175 4908
rect 231 4852 317 4908
rect 373 4852 383 4908
rect 165 4548 383 4852
rect 165 4492 175 4548
rect 231 4492 317 4548
rect 373 4492 383 4548
rect 165 4406 383 4492
rect 165 4350 175 4406
rect 231 4350 317 4406
rect 373 4350 383 4406
rect 165 4264 383 4350
rect 165 4208 175 4264
rect 231 4208 317 4264
rect 373 4208 383 4264
rect 165 4122 383 4208
rect 165 4066 175 4122
rect 231 4066 317 4122
rect 373 4066 383 4122
rect 165 3980 383 4066
rect 165 3924 175 3980
rect 231 3924 317 3980
rect 373 3924 383 3980
rect 165 3838 383 3924
rect 165 3782 175 3838
rect 231 3782 317 3838
rect 373 3782 383 3838
rect 165 3696 383 3782
rect 165 3640 175 3696
rect 231 3640 317 3696
rect 373 3640 383 3696
rect 165 3554 383 3640
rect 165 3498 175 3554
rect 231 3498 317 3554
rect 373 3498 383 3554
rect 165 3412 383 3498
rect 165 3356 175 3412
rect 231 3356 317 3412
rect 373 3356 383 3412
rect 165 3270 383 3356
rect 165 3214 175 3270
rect 231 3214 317 3270
rect 373 3214 383 3270
rect 165 3128 383 3214
rect 165 3072 175 3128
rect 231 3072 317 3128
rect 373 3072 383 3128
rect 165 2986 383 3072
rect 165 2930 175 2986
rect 231 2930 317 2986
rect 373 2930 383 2986
rect 165 2844 383 2930
rect 165 2788 175 2844
rect 231 2788 317 2844
rect 373 2788 383 2844
rect 165 2702 383 2788
rect 165 2646 175 2702
rect 231 2646 317 2702
rect 373 2646 383 2702
rect 165 2560 383 2646
rect 165 2504 175 2560
rect 231 2504 317 2560
rect 373 2504 383 2560
rect 165 2418 383 2504
rect 165 2362 175 2418
rect 231 2362 317 2418
rect 373 2362 383 2418
rect 165 2276 383 2362
rect 165 2220 175 2276
rect 231 2220 317 2276
rect 373 2220 383 2276
rect 165 2134 383 2220
rect 165 2078 175 2134
rect 231 2078 317 2134
rect 373 2078 383 2134
rect 165 1992 383 2078
rect 165 1936 175 1992
rect 231 1936 317 1992
rect 373 1936 383 1992
rect 165 1850 383 1936
rect 165 1794 175 1850
rect 231 1794 317 1850
rect 373 1794 383 1850
rect 165 1708 383 1794
rect 165 1652 175 1708
rect 231 1652 317 1708
rect 373 1652 383 1708
rect 165 1600 383 1652
<< via2 >>
rect 56 52543 112 52567
rect 56 52511 58 52543
rect 58 52511 110 52543
rect 110 52511 112 52543
rect 56 52369 58 52425
rect 58 52369 110 52425
rect 110 52369 112 52425
rect 56 52227 58 52283
rect 58 52227 110 52283
rect 110 52227 112 52283
rect 56 52085 58 52141
rect 58 52085 110 52141
rect 110 52085 112 52141
rect 56 51943 58 51999
rect 58 51943 110 51999
rect 110 51943 112 51999
rect 56 51801 58 51857
rect 58 51801 110 51857
rect 110 51801 112 51857
rect 56 51659 58 51715
rect 58 51659 110 51715
rect 110 51659 112 51715
rect 56 51517 58 51573
rect 58 51517 110 51573
rect 110 51517 112 51573
rect 56 51375 58 51431
rect 58 51375 110 51431
rect 110 51375 112 51431
rect 56 51243 58 51289
rect 58 51243 110 51289
rect 110 51243 112 51289
rect 56 51233 112 51243
rect 214 50904 270 50960
rect 356 50904 412 50960
rect 498 50904 554 50960
rect 214 50762 270 50818
rect 356 50762 412 50818
rect 498 50762 554 50818
rect 214 50620 270 50676
rect 356 50620 412 50676
rect 498 50620 554 50676
rect 214 50478 270 50534
rect 356 50478 412 50534
rect 498 50478 554 50534
rect 214 50336 270 50392
rect 356 50336 412 50392
rect 498 50336 554 50392
rect 214 50194 270 50250
rect 356 50194 412 50250
rect 498 50194 554 50250
rect 214 50052 270 50108
rect 356 50052 412 50108
rect 498 50052 554 50108
rect 214 49910 270 49966
rect 356 49910 412 49966
rect 498 49910 554 49966
rect 214 49768 270 49824
rect 356 49768 412 49824
rect 498 49768 554 49824
rect 214 49626 270 49682
rect 356 49626 412 49682
rect 498 49626 554 49682
rect 214 39704 270 39760
rect 356 39704 412 39760
rect 498 39704 554 39760
rect 214 39562 270 39618
rect 356 39562 412 39618
rect 498 39562 554 39618
rect 214 39420 270 39476
rect 356 39420 412 39476
rect 498 39420 554 39476
rect 214 39278 270 39334
rect 356 39278 412 39334
rect 498 39278 554 39334
rect 214 39136 270 39192
rect 356 39136 412 39192
rect 498 39136 554 39192
rect 214 38994 270 39050
rect 356 38994 412 39050
rect 498 38994 554 39050
rect 214 38852 270 38908
rect 356 38852 412 38908
rect 498 38852 554 38908
rect 214 38710 270 38766
rect 356 38710 412 38766
rect 498 38710 554 38766
rect 214 38568 270 38624
rect 356 38568 412 38624
rect 498 38568 554 38624
rect 214 38426 270 38482
rect 356 38426 412 38482
rect 498 38426 554 38482
rect 734 52504 790 52560
rect 876 52504 932 52560
rect 1018 52504 1074 52560
rect 734 52362 790 52418
rect 876 52362 932 52418
rect 1018 52362 1074 52418
rect 734 52220 790 52276
rect 876 52220 932 52276
rect 1018 52220 1074 52276
rect 734 52078 790 52134
rect 876 52078 932 52134
rect 1018 52078 1074 52134
rect 734 51936 790 51992
rect 876 51936 932 51992
rect 1018 51936 1074 51992
rect 734 51794 790 51850
rect 876 51794 932 51850
rect 1018 51794 1074 51850
rect 734 51652 790 51708
rect 876 51652 932 51708
rect 1018 51652 1074 51708
rect 734 51510 790 51566
rect 876 51510 932 51566
rect 1018 51510 1074 51566
rect 734 51368 790 51424
rect 876 51368 932 51424
rect 1018 51368 1074 51424
rect 734 51226 790 51282
rect 876 51226 932 51282
rect 1018 51226 1074 51282
rect 1896 57179 1952 57235
rect 1896 57037 1952 57093
rect 1896 56895 1952 56951
rect 1896 56753 1952 56809
rect 1896 56611 1952 56667
rect 1896 56469 1952 56525
rect 1896 56327 1952 56383
rect 1896 56185 1952 56241
rect 1896 56043 1952 56099
rect 1896 54104 1952 54160
rect 1896 53962 1952 54018
rect 1896 53820 1952 53876
rect 1896 53678 1952 53734
rect 1896 53536 1952 53592
rect 2500 57160 2556 57180
rect 2642 57160 2698 57180
rect 2784 57160 2840 57180
rect 2926 57160 2982 57180
rect 3068 57160 3124 57180
rect 2500 57124 2522 57160
rect 2522 57124 2556 57160
rect 2642 57124 2646 57160
rect 2646 57124 2698 57160
rect 2784 57124 2822 57160
rect 2822 57124 2840 57160
rect 2926 57124 2946 57160
rect 2946 57124 2982 57160
rect 3068 57124 3070 57160
rect 3070 57124 3124 57160
rect 3210 57124 3266 57180
rect 3352 57160 3408 57180
rect 3494 57160 3550 57180
rect 3636 57160 3692 57180
rect 3778 57160 3834 57180
rect 3920 57160 3976 57180
rect 3352 57124 3390 57160
rect 3390 57124 3408 57160
rect 3494 57124 3514 57160
rect 3514 57124 3550 57160
rect 3636 57124 3638 57160
rect 3638 57124 3690 57160
rect 3690 57124 3692 57160
rect 3778 57124 3814 57160
rect 3814 57124 3834 57160
rect 3920 57124 3938 57160
rect 3938 57124 3976 57160
rect 4062 57124 4118 57180
rect 4204 57160 4260 57180
rect 4346 57160 4402 57180
rect 4488 57160 4544 57180
rect 4630 57160 4686 57180
rect 4772 57160 4828 57180
rect 4914 57160 4970 57180
rect 4204 57124 4258 57160
rect 4258 57124 4260 57160
rect 4346 57124 4382 57160
rect 4382 57124 4402 57160
rect 4488 57124 4506 57160
rect 4506 57124 4544 57160
rect 4630 57124 4682 57160
rect 4682 57124 4686 57160
rect 4772 57124 4806 57160
rect 4806 57124 4828 57160
rect 4914 57124 4930 57160
rect 4930 57124 4970 57160
rect 5056 57124 5112 57180
rect 5198 57160 5254 57180
rect 5340 57160 5396 57180
rect 5482 57160 5538 57180
rect 5624 57160 5680 57180
rect 5766 57160 5822 57180
rect 5908 57160 5964 57180
rect 5198 57124 5250 57160
rect 5250 57124 5254 57160
rect 5340 57124 5374 57160
rect 5374 57124 5396 57160
rect 5482 57124 5498 57160
rect 5498 57124 5538 57160
rect 5624 57124 5674 57160
rect 5674 57124 5680 57160
rect 5766 57124 5798 57160
rect 5798 57124 5822 57160
rect 5908 57124 5922 57160
rect 5922 57124 5964 57160
rect 6050 57124 6106 57180
rect 6192 57160 6248 57180
rect 6334 57160 6390 57180
rect 6476 57160 6532 57180
rect 6618 57160 6674 57180
rect 6760 57160 6816 57180
rect 6902 57160 6958 57180
rect 6192 57124 6242 57160
rect 6242 57124 6248 57160
rect 6334 57124 6366 57160
rect 6366 57124 6390 57160
rect 6476 57124 6490 57160
rect 6490 57124 6532 57160
rect 6618 57124 6666 57160
rect 6666 57124 6674 57160
rect 6760 57124 6790 57160
rect 6790 57124 6816 57160
rect 6902 57124 6914 57160
rect 6914 57124 6958 57160
rect 7044 57124 7100 57180
rect 7186 57160 7242 57180
rect 7328 57160 7384 57180
rect 7470 57160 7526 57180
rect 7612 57160 7668 57180
rect 7754 57160 7810 57180
rect 7896 57160 7952 57180
rect 7186 57124 7234 57160
rect 7234 57124 7242 57160
rect 7328 57124 7358 57160
rect 7358 57124 7384 57160
rect 7470 57124 7482 57160
rect 7482 57124 7526 57160
rect 7612 57124 7658 57160
rect 7658 57124 7668 57160
rect 7754 57124 7782 57160
rect 7782 57124 7810 57160
rect 7896 57124 7906 57160
rect 7906 57124 7952 57160
rect 8038 57124 8094 57180
rect 8180 57160 8236 57180
rect 8322 57160 8378 57180
rect 8464 57160 8520 57180
rect 8606 57160 8662 57180
rect 8748 57160 8804 57180
rect 8890 57160 8946 57180
rect 8180 57124 8226 57160
rect 8226 57124 8236 57160
rect 8322 57124 8350 57160
rect 8350 57124 8378 57160
rect 8464 57124 8474 57160
rect 8474 57124 8520 57160
rect 8606 57124 8650 57160
rect 8650 57124 8662 57160
rect 8748 57124 8774 57160
rect 8774 57124 8804 57160
rect 8890 57124 8898 57160
rect 8898 57124 8946 57160
rect 9032 57124 9088 57180
rect 9174 57160 9230 57180
rect 9316 57160 9372 57180
rect 9458 57160 9514 57180
rect 9600 57160 9656 57180
rect 9742 57160 9798 57180
rect 9884 57160 9940 57180
rect 9174 57124 9218 57160
rect 9218 57124 9230 57160
rect 9316 57124 9342 57160
rect 9342 57124 9372 57160
rect 9458 57124 9466 57160
rect 9466 57124 9514 57160
rect 9600 57124 9642 57160
rect 9642 57124 9656 57160
rect 9742 57124 9766 57160
rect 9766 57124 9798 57160
rect 9884 57124 9890 57160
rect 9890 57124 9940 57160
rect 10026 57124 10082 57180
rect 10168 57160 10224 57180
rect 10310 57160 10366 57180
rect 10452 57160 10508 57180
rect 10594 57160 10650 57180
rect 10736 57160 10792 57180
rect 10878 57160 10934 57180
rect 10168 57124 10210 57160
rect 10210 57124 10224 57160
rect 10310 57124 10334 57160
rect 10334 57124 10366 57160
rect 10452 57124 10458 57160
rect 10458 57124 10508 57160
rect 10594 57124 10634 57160
rect 10634 57124 10650 57160
rect 10736 57124 10758 57160
rect 10758 57124 10792 57160
rect 10878 57124 10882 57160
rect 10882 57124 10934 57160
rect 11020 57124 11076 57180
rect 11162 57160 11218 57180
rect 11304 57160 11360 57180
rect 11446 57160 11502 57180
rect 11588 57160 11644 57180
rect 11730 57160 11786 57180
rect 11872 57160 11928 57180
rect 11162 57124 11202 57160
rect 11202 57124 11218 57160
rect 11304 57124 11326 57160
rect 11326 57124 11360 57160
rect 11446 57124 11450 57160
rect 11450 57124 11502 57160
rect 11588 57124 11626 57160
rect 11626 57124 11644 57160
rect 11730 57124 11750 57160
rect 11750 57124 11786 57160
rect 11872 57124 11874 57160
rect 11874 57124 11928 57160
rect 12014 57124 12070 57180
rect 12156 57160 12212 57180
rect 12298 57160 12354 57180
rect 12440 57160 12496 57180
rect 12582 57160 12638 57180
rect 12724 57160 12780 57180
rect 12156 57124 12194 57160
rect 12194 57124 12212 57160
rect 12298 57124 12318 57160
rect 12318 57124 12354 57160
rect 12440 57124 12442 57160
rect 12442 57124 12494 57160
rect 12494 57124 12496 57160
rect 12582 57124 12618 57160
rect 12618 57124 12638 57160
rect 12724 57124 12742 57160
rect 12742 57124 12780 57160
rect 12866 57124 12922 57180
rect 13008 57160 13064 57180
rect 13150 57160 13206 57180
rect 13292 57160 13348 57180
rect 13434 57160 13490 57180
rect 13576 57160 13632 57180
rect 13008 57124 13062 57160
rect 13062 57124 13064 57160
rect 13150 57124 13186 57160
rect 13186 57124 13206 57160
rect 13292 57124 13310 57160
rect 13310 57124 13348 57160
rect 13434 57124 13486 57160
rect 13486 57124 13490 57160
rect 13576 57124 13610 57160
rect 13610 57124 13632 57160
rect 2500 57036 2556 57038
rect 2642 57036 2698 57038
rect 2784 57036 2840 57038
rect 2926 57036 2982 57038
rect 3068 57036 3124 57038
rect 2500 56984 2522 57036
rect 2522 56984 2556 57036
rect 2642 56984 2646 57036
rect 2646 56984 2698 57036
rect 2784 56984 2822 57036
rect 2822 56984 2840 57036
rect 2926 56984 2946 57036
rect 2946 56984 2982 57036
rect 3068 56984 3070 57036
rect 3070 56984 3124 57036
rect 2500 56982 2556 56984
rect 2642 56982 2698 56984
rect 2784 56982 2840 56984
rect 2926 56982 2982 56984
rect 3068 56982 3124 56984
rect 3210 56982 3266 57038
rect 3352 57036 3408 57038
rect 3494 57036 3550 57038
rect 3636 57036 3692 57038
rect 3778 57036 3834 57038
rect 3920 57036 3976 57038
rect 3352 56984 3390 57036
rect 3390 56984 3408 57036
rect 3494 56984 3514 57036
rect 3514 56984 3550 57036
rect 3636 56984 3638 57036
rect 3638 56984 3690 57036
rect 3690 56984 3692 57036
rect 3778 56984 3814 57036
rect 3814 56984 3834 57036
rect 3920 56984 3938 57036
rect 3938 56984 3976 57036
rect 3352 56982 3408 56984
rect 3494 56982 3550 56984
rect 3636 56982 3692 56984
rect 3778 56982 3834 56984
rect 3920 56982 3976 56984
rect 4062 56982 4118 57038
rect 4204 57036 4260 57038
rect 4346 57036 4402 57038
rect 4488 57036 4544 57038
rect 4630 57036 4686 57038
rect 4772 57036 4828 57038
rect 4914 57036 4970 57038
rect 4204 56984 4258 57036
rect 4258 56984 4260 57036
rect 4346 56984 4382 57036
rect 4382 56984 4402 57036
rect 4488 56984 4506 57036
rect 4506 56984 4544 57036
rect 4630 56984 4682 57036
rect 4682 56984 4686 57036
rect 4772 56984 4806 57036
rect 4806 56984 4828 57036
rect 4914 56984 4930 57036
rect 4930 56984 4970 57036
rect 4204 56982 4260 56984
rect 4346 56982 4402 56984
rect 4488 56982 4544 56984
rect 4630 56982 4686 56984
rect 4772 56982 4828 56984
rect 4914 56982 4970 56984
rect 5056 56982 5112 57038
rect 5198 57036 5254 57038
rect 5340 57036 5396 57038
rect 5482 57036 5538 57038
rect 5624 57036 5680 57038
rect 5766 57036 5822 57038
rect 5908 57036 5964 57038
rect 5198 56984 5250 57036
rect 5250 56984 5254 57036
rect 5340 56984 5374 57036
rect 5374 56984 5396 57036
rect 5482 56984 5498 57036
rect 5498 56984 5538 57036
rect 5624 56984 5674 57036
rect 5674 56984 5680 57036
rect 5766 56984 5798 57036
rect 5798 56984 5822 57036
rect 5908 56984 5922 57036
rect 5922 56984 5964 57036
rect 5198 56982 5254 56984
rect 5340 56982 5396 56984
rect 5482 56982 5538 56984
rect 5624 56982 5680 56984
rect 5766 56982 5822 56984
rect 5908 56982 5964 56984
rect 6050 56982 6106 57038
rect 6192 57036 6248 57038
rect 6334 57036 6390 57038
rect 6476 57036 6532 57038
rect 6618 57036 6674 57038
rect 6760 57036 6816 57038
rect 6902 57036 6958 57038
rect 6192 56984 6242 57036
rect 6242 56984 6248 57036
rect 6334 56984 6366 57036
rect 6366 56984 6390 57036
rect 6476 56984 6490 57036
rect 6490 56984 6532 57036
rect 6618 56984 6666 57036
rect 6666 56984 6674 57036
rect 6760 56984 6790 57036
rect 6790 56984 6816 57036
rect 6902 56984 6914 57036
rect 6914 56984 6958 57036
rect 6192 56982 6248 56984
rect 6334 56982 6390 56984
rect 6476 56982 6532 56984
rect 6618 56982 6674 56984
rect 6760 56982 6816 56984
rect 6902 56982 6958 56984
rect 7044 56982 7100 57038
rect 7186 57036 7242 57038
rect 7328 57036 7384 57038
rect 7470 57036 7526 57038
rect 7612 57036 7668 57038
rect 7754 57036 7810 57038
rect 7896 57036 7952 57038
rect 7186 56984 7234 57036
rect 7234 56984 7242 57036
rect 7328 56984 7358 57036
rect 7358 56984 7384 57036
rect 7470 56984 7482 57036
rect 7482 56984 7526 57036
rect 7612 56984 7658 57036
rect 7658 56984 7668 57036
rect 7754 56984 7782 57036
rect 7782 56984 7810 57036
rect 7896 56984 7906 57036
rect 7906 56984 7952 57036
rect 7186 56982 7242 56984
rect 7328 56982 7384 56984
rect 7470 56982 7526 56984
rect 7612 56982 7668 56984
rect 7754 56982 7810 56984
rect 7896 56982 7952 56984
rect 8038 56982 8094 57038
rect 8180 57036 8236 57038
rect 8322 57036 8378 57038
rect 8464 57036 8520 57038
rect 8606 57036 8662 57038
rect 8748 57036 8804 57038
rect 8890 57036 8946 57038
rect 8180 56984 8226 57036
rect 8226 56984 8236 57036
rect 8322 56984 8350 57036
rect 8350 56984 8378 57036
rect 8464 56984 8474 57036
rect 8474 56984 8520 57036
rect 8606 56984 8650 57036
rect 8650 56984 8662 57036
rect 8748 56984 8774 57036
rect 8774 56984 8804 57036
rect 8890 56984 8898 57036
rect 8898 56984 8946 57036
rect 8180 56982 8236 56984
rect 8322 56982 8378 56984
rect 8464 56982 8520 56984
rect 8606 56982 8662 56984
rect 8748 56982 8804 56984
rect 8890 56982 8946 56984
rect 9032 56982 9088 57038
rect 9174 57036 9230 57038
rect 9316 57036 9372 57038
rect 9458 57036 9514 57038
rect 9600 57036 9656 57038
rect 9742 57036 9798 57038
rect 9884 57036 9940 57038
rect 9174 56984 9218 57036
rect 9218 56984 9230 57036
rect 9316 56984 9342 57036
rect 9342 56984 9372 57036
rect 9458 56984 9466 57036
rect 9466 56984 9514 57036
rect 9600 56984 9642 57036
rect 9642 56984 9656 57036
rect 9742 56984 9766 57036
rect 9766 56984 9798 57036
rect 9884 56984 9890 57036
rect 9890 56984 9940 57036
rect 9174 56982 9230 56984
rect 9316 56982 9372 56984
rect 9458 56982 9514 56984
rect 9600 56982 9656 56984
rect 9742 56982 9798 56984
rect 9884 56982 9940 56984
rect 10026 56982 10082 57038
rect 10168 57036 10224 57038
rect 10310 57036 10366 57038
rect 10452 57036 10508 57038
rect 10594 57036 10650 57038
rect 10736 57036 10792 57038
rect 10878 57036 10934 57038
rect 10168 56984 10210 57036
rect 10210 56984 10224 57036
rect 10310 56984 10334 57036
rect 10334 56984 10366 57036
rect 10452 56984 10458 57036
rect 10458 56984 10508 57036
rect 10594 56984 10634 57036
rect 10634 56984 10650 57036
rect 10736 56984 10758 57036
rect 10758 56984 10792 57036
rect 10878 56984 10882 57036
rect 10882 56984 10934 57036
rect 10168 56982 10224 56984
rect 10310 56982 10366 56984
rect 10452 56982 10508 56984
rect 10594 56982 10650 56984
rect 10736 56982 10792 56984
rect 10878 56982 10934 56984
rect 11020 56982 11076 57038
rect 11162 57036 11218 57038
rect 11304 57036 11360 57038
rect 11446 57036 11502 57038
rect 11588 57036 11644 57038
rect 11730 57036 11786 57038
rect 11872 57036 11928 57038
rect 11162 56984 11202 57036
rect 11202 56984 11218 57036
rect 11304 56984 11326 57036
rect 11326 56984 11360 57036
rect 11446 56984 11450 57036
rect 11450 56984 11502 57036
rect 11588 56984 11626 57036
rect 11626 56984 11644 57036
rect 11730 56984 11750 57036
rect 11750 56984 11786 57036
rect 11872 56984 11874 57036
rect 11874 56984 11928 57036
rect 11162 56982 11218 56984
rect 11304 56982 11360 56984
rect 11446 56982 11502 56984
rect 11588 56982 11644 56984
rect 11730 56982 11786 56984
rect 11872 56982 11928 56984
rect 12014 56982 12070 57038
rect 12156 57036 12212 57038
rect 12298 57036 12354 57038
rect 12440 57036 12496 57038
rect 12582 57036 12638 57038
rect 12724 57036 12780 57038
rect 12156 56984 12194 57036
rect 12194 56984 12212 57036
rect 12298 56984 12318 57036
rect 12318 56984 12354 57036
rect 12440 56984 12442 57036
rect 12442 56984 12494 57036
rect 12494 56984 12496 57036
rect 12582 56984 12618 57036
rect 12618 56984 12638 57036
rect 12724 56984 12742 57036
rect 12742 56984 12780 57036
rect 12156 56982 12212 56984
rect 12298 56982 12354 56984
rect 12440 56982 12496 56984
rect 12582 56982 12638 56984
rect 12724 56982 12780 56984
rect 12866 56982 12922 57038
rect 13008 57036 13064 57038
rect 13150 57036 13206 57038
rect 13292 57036 13348 57038
rect 13434 57036 13490 57038
rect 13576 57036 13632 57038
rect 13008 56984 13062 57036
rect 13062 56984 13064 57036
rect 13150 56984 13186 57036
rect 13186 56984 13206 57036
rect 13292 56984 13310 57036
rect 13310 56984 13348 57036
rect 13434 56984 13486 57036
rect 13486 56984 13490 57036
rect 13576 56984 13610 57036
rect 13610 56984 13632 57036
rect 13008 56982 13064 56984
rect 13150 56982 13206 56984
rect 13292 56982 13348 56984
rect 13434 56982 13490 56984
rect 13576 56982 13632 56984
rect 2500 56860 2522 56896
rect 2522 56860 2556 56896
rect 2642 56860 2646 56896
rect 2646 56860 2698 56896
rect 2784 56860 2822 56896
rect 2822 56860 2840 56896
rect 2926 56860 2946 56896
rect 2946 56860 2982 56896
rect 3068 56860 3070 56896
rect 3070 56860 3124 56896
rect 2500 56840 2556 56860
rect 2642 56840 2698 56860
rect 2784 56840 2840 56860
rect 2926 56840 2982 56860
rect 3068 56840 3124 56860
rect 3210 56840 3266 56896
rect 3352 56860 3390 56896
rect 3390 56860 3408 56896
rect 3494 56860 3514 56896
rect 3514 56860 3550 56896
rect 3636 56860 3638 56896
rect 3638 56860 3690 56896
rect 3690 56860 3692 56896
rect 3778 56860 3814 56896
rect 3814 56860 3834 56896
rect 3920 56860 3938 56896
rect 3938 56860 3976 56896
rect 3352 56840 3408 56860
rect 3494 56840 3550 56860
rect 3636 56840 3692 56860
rect 3778 56840 3834 56860
rect 3920 56840 3976 56860
rect 4062 56840 4118 56896
rect 4204 56860 4258 56896
rect 4258 56860 4260 56896
rect 4346 56860 4382 56896
rect 4382 56860 4402 56896
rect 4488 56860 4506 56896
rect 4506 56860 4544 56896
rect 4630 56860 4682 56896
rect 4682 56860 4686 56896
rect 4772 56860 4806 56896
rect 4806 56860 4828 56896
rect 4914 56860 4930 56896
rect 4930 56860 4970 56896
rect 4204 56840 4260 56860
rect 4346 56840 4402 56860
rect 4488 56840 4544 56860
rect 4630 56840 4686 56860
rect 4772 56840 4828 56860
rect 4914 56840 4970 56860
rect 5056 56840 5112 56896
rect 5198 56860 5250 56896
rect 5250 56860 5254 56896
rect 5340 56860 5374 56896
rect 5374 56860 5396 56896
rect 5482 56860 5498 56896
rect 5498 56860 5538 56896
rect 5624 56860 5674 56896
rect 5674 56860 5680 56896
rect 5766 56860 5798 56896
rect 5798 56860 5822 56896
rect 5908 56860 5922 56896
rect 5922 56860 5964 56896
rect 5198 56840 5254 56860
rect 5340 56840 5396 56860
rect 5482 56840 5538 56860
rect 5624 56840 5680 56860
rect 5766 56840 5822 56860
rect 5908 56840 5964 56860
rect 6050 56840 6106 56896
rect 6192 56860 6242 56896
rect 6242 56860 6248 56896
rect 6334 56860 6366 56896
rect 6366 56860 6390 56896
rect 6476 56860 6490 56896
rect 6490 56860 6532 56896
rect 6618 56860 6666 56896
rect 6666 56860 6674 56896
rect 6760 56860 6790 56896
rect 6790 56860 6816 56896
rect 6902 56860 6914 56896
rect 6914 56860 6958 56896
rect 6192 56840 6248 56860
rect 6334 56840 6390 56860
rect 6476 56840 6532 56860
rect 6618 56840 6674 56860
rect 6760 56840 6816 56860
rect 6902 56840 6958 56860
rect 7044 56840 7100 56896
rect 7186 56860 7234 56896
rect 7234 56860 7242 56896
rect 7328 56860 7358 56896
rect 7358 56860 7384 56896
rect 7470 56860 7482 56896
rect 7482 56860 7526 56896
rect 7612 56860 7658 56896
rect 7658 56860 7668 56896
rect 7754 56860 7782 56896
rect 7782 56860 7810 56896
rect 7896 56860 7906 56896
rect 7906 56860 7952 56896
rect 7186 56840 7242 56860
rect 7328 56840 7384 56860
rect 7470 56840 7526 56860
rect 7612 56840 7668 56860
rect 7754 56840 7810 56860
rect 7896 56840 7952 56860
rect 8038 56840 8094 56896
rect 8180 56860 8226 56896
rect 8226 56860 8236 56896
rect 8322 56860 8350 56896
rect 8350 56860 8378 56896
rect 8464 56860 8474 56896
rect 8474 56860 8520 56896
rect 8606 56860 8650 56896
rect 8650 56860 8662 56896
rect 8748 56860 8774 56896
rect 8774 56860 8804 56896
rect 8890 56860 8898 56896
rect 8898 56860 8946 56896
rect 8180 56840 8236 56860
rect 8322 56840 8378 56860
rect 8464 56840 8520 56860
rect 8606 56840 8662 56860
rect 8748 56840 8804 56860
rect 8890 56840 8946 56860
rect 9032 56840 9088 56896
rect 9174 56860 9218 56896
rect 9218 56860 9230 56896
rect 9316 56860 9342 56896
rect 9342 56860 9372 56896
rect 9458 56860 9466 56896
rect 9466 56860 9514 56896
rect 9600 56860 9642 56896
rect 9642 56860 9656 56896
rect 9742 56860 9766 56896
rect 9766 56860 9798 56896
rect 9884 56860 9890 56896
rect 9890 56860 9940 56896
rect 9174 56840 9230 56860
rect 9316 56840 9372 56860
rect 9458 56840 9514 56860
rect 9600 56840 9656 56860
rect 9742 56840 9798 56860
rect 9884 56840 9940 56860
rect 10026 56840 10082 56896
rect 10168 56860 10210 56896
rect 10210 56860 10224 56896
rect 10310 56860 10334 56896
rect 10334 56860 10366 56896
rect 10452 56860 10458 56896
rect 10458 56860 10508 56896
rect 10594 56860 10634 56896
rect 10634 56860 10650 56896
rect 10736 56860 10758 56896
rect 10758 56860 10792 56896
rect 10878 56860 10882 56896
rect 10882 56860 10934 56896
rect 10168 56840 10224 56860
rect 10310 56840 10366 56860
rect 10452 56840 10508 56860
rect 10594 56840 10650 56860
rect 10736 56840 10792 56860
rect 10878 56840 10934 56860
rect 11020 56840 11076 56896
rect 11162 56860 11202 56896
rect 11202 56860 11218 56896
rect 11304 56860 11326 56896
rect 11326 56860 11360 56896
rect 11446 56860 11450 56896
rect 11450 56860 11502 56896
rect 11588 56860 11626 56896
rect 11626 56860 11644 56896
rect 11730 56860 11750 56896
rect 11750 56860 11786 56896
rect 11872 56860 11874 56896
rect 11874 56860 11928 56896
rect 11162 56840 11218 56860
rect 11304 56840 11360 56860
rect 11446 56840 11502 56860
rect 11588 56840 11644 56860
rect 11730 56840 11786 56860
rect 11872 56840 11928 56860
rect 12014 56840 12070 56896
rect 12156 56860 12194 56896
rect 12194 56860 12212 56896
rect 12298 56860 12318 56896
rect 12318 56860 12354 56896
rect 12440 56860 12442 56896
rect 12442 56860 12494 56896
rect 12494 56860 12496 56896
rect 12582 56860 12618 56896
rect 12618 56860 12638 56896
rect 12724 56860 12742 56896
rect 12742 56860 12780 56896
rect 12156 56840 12212 56860
rect 12298 56840 12354 56860
rect 12440 56840 12496 56860
rect 12582 56840 12638 56860
rect 12724 56840 12780 56860
rect 12866 56840 12922 56896
rect 13008 56860 13062 56896
rect 13062 56860 13064 56896
rect 13150 56860 13186 56896
rect 13186 56860 13206 56896
rect 13292 56860 13310 56896
rect 13310 56860 13348 56896
rect 13434 56860 13486 56896
rect 13486 56860 13490 56896
rect 13576 56860 13610 56896
rect 13610 56860 13632 56896
rect 13008 56840 13064 56860
rect 13150 56840 13206 56860
rect 13292 56840 13348 56860
rect 13434 56840 13490 56860
rect 13576 56840 13632 56860
rect 2500 56418 2556 56438
rect 2642 56418 2698 56438
rect 2784 56418 2840 56438
rect 2926 56418 2982 56438
rect 3068 56418 3124 56438
rect 2500 56382 2522 56418
rect 2522 56382 2556 56418
rect 2642 56382 2646 56418
rect 2646 56382 2698 56418
rect 2784 56382 2822 56418
rect 2822 56382 2840 56418
rect 2926 56382 2946 56418
rect 2946 56382 2982 56418
rect 3068 56382 3070 56418
rect 3070 56382 3124 56418
rect 3210 56382 3266 56438
rect 3352 56418 3408 56438
rect 3494 56418 3550 56438
rect 3636 56418 3692 56438
rect 3778 56418 3834 56438
rect 3920 56418 3976 56438
rect 3352 56382 3390 56418
rect 3390 56382 3408 56418
rect 3494 56382 3514 56418
rect 3514 56382 3550 56418
rect 3636 56382 3638 56418
rect 3638 56382 3690 56418
rect 3690 56382 3692 56418
rect 3778 56382 3814 56418
rect 3814 56382 3834 56418
rect 3920 56382 3938 56418
rect 3938 56382 3976 56418
rect 4062 56382 4118 56438
rect 4204 56418 4260 56438
rect 4346 56418 4402 56438
rect 4488 56418 4544 56438
rect 4630 56418 4686 56438
rect 4772 56418 4828 56438
rect 4914 56418 4970 56438
rect 4204 56382 4258 56418
rect 4258 56382 4260 56418
rect 4346 56382 4382 56418
rect 4382 56382 4402 56418
rect 4488 56382 4506 56418
rect 4506 56382 4544 56418
rect 4630 56382 4682 56418
rect 4682 56382 4686 56418
rect 4772 56382 4806 56418
rect 4806 56382 4828 56418
rect 4914 56382 4930 56418
rect 4930 56382 4970 56418
rect 5056 56382 5112 56438
rect 5198 56418 5254 56438
rect 5340 56418 5396 56438
rect 5482 56418 5538 56438
rect 5624 56418 5680 56438
rect 5766 56418 5822 56438
rect 5908 56418 5964 56438
rect 5198 56382 5250 56418
rect 5250 56382 5254 56418
rect 5340 56382 5374 56418
rect 5374 56382 5396 56418
rect 5482 56382 5498 56418
rect 5498 56382 5538 56418
rect 5624 56382 5674 56418
rect 5674 56382 5680 56418
rect 5766 56382 5798 56418
rect 5798 56382 5822 56418
rect 5908 56382 5922 56418
rect 5922 56382 5964 56418
rect 6050 56382 6106 56438
rect 6192 56418 6248 56438
rect 6334 56418 6390 56438
rect 6476 56418 6532 56438
rect 6618 56418 6674 56438
rect 6760 56418 6816 56438
rect 6902 56418 6958 56438
rect 6192 56382 6242 56418
rect 6242 56382 6248 56418
rect 6334 56382 6366 56418
rect 6366 56382 6390 56418
rect 6476 56382 6490 56418
rect 6490 56382 6532 56418
rect 6618 56382 6666 56418
rect 6666 56382 6674 56418
rect 6760 56382 6790 56418
rect 6790 56382 6816 56418
rect 6902 56382 6914 56418
rect 6914 56382 6958 56418
rect 7044 56382 7100 56438
rect 7186 56418 7242 56438
rect 7328 56418 7384 56438
rect 7470 56418 7526 56438
rect 7612 56418 7668 56438
rect 7754 56418 7810 56438
rect 7896 56418 7952 56438
rect 7186 56382 7234 56418
rect 7234 56382 7242 56418
rect 7328 56382 7358 56418
rect 7358 56382 7384 56418
rect 7470 56382 7482 56418
rect 7482 56382 7526 56418
rect 7612 56382 7658 56418
rect 7658 56382 7668 56418
rect 7754 56382 7782 56418
rect 7782 56382 7810 56418
rect 7896 56382 7906 56418
rect 7906 56382 7952 56418
rect 8038 56382 8094 56438
rect 8180 56418 8236 56438
rect 8322 56418 8378 56438
rect 8464 56418 8520 56438
rect 8606 56418 8662 56438
rect 8748 56418 8804 56438
rect 8890 56418 8946 56438
rect 8180 56382 8226 56418
rect 8226 56382 8236 56418
rect 8322 56382 8350 56418
rect 8350 56382 8378 56418
rect 8464 56382 8474 56418
rect 8474 56382 8520 56418
rect 8606 56382 8650 56418
rect 8650 56382 8662 56418
rect 8748 56382 8774 56418
rect 8774 56382 8804 56418
rect 8890 56382 8898 56418
rect 8898 56382 8946 56418
rect 9032 56382 9088 56438
rect 9174 56418 9230 56438
rect 9316 56418 9372 56438
rect 9458 56418 9514 56438
rect 9600 56418 9656 56438
rect 9742 56418 9798 56438
rect 9884 56418 9940 56438
rect 9174 56382 9218 56418
rect 9218 56382 9230 56418
rect 9316 56382 9342 56418
rect 9342 56382 9372 56418
rect 9458 56382 9466 56418
rect 9466 56382 9514 56418
rect 9600 56382 9642 56418
rect 9642 56382 9656 56418
rect 9742 56382 9766 56418
rect 9766 56382 9798 56418
rect 9884 56382 9890 56418
rect 9890 56382 9940 56418
rect 10026 56382 10082 56438
rect 10168 56418 10224 56438
rect 10310 56418 10366 56438
rect 10452 56418 10508 56438
rect 10594 56418 10650 56438
rect 10736 56418 10792 56438
rect 10878 56418 10934 56438
rect 10168 56382 10210 56418
rect 10210 56382 10224 56418
rect 10310 56382 10334 56418
rect 10334 56382 10366 56418
rect 10452 56382 10458 56418
rect 10458 56382 10508 56418
rect 10594 56382 10634 56418
rect 10634 56382 10650 56418
rect 10736 56382 10758 56418
rect 10758 56382 10792 56418
rect 10878 56382 10882 56418
rect 10882 56382 10934 56418
rect 11020 56382 11076 56438
rect 11162 56418 11218 56438
rect 11304 56418 11360 56438
rect 11446 56418 11502 56438
rect 11588 56418 11644 56438
rect 11730 56418 11786 56438
rect 11872 56418 11928 56438
rect 11162 56382 11202 56418
rect 11202 56382 11218 56418
rect 11304 56382 11326 56418
rect 11326 56382 11360 56418
rect 11446 56382 11450 56418
rect 11450 56382 11502 56418
rect 11588 56382 11626 56418
rect 11626 56382 11644 56418
rect 11730 56382 11750 56418
rect 11750 56382 11786 56418
rect 11872 56382 11874 56418
rect 11874 56382 11928 56418
rect 12014 56382 12070 56438
rect 12156 56418 12212 56438
rect 12298 56418 12354 56438
rect 12440 56418 12496 56438
rect 12582 56418 12638 56438
rect 12724 56418 12780 56438
rect 12156 56382 12194 56418
rect 12194 56382 12212 56418
rect 12298 56382 12318 56418
rect 12318 56382 12354 56418
rect 12440 56382 12442 56418
rect 12442 56382 12494 56418
rect 12494 56382 12496 56418
rect 12582 56382 12618 56418
rect 12618 56382 12638 56418
rect 12724 56382 12742 56418
rect 12742 56382 12780 56418
rect 12866 56382 12922 56438
rect 13008 56418 13064 56438
rect 13150 56418 13206 56438
rect 13292 56418 13348 56438
rect 13434 56418 13490 56438
rect 13576 56418 13632 56438
rect 13008 56382 13062 56418
rect 13062 56382 13064 56418
rect 13150 56382 13186 56418
rect 13186 56382 13206 56418
rect 13292 56382 13310 56418
rect 13310 56382 13348 56418
rect 13434 56382 13486 56418
rect 13486 56382 13490 56418
rect 13576 56382 13610 56418
rect 13610 56382 13632 56418
rect 2500 56294 2556 56296
rect 2642 56294 2698 56296
rect 2784 56294 2840 56296
rect 2926 56294 2982 56296
rect 3068 56294 3124 56296
rect 2500 56242 2522 56294
rect 2522 56242 2556 56294
rect 2642 56242 2646 56294
rect 2646 56242 2698 56294
rect 2784 56242 2822 56294
rect 2822 56242 2840 56294
rect 2926 56242 2946 56294
rect 2946 56242 2982 56294
rect 3068 56242 3070 56294
rect 3070 56242 3124 56294
rect 2500 56240 2556 56242
rect 2642 56240 2698 56242
rect 2784 56240 2840 56242
rect 2926 56240 2982 56242
rect 3068 56240 3124 56242
rect 3210 56240 3266 56296
rect 3352 56294 3408 56296
rect 3494 56294 3550 56296
rect 3636 56294 3692 56296
rect 3778 56294 3834 56296
rect 3920 56294 3976 56296
rect 3352 56242 3390 56294
rect 3390 56242 3408 56294
rect 3494 56242 3514 56294
rect 3514 56242 3550 56294
rect 3636 56242 3638 56294
rect 3638 56242 3690 56294
rect 3690 56242 3692 56294
rect 3778 56242 3814 56294
rect 3814 56242 3834 56294
rect 3920 56242 3938 56294
rect 3938 56242 3976 56294
rect 3352 56240 3408 56242
rect 3494 56240 3550 56242
rect 3636 56240 3692 56242
rect 3778 56240 3834 56242
rect 3920 56240 3976 56242
rect 4062 56240 4118 56296
rect 4204 56294 4260 56296
rect 4346 56294 4402 56296
rect 4488 56294 4544 56296
rect 4630 56294 4686 56296
rect 4772 56294 4828 56296
rect 4914 56294 4970 56296
rect 4204 56242 4258 56294
rect 4258 56242 4260 56294
rect 4346 56242 4382 56294
rect 4382 56242 4402 56294
rect 4488 56242 4506 56294
rect 4506 56242 4544 56294
rect 4630 56242 4682 56294
rect 4682 56242 4686 56294
rect 4772 56242 4806 56294
rect 4806 56242 4828 56294
rect 4914 56242 4930 56294
rect 4930 56242 4970 56294
rect 4204 56240 4260 56242
rect 4346 56240 4402 56242
rect 4488 56240 4544 56242
rect 4630 56240 4686 56242
rect 4772 56240 4828 56242
rect 4914 56240 4970 56242
rect 5056 56240 5112 56296
rect 5198 56294 5254 56296
rect 5340 56294 5396 56296
rect 5482 56294 5538 56296
rect 5624 56294 5680 56296
rect 5766 56294 5822 56296
rect 5908 56294 5964 56296
rect 5198 56242 5250 56294
rect 5250 56242 5254 56294
rect 5340 56242 5374 56294
rect 5374 56242 5396 56294
rect 5482 56242 5498 56294
rect 5498 56242 5538 56294
rect 5624 56242 5674 56294
rect 5674 56242 5680 56294
rect 5766 56242 5798 56294
rect 5798 56242 5822 56294
rect 5908 56242 5922 56294
rect 5922 56242 5964 56294
rect 5198 56240 5254 56242
rect 5340 56240 5396 56242
rect 5482 56240 5538 56242
rect 5624 56240 5680 56242
rect 5766 56240 5822 56242
rect 5908 56240 5964 56242
rect 6050 56240 6106 56296
rect 6192 56294 6248 56296
rect 6334 56294 6390 56296
rect 6476 56294 6532 56296
rect 6618 56294 6674 56296
rect 6760 56294 6816 56296
rect 6902 56294 6958 56296
rect 6192 56242 6242 56294
rect 6242 56242 6248 56294
rect 6334 56242 6366 56294
rect 6366 56242 6390 56294
rect 6476 56242 6490 56294
rect 6490 56242 6532 56294
rect 6618 56242 6666 56294
rect 6666 56242 6674 56294
rect 6760 56242 6790 56294
rect 6790 56242 6816 56294
rect 6902 56242 6914 56294
rect 6914 56242 6958 56294
rect 6192 56240 6248 56242
rect 6334 56240 6390 56242
rect 6476 56240 6532 56242
rect 6618 56240 6674 56242
rect 6760 56240 6816 56242
rect 6902 56240 6958 56242
rect 7044 56240 7100 56296
rect 7186 56294 7242 56296
rect 7328 56294 7384 56296
rect 7470 56294 7526 56296
rect 7612 56294 7668 56296
rect 7754 56294 7810 56296
rect 7896 56294 7952 56296
rect 7186 56242 7234 56294
rect 7234 56242 7242 56294
rect 7328 56242 7358 56294
rect 7358 56242 7384 56294
rect 7470 56242 7482 56294
rect 7482 56242 7526 56294
rect 7612 56242 7658 56294
rect 7658 56242 7668 56294
rect 7754 56242 7782 56294
rect 7782 56242 7810 56294
rect 7896 56242 7906 56294
rect 7906 56242 7952 56294
rect 7186 56240 7242 56242
rect 7328 56240 7384 56242
rect 7470 56240 7526 56242
rect 7612 56240 7668 56242
rect 7754 56240 7810 56242
rect 7896 56240 7952 56242
rect 8038 56240 8094 56296
rect 8180 56294 8236 56296
rect 8322 56294 8378 56296
rect 8464 56294 8520 56296
rect 8606 56294 8662 56296
rect 8748 56294 8804 56296
rect 8890 56294 8946 56296
rect 8180 56242 8226 56294
rect 8226 56242 8236 56294
rect 8322 56242 8350 56294
rect 8350 56242 8378 56294
rect 8464 56242 8474 56294
rect 8474 56242 8520 56294
rect 8606 56242 8650 56294
rect 8650 56242 8662 56294
rect 8748 56242 8774 56294
rect 8774 56242 8804 56294
rect 8890 56242 8898 56294
rect 8898 56242 8946 56294
rect 8180 56240 8236 56242
rect 8322 56240 8378 56242
rect 8464 56240 8520 56242
rect 8606 56240 8662 56242
rect 8748 56240 8804 56242
rect 8890 56240 8946 56242
rect 9032 56240 9088 56296
rect 9174 56294 9230 56296
rect 9316 56294 9372 56296
rect 9458 56294 9514 56296
rect 9600 56294 9656 56296
rect 9742 56294 9798 56296
rect 9884 56294 9940 56296
rect 9174 56242 9218 56294
rect 9218 56242 9230 56294
rect 9316 56242 9342 56294
rect 9342 56242 9372 56294
rect 9458 56242 9466 56294
rect 9466 56242 9514 56294
rect 9600 56242 9642 56294
rect 9642 56242 9656 56294
rect 9742 56242 9766 56294
rect 9766 56242 9798 56294
rect 9884 56242 9890 56294
rect 9890 56242 9940 56294
rect 9174 56240 9230 56242
rect 9316 56240 9372 56242
rect 9458 56240 9514 56242
rect 9600 56240 9656 56242
rect 9742 56240 9798 56242
rect 9884 56240 9940 56242
rect 10026 56240 10082 56296
rect 10168 56294 10224 56296
rect 10310 56294 10366 56296
rect 10452 56294 10508 56296
rect 10594 56294 10650 56296
rect 10736 56294 10792 56296
rect 10878 56294 10934 56296
rect 10168 56242 10210 56294
rect 10210 56242 10224 56294
rect 10310 56242 10334 56294
rect 10334 56242 10366 56294
rect 10452 56242 10458 56294
rect 10458 56242 10508 56294
rect 10594 56242 10634 56294
rect 10634 56242 10650 56294
rect 10736 56242 10758 56294
rect 10758 56242 10792 56294
rect 10878 56242 10882 56294
rect 10882 56242 10934 56294
rect 10168 56240 10224 56242
rect 10310 56240 10366 56242
rect 10452 56240 10508 56242
rect 10594 56240 10650 56242
rect 10736 56240 10792 56242
rect 10878 56240 10934 56242
rect 11020 56240 11076 56296
rect 11162 56294 11218 56296
rect 11304 56294 11360 56296
rect 11446 56294 11502 56296
rect 11588 56294 11644 56296
rect 11730 56294 11786 56296
rect 11872 56294 11928 56296
rect 11162 56242 11202 56294
rect 11202 56242 11218 56294
rect 11304 56242 11326 56294
rect 11326 56242 11360 56294
rect 11446 56242 11450 56294
rect 11450 56242 11502 56294
rect 11588 56242 11626 56294
rect 11626 56242 11644 56294
rect 11730 56242 11750 56294
rect 11750 56242 11786 56294
rect 11872 56242 11874 56294
rect 11874 56242 11928 56294
rect 11162 56240 11218 56242
rect 11304 56240 11360 56242
rect 11446 56240 11502 56242
rect 11588 56240 11644 56242
rect 11730 56240 11786 56242
rect 11872 56240 11928 56242
rect 12014 56240 12070 56296
rect 12156 56294 12212 56296
rect 12298 56294 12354 56296
rect 12440 56294 12496 56296
rect 12582 56294 12638 56296
rect 12724 56294 12780 56296
rect 12156 56242 12194 56294
rect 12194 56242 12212 56294
rect 12298 56242 12318 56294
rect 12318 56242 12354 56294
rect 12440 56242 12442 56294
rect 12442 56242 12494 56294
rect 12494 56242 12496 56294
rect 12582 56242 12618 56294
rect 12618 56242 12638 56294
rect 12724 56242 12742 56294
rect 12742 56242 12780 56294
rect 12156 56240 12212 56242
rect 12298 56240 12354 56242
rect 12440 56240 12496 56242
rect 12582 56240 12638 56242
rect 12724 56240 12780 56242
rect 12866 56240 12922 56296
rect 13008 56294 13064 56296
rect 13150 56294 13206 56296
rect 13292 56294 13348 56296
rect 13434 56294 13490 56296
rect 13576 56294 13632 56296
rect 13008 56242 13062 56294
rect 13062 56242 13064 56294
rect 13150 56242 13186 56294
rect 13186 56242 13206 56294
rect 13292 56242 13310 56294
rect 13310 56242 13348 56294
rect 13434 56242 13486 56294
rect 13486 56242 13490 56294
rect 13576 56242 13610 56294
rect 13610 56242 13632 56294
rect 13008 56240 13064 56242
rect 13150 56240 13206 56242
rect 13292 56240 13348 56242
rect 13434 56240 13490 56242
rect 13576 56240 13632 56242
rect 2500 56118 2522 56154
rect 2522 56118 2556 56154
rect 2642 56118 2646 56154
rect 2646 56118 2698 56154
rect 2784 56118 2822 56154
rect 2822 56118 2840 56154
rect 2926 56118 2946 56154
rect 2946 56118 2982 56154
rect 3068 56118 3070 56154
rect 3070 56118 3124 56154
rect 2500 56098 2556 56118
rect 2642 56098 2698 56118
rect 2784 56098 2840 56118
rect 2926 56098 2982 56118
rect 3068 56098 3124 56118
rect 3210 56098 3266 56154
rect 3352 56118 3390 56154
rect 3390 56118 3408 56154
rect 3494 56118 3514 56154
rect 3514 56118 3550 56154
rect 3636 56118 3638 56154
rect 3638 56118 3690 56154
rect 3690 56118 3692 56154
rect 3778 56118 3814 56154
rect 3814 56118 3834 56154
rect 3920 56118 3938 56154
rect 3938 56118 3976 56154
rect 3352 56098 3408 56118
rect 3494 56098 3550 56118
rect 3636 56098 3692 56118
rect 3778 56098 3834 56118
rect 3920 56098 3976 56118
rect 4062 56098 4118 56154
rect 4204 56118 4258 56154
rect 4258 56118 4260 56154
rect 4346 56118 4382 56154
rect 4382 56118 4402 56154
rect 4488 56118 4506 56154
rect 4506 56118 4544 56154
rect 4630 56118 4682 56154
rect 4682 56118 4686 56154
rect 4772 56118 4806 56154
rect 4806 56118 4828 56154
rect 4914 56118 4930 56154
rect 4930 56118 4970 56154
rect 4204 56098 4260 56118
rect 4346 56098 4402 56118
rect 4488 56098 4544 56118
rect 4630 56098 4686 56118
rect 4772 56098 4828 56118
rect 4914 56098 4970 56118
rect 5056 56098 5112 56154
rect 5198 56118 5250 56154
rect 5250 56118 5254 56154
rect 5340 56118 5374 56154
rect 5374 56118 5396 56154
rect 5482 56118 5498 56154
rect 5498 56118 5538 56154
rect 5624 56118 5674 56154
rect 5674 56118 5680 56154
rect 5766 56118 5798 56154
rect 5798 56118 5822 56154
rect 5908 56118 5922 56154
rect 5922 56118 5964 56154
rect 5198 56098 5254 56118
rect 5340 56098 5396 56118
rect 5482 56098 5538 56118
rect 5624 56098 5680 56118
rect 5766 56098 5822 56118
rect 5908 56098 5964 56118
rect 6050 56098 6106 56154
rect 6192 56118 6242 56154
rect 6242 56118 6248 56154
rect 6334 56118 6366 56154
rect 6366 56118 6390 56154
rect 6476 56118 6490 56154
rect 6490 56118 6532 56154
rect 6618 56118 6666 56154
rect 6666 56118 6674 56154
rect 6760 56118 6790 56154
rect 6790 56118 6816 56154
rect 6902 56118 6914 56154
rect 6914 56118 6958 56154
rect 6192 56098 6248 56118
rect 6334 56098 6390 56118
rect 6476 56098 6532 56118
rect 6618 56098 6674 56118
rect 6760 56098 6816 56118
rect 6902 56098 6958 56118
rect 7044 56098 7100 56154
rect 7186 56118 7234 56154
rect 7234 56118 7242 56154
rect 7328 56118 7358 56154
rect 7358 56118 7384 56154
rect 7470 56118 7482 56154
rect 7482 56118 7526 56154
rect 7612 56118 7658 56154
rect 7658 56118 7668 56154
rect 7754 56118 7782 56154
rect 7782 56118 7810 56154
rect 7896 56118 7906 56154
rect 7906 56118 7952 56154
rect 7186 56098 7242 56118
rect 7328 56098 7384 56118
rect 7470 56098 7526 56118
rect 7612 56098 7668 56118
rect 7754 56098 7810 56118
rect 7896 56098 7952 56118
rect 8038 56098 8094 56154
rect 8180 56118 8226 56154
rect 8226 56118 8236 56154
rect 8322 56118 8350 56154
rect 8350 56118 8378 56154
rect 8464 56118 8474 56154
rect 8474 56118 8520 56154
rect 8606 56118 8650 56154
rect 8650 56118 8662 56154
rect 8748 56118 8774 56154
rect 8774 56118 8804 56154
rect 8890 56118 8898 56154
rect 8898 56118 8946 56154
rect 8180 56098 8236 56118
rect 8322 56098 8378 56118
rect 8464 56098 8520 56118
rect 8606 56098 8662 56118
rect 8748 56098 8804 56118
rect 8890 56098 8946 56118
rect 9032 56098 9088 56154
rect 9174 56118 9218 56154
rect 9218 56118 9230 56154
rect 9316 56118 9342 56154
rect 9342 56118 9372 56154
rect 9458 56118 9466 56154
rect 9466 56118 9514 56154
rect 9600 56118 9642 56154
rect 9642 56118 9656 56154
rect 9742 56118 9766 56154
rect 9766 56118 9798 56154
rect 9884 56118 9890 56154
rect 9890 56118 9940 56154
rect 9174 56098 9230 56118
rect 9316 56098 9372 56118
rect 9458 56098 9514 56118
rect 9600 56098 9656 56118
rect 9742 56098 9798 56118
rect 9884 56098 9940 56118
rect 10026 56098 10082 56154
rect 10168 56118 10210 56154
rect 10210 56118 10224 56154
rect 10310 56118 10334 56154
rect 10334 56118 10366 56154
rect 10452 56118 10458 56154
rect 10458 56118 10508 56154
rect 10594 56118 10634 56154
rect 10634 56118 10650 56154
rect 10736 56118 10758 56154
rect 10758 56118 10792 56154
rect 10878 56118 10882 56154
rect 10882 56118 10934 56154
rect 10168 56098 10224 56118
rect 10310 56098 10366 56118
rect 10452 56098 10508 56118
rect 10594 56098 10650 56118
rect 10736 56098 10792 56118
rect 10878 56098 10934 56118
rect 11020 56098 11076 56154
rect 11162 56118 11202 56154
rect 11202 56118 11218 56154
rect 11304 56118 11326 56154
rect 11326 56118 11360 56154
rect 11446 56118 11450 56154
rect 11450 56118 11502 56154
rect 11588 56118 11626 56154
rect 11626 56118 11644 56154
rect 11730 56118 11750 56154
rect 11750 56118 11786 56154
rect 11872 56118 11874 56154
rect 11874 56118 11928 56154
rect 11162 56098 11218 56118
rect 11304 56098 11360 56118
rect 11446 56098 11502 56118
rect 11588 56098 11644 56118
rect 11730 56098 11786 56118
rect 11872 56098 11928 56118
rect 12014 56098 12070 56154
rect 12156 56118 12194 56154
rect 12194 56118 12212 56154
rect 12298 56118 12318 56154
rect 12318 56118 12354 56154
rect 12440 56118 12442 56154
rect 12442 56118 12494 56154
rect 12494 56118 12496 56154
rect 12582 56118 12618 56154
rect 12618 56118 12638 56154
rect 12724 56118 12742 56154
rect 12742 56118 12780 56154
rect 12156 56098 12212 56118
rect 12298 56098 12354 56118
rect 12440 56098 12496 56118
rect 12582 56098 12638 56118
rect 12724 56098 12780 56118
rect 12866 56098 12922 56154
rect 13008 56118 13062 56154
rect 13062 56118 13064 56154
rect 13150 56118 13186 56154
rect 13186 56118 13206 56154
rect 13292 56118 13310 56154
rect 13310 56118 13348 56154
rect 13434 56118 13486 56154
rect 13486 56118 13490 56154
rect 13576 56118 13610 56154
rect 13610 56118 13632 56154
rect 13008 56098 13064 56118
rect 13150 56098 13206 56118
rect 13292 56098 13348 56118
rect 13434 56098 13490 56118
rect 13576 56098 13632 56118
rect 4760 55729 4816 55741
rect 4760 55685 4762 55729
rect 4762 55685 4814 55729
rect 4814 55685 4816 55729
rect 4760 55543 4762 55599
rect 4762 55543 4814 55599
rect 4814 55543 4816 55599
rect 4760 55401 4762 55457
rect 4762 55401 4814 55457
rect 4814 55401 4816 55457
rect 4760 55259 4762 55315
rect 4762 55259 4814 55315
rect 4814 55259 4816 55315
rect 4760 55117 4762 55173
rect 4762 55117 4814 55173
rect 4814 55117 4816 55173
rect 4760 54975 4762 55031
rect 4762 54975 4814 55031
rect 4814 54975 4816 55031
rect 4948 55695 4950 55751
rect 4950 55695 5002 55751
rect 5002 55695 5004 55751
rect 4948 55553 4950 55609
rect 4950 55553 5002 55609
rect 5002 55553 5004 55609
rect 4948 55411 4950 55467
rect 4950 55411 5002 55467
rect 5002 55411 5004 55467
rect 4948 55269 4950 55325
rect 4950 55269 5002 55325
rect 5002 55269 5004 55325
rect 4948 55127 4950 55183
rect 4950 55127 5002 55183
rect 5002 55127 5004 55183
rect 4948 54985 4950 55041
rect 4950 54985 5002 55041
rect 5002 54985 5004 55041
rect 5436 55704 5438 55760
rect 5438 55704 5490 55760
rect 5490 55704 5492 55760
rect 5436 55562 5438 55618
rect 5438 55562 5490 55618
rect 5490 55562 5492 55618
rect 5436 55420 5438 55476
rect 5438 55420 5490 55476
rect 5490 55420 5492 55476
rect 5436 55278 5438 55334
rect 5438 55278 5490 55334
rect 5490 55278 5492 55334
rect 5436 55136 5438 55192
rect 5438 55136 5490 55192
rect 5490 55136 5492 55192
rect 5436 54994 5438 55050
rect 5438 54994 5490 55050
rect 5490 54994 5492 55050
rect 5924 55704 5926 55760
rect 5926 55704 5978 55760
rect 5978 55704 5980 55760
rect 5924 55562 5926 55618
rect 5926 55562 5978 55618
rect 5978 55562 5980 55618
rect 5924 55420 5926 55476
rect 5926 55420 5978 55476
rect 5978 55420 5980 55476
rect 5924 55278 5926 55334
rect 5926 55278 5978 55334
rect 5978 55278 5980 55334
rect 5924 55136 5926 55192
rect 5926 55136 5978 55192
rect 5978 55136 5980 55192
rect 5924 54994 5926 55050
rect 5926 54994 5978 55050
rect 5978 54994 5980 55050
rect 6106 55729 6162 55741
rect 6106 55685 6108 55729
rect 6108 55685 6160 55729
rect 6160 55685 6162 55729
rect 6106 55543 6108 55599
rect 6108 55543 6160 55599
rect 6160 55543 6162 55599
rect 6106 55401 6108 55457
rect 6108 55401 6160 55457
rect 6160 55401 6162 55457
rect 6106 55259 6108 55315
rect 6108 55259 6160 55315
rect 6160 55259 6162 55315
rect 6106 55117 6108 55173
rect 6108 55117 6160 55173
rect 6160 55117 6162 55173
rect 6106 54975 6108 55031
rect 6108 54975 6160 55031
rect 6160 54975 6162 55031
rect 6288 55704 6290 55760
rect 6290 55704 6342 55760
rect 6342 55704 6344 55760
rect 6288 55562 6290 55618
rect 6290 55562 6342 55618
rect 6342 55562 6344 55618
rect 6288 55420 6290 55476
rect 6290 55420 6342 55476
rect 6342 55420 6344 55476
rect 6288 55278 6290 55334
rect 6290 55278 6342 55334
rect 6342 55278 6344 55334
rect 6288 55136 6290 55192
rect 6290 55136 6342 55192
rect 6342 55136 6344 55192
rect 6288 54994 6290 55050
rect 6290 54994 6342 55050
rect 6342 54994 6344 55050
rect 6776 55704 6778 55760
rect 6778 55704 6830 55760
rect 6830 55704 6832 55760
rect 6776 55562 6778 55618
rect 6778 55562 6830 55618
rect 6830 55562 6832 55618
rect 6776 55420 6778 55476
rect 6778 55420 6830 55476
rect 6830 55420 6832 55476
rect 6776 55278 6778 55334
rect 6778 55278 6830 55334
rect 6830 55278 6832 55334
rect 6776 55136 6778 55192
rect 6778 55136 6830 55192
rect 6830 55136 6832 55192
rect 6776 54994 6778 55050
rect 6778 54994 6830 55050
rect 6830 54994 6832 55050
rect 7264 55704 7266 55760
rect 7266 55704 7318 55760
rect 7318 55704 7320 55760
rect 7264 55562 7266 55618
rect 7266 55562 7318 55618
rect 7318 55562 7320 55618
rect 7264 55420 7266 55476
rect 7266 55420 7318 55476
rect 7318 55420 7320 55476
rect 7264 55278 7266 55334
rect 7266 55278 7318 55334
rect 7318 55278 7320 55334
rect 7264 55136 7266 55192
rect 7266 55136 7318 55192
rect 7318 55136 7320 55192
rect 7264 54994 7266 55050
rect 7266 54994 7318 55050
rect 7318 54994 7320 55050
rect 7452 55729 7508 55741
rect 7452 55685 7454 55729
rect 7454 55685 7506 55729
rect 7506 55685 7508 55729
rect 7452 55543 7454 55599
rect 7454 55543 7506 55599
rect 7506 55543 7508 55599
rect 7452 55401 7454 55457
rect 7454 55401 7506 55457
rect 7506 55401 7508 55457
rect 7452 55259 7454 55315
rect 7454 55259 7506 55315
rect 7506 55259 7508 55315
rect 7452 55117 7454 55173
rect 7454 55117 7506 55173
rect 7506 55117 7508 55173
rect 7452 54975 7454 55031
rect 7454 54975 7506 55031
rect 7506 54975 7508 55031
rect 4760 54845 4762 54889
rect 4762 54845 4814 54889
rect 4814 54845 4816 54889
rect 4760 54833 4816 54845
rect 6106 54845 6108 54889
rect 6108 54845 6160 54889
rect 6160 54845 6162 54889
rect 6106 54833 6162 54845
rect 7452 54845 7454 54889
rect 7454 54845 7506 54889
rect 7506 54845 7508 54889
rect 7452 54833 7508 54845
rect 10004 55729 10060 55741
rect 10004 55685 10006 55729
rect 10006 55685 10058 55729
rect 10058 55685 10060 55729
rect 10004 55543 10006 55599
rect 10006 55543 10058 55599
rect 10058 55543 10060 55599
rect 10004 55401 10006 55457
rect 10006 55401 10058 55457
rect 10058 55401 10060 55457
rect 10004 55259 10006 55315
rect 10006 55259 10058 55315
rect 10058 55259 10060 55315
rect 10004 55117 10006 55173
rect 10006 55117 10058 55173
rect 10058 55117 10060 55173
rect 10004 54975 10006 55031
rect 10006 54975 10058 55031
rect 10058 54975 10060 55031
rect 10192 55704 10194 55760
rect 10194 55704 10246 55760
rect 10246 55704 10248 55760
rect 10192 55562 10194 55618
rect 10194 55562 10246 55618
rect 10246 55562 10248 55618
rect 10192 55420 10194 55476
rect 10194 55420 10246 55476
rect 10246 55420 10248 55476
rect 10192 55278 10194 55334
rect 10194 55278 10246 55334
rect 10246 55278 10248 55334
rect 10192 55136 10194 55192
rect 10194 55136 10246 55192
rect 10246 55136 10248 55192
rect 10192 54994 10194 55050
rect 10194 54994 10246 55050
rect 10246 54994 10248 55050
rect 10680 55704 10682 55760
rect 10682 55704 10734 55760
rect 10734 55704 10736 55760
rect 10680 55562 10682 55618
rect 10682 55562 10734 55618
rect 10734 55562 10736 55618
rect 10680 55420 10682 55476
rect 10682 55420 10734 55476
rect 10734 55420 10736 55476
rect 10680 55278 10682 55334
rect 10682 55278 10734 55334
rect 10734 55278 10736 55334
rect 10680 55136 10682 55192
rect 10682 55136 10734 55192
rect 10734 55136 10736 55192
rect 10680 54994 10682 55050
rect 10682 54994 10734 55050
rect 10734 54994 10736 55050
rect 11168 55704 11170 55760
rect 11170 55704 11222 55760
rect 11222 55704 11224 55760
rect 11168 55562 11170 55618
rect 11170 55562 11222 55618
rect 11222 55562 11224 55618
rect 11168 55420 11170 55476
rect 11170 55420 11222 55476
rect 11222 55420 11224 55476
rect 11168 55278 11170 55334
rect 11170 55278 11222 55334
rect 11222 55278 11224 55334
rect 11168 55136 11170 55192
rect 11170 55136 11222 55192
rect 11222 55136 11224 55192
rect 11168 54994 11170 55050
rect 11170 54994 11222 55050
rect 11222 54994 11224 55050
rect 11350 55729 11406 55741
rect 11350 55685 11352 55729
rect 11352 55685 11404 55729
rect 11404 55685 11406 55729
rect 11350 55543 11352 55599
rect 11352 55543 11404 55599
rect 11404 55543 11406 55599
rect 11350 55401 11352 55457
rect 11352 55401 11404 55457
rect 11404 55401 11406 55457
rect 11350 55259 11352 55315
rect 11352 55259 11404 55315
rect 11404 55259 11406 55315
rect 11350 55117 11352 55173
rect 11352 55117 11404 55173
rect 11404 55117 11406 55173
rect 11350 54975 11352 55031
rect 11352 54975 11404 55031
rect 11404 54975 11406 55031
rect 11532 55704 11534 55760
rect 11534 55704 11586 55760
rect 11586 55704 11588 55760
rect 11532 55562 11534 55618
rect 11534 55562 11586 55618
rect 11586 55562 11588 55618
rect 11532 55420 11534 55476
rect 11534 55420 11586 55476
rect 11586 55420 11588 55476
rect 11532 55278 11534 55334
rect 11534 55278 11586 55334
rect 11586 55278 11588 55334
rect 11532 55136 11534 55192
rect 11534 55136 11586 55192
rect 11586 55136 11588 55192
rect 11532 54994 11534 55050
rect 11534 54994 11586 55050
rect 11586 54994 11588 55050
rect 12020 55704 12022 55760
rect 12022 55704 12074 55760
rect 12074 55704 12076 55760
rect 12020 55562 12022 55618
rect 12022 55562 12074 55618
rect 12074 55562 12076 55618
rect 12020 55420 12022 55476
rect 12022 55420 12074 55476
rect 12074 55420 12076 55476
rect 12020 55278 12022 55334
rect 12022 55278 12074 55334
rect 12074 55278 12076 55334
rect 12020 55136 12022 55192
rect 12022 55136 12074 55192
rect 12074 55136 12076 55192
rect 12020 54994 12022 55050
rect 12022 54994 12074 55050
rect 12074 54994 12076 55050
rect 12508 55704 12510 55760
rect 12510 55704 12562 55760
rect 12562 55704 12564 55760
rect 12508 55562 12510 55618
rect 12510 55562 12562 55618
rect 12562 55562 12564 55618
rect 12508 55420 12510 55476
rect 12510 55420 12562 55476
rect 12562 55420 12564 55476
rect 12508 55278 12510 55334
rect 12510 55278 12562 55334
rect 12562 55278 12564 55334
rect 12508 55136 12510 55192
rect 12510 55136 12562 55192
rect 12562 55136 12564 55192
rect 12508 54994 12510 55050
rect 12510 54994 12562 55050
rect 12562 54994 12564 55050
rect 12696 55729 12752 55741
rect 12696 55685 12698 55729
rect 12698 55685 12750 55729
rect 12750 55685 12752 55729
rect 12696 55543 12698 55599
rect 12698 55543 12750 55599
rect 12750 55543 12752 55599
rect 12696 55401 12698 55457
rect 12698 55401 12750 55457
rect 12750 55401 12752 55457
rect 12696 55259 12698 55315
rect 12698 55259 12750 55315
rect 12750 55259 12752 55315
rect 12696 55117 12698 55173
rect 12698 55117 12750 55173
rect 12750 55117 12752 55173
rect 12696 54975 12698 55031
rect 12698 54975 12750 55031
rect 12750 54975 12752 55031
rect 10004 54845 10006 54889
rect 10006 54845 10058 54889
rect 10058 54845 10060 54889
rect 10004 54833 10060 54845
rect 11350 54845 11352 54889
rect 11352 54845 11404 54889
rect 11404 54845 11406 54889
rect 11350 54833 11406 54845
rect 12696 54845 12698 54889
rect 12698 54845 12750 54889
rect 12750 54845 12752 54889
rect 12696 54833 12752 54845
rect 1896 53394 1952 53450
rect 1896 53252 1952 53308
rect 1896 53110 1952 53166
rect 1896 52968 1952 53024
rect 4760 54104 4762 54160
rect 4762 54104 4814 54160
rect 4814 54104 4816 54160
rect 4760 53962 4762 54018
rect 4762 53962 4814 54018
rect 4814 53962 4816 54018
rect 4760 53820 4762 53876
rect 4762 53820 4814 53876
rect 4814 53820 4816 53876
rect 4760 53678 4762 53734
rect 4762 53678 4814 53734
rect 4814 53678 4816 53734
rect 4760 53536 4762 53592
rect 4762 53536 4814 53592
rect 4814 53536 4816 53592
rect 4760 53394 4762 53450
rect 4762 53394 4814 53450
rect 4814 53394 4816 53450
rect 4760 53252 4816 53308
rect 4948 54043 5004 54099
rect 4948 53901 4950 53957
rect 4950 53901 5002 53957
rect 5002 53901 5004 53957
rect 4948 53759 4950 53815
rect 4950 53759 5002 53815
rect 5002 53759 5004 53815
rect 4948 53617 4950 53673
rect 4950 53617 5002 53673
rect 5002 53617 5004 53673
rect 4948 53475 4950 53531
rect 4950 53475 5002 53531
rect 5002 53475 5004 53531
rect 4948 53333 5004 53389
rect 1896 52826 1952 52882
rect 5436 54043 5492 54099
rect 5436 53901 5438 53957
rect 5438 53901 5490 53957
rect 5490 53901 5492 53957
rect 5436 53759 5438 53815
rect 5438 53759 5490 53815
rect 5490 53759 5492 53815
rect 5436 53617 5438 53673
rect 5438 53617 5490 53673
rect 5490 53617 5492 53673
rect 5436 53475 5438 53531
rect 5438 53475 5490 53531
rect 5490 53475 5492 53531
rect 5436 53333 5492 53389
rect 5924 54043 5980 54099
rect 5924 53901 5926 53957
rect 5926 53901 5978 53957
rect 5978 53901 5980 53957
rect 5924 53759 5926 53815
rect 5926 53759 5978 53815
rect 5978 53759 5980 53815
rect 5924 53617 5926 53673
rect 5926 53617 5978 53673
rect 5978 53617 5980 53673
rect 5924 53475 5926 53531
rect 5926 53475 5978 53531
rect 5978 53475 5980 53531
rect 5924 53333 5980 53389
rect 6106 54104 6108 54160
rect 6108 54104 6160 54160
rect 6160 54104 6162 54160
rect 6106 53962 6108 54018
rect 6108 53962 6160 54018
rect 6160 53962 6162 54018
rect 6106 53820 6108 53876
rect 6108 53820 6160 53876
rect 6160 53820 6162 53876
rect 6106 53678 6108 53734
rect 6108 53678 6160 53734
rect 6160 53678 6162 53734
rect 6106 53536 6108 53592
rect 6108 53536 6160 53592
rect 6160 53536 6162 53592
rect 6106 53394 6108 53450
rect 6108 53394 6160 53450
rect 6160 53394 6162 53450
rect 6288 54043 6344 54099
rect 6288 53901 6290 53957
rect 6290 53901 6342 53957
rect 6342 53901 6344 53957
rect 6288 53759 6290 53815
rect 6290 53759 6342 53815
rect 6342 53759 6344 53815
rect 6288 53617 6290 53673
rect 6290 53617 6342 53673
rect 6342 53617 6344 53673
rect 6288 53475 6290 53531
rect 6290 53475 6342 53531
rect 6342 53475 6344 53531
rect 6288 53333 6344 53389
rect 6776 54043 6832 54099
rect 6776 53901 6778 53957
rect 6778 53901 6830 53957
rect 6830 53901 6832 53957
rect 6776 53759 6778 53815
rect 6778 53759 6830 53815
rect 6830 53759 6832 53815
rect 6776 53617 6778 53673
rect 6778 53617 6830 53673
rect 6830 53617 6832 53673
rect 6776 53475 6778 53531
rect 6778 53475 6830 53531
rect 6830 53475 6832 53531
rect 6776 53333 6832 53389
rect 6106 53252 6162 53308
rect 7264 54043 7320 54099
rect 7264 53901 7266 53957
rect 7266 53901 7318 53957
rect 7318 53901 7320 53957
rect 7264 53759 7266 53815
rect 7266 53759 7318 53815
rect 7318 53759 7320 53815
rect 7264 53617 7266 53673
rect 7266 53617 7318 53673
rect 7318 53617 7320 53673
rect 7264 53475 7266 53531
rect 7266 53475 7318 53531
rect 7318 53475 7320 53531
rect 7264 53333 7320 53389
rect 7452 54104 7454 54160
rect 7454 54104 7506 54160
rect 7506 54104 7508 54160
rect 7452 53962 7454 54018
rect 7454 53962 7506 54018
rect 7506 53962 7508 54018
rect 7452 53820 7454 53876
rect 7454 53820 7506 53876
rect 7506 53820 7508 53876
rect 7452 53678 7454 53734
rect 7454 53678 7506 53734
rect 7506 53678 7508 53734
rect 7452 53536 7454 53592
rect 7454 53536 7506 53592
rect 7506 53536 7508 53592
rect 7452 53394 7454 53450
rect 7454 53394 7506 53450
rect 7506 53394 7508 53450
rect 7452 53252 7508 53308
rect 9179 54104 9235 54160
rect 9321 54104 9377 54160
rect 9463 54104 9519 54160
rect 9179 53962 9235 54018
rect 9321 53962 9377 54018
rect 9463 53962 9519 54018
rect 9179 53820 9235 53876
rect 9321 53820 9377 53876
rect 9463 53820 9519 53876
rect 9179 53678 9235 53734
rect 9321 53678 9377 53734
rect 9463 53678 9519 53734
rect 9179 53536 9235 53592
rect 9321 53536 9377 53592
rect 9463 53536 9519 53592
rect 9179 53394 9235 53450
rect 9321 53394 9377 53450
rect 9463 53394 9519 53450
rect 9179 53252 9235 53308
rect 9321 53252 9377 53308
rect 9463 53252 9519 53308
rect 10004 54104 10006 54160
rect 10006 54104 10058 54160
rect 10058 54104 10060 54160
rect 10004 53962 10006 54018
rect 10006 53962 10058 54018
rect 10058 53962 10060 54018
rect 10004 53820 10006 53876
rect 10006 53820 10058 53876
rect 10058 53820 10060 53876
rect 10004 53678 10006 53734
rect 10006 53678 10058 53734
rect 10058 53678 10060 53734
rect 10004 53536 10006 53592
rect 10006 53536 10058 53592
rect 10058 53536 10060 53592
rect 10004 53394 10006 53450
rect 10006 53394 10058 53450
rect 10058 53394 10060 53450
rect 10192 54043 10248 54099
rect 10192 53901 10194 53957
rect 10194 53901 10246 53957
rect 10246 53901 10248 53957
rect 10192 53759 10194 53815
rect 10194 53759 10246 53815
rect 10246 53759 10248 53815
rect 10192 53617 10194 53673
rect 10194 53617 10246 53673
rect 10246 53617 10248 53673
rect 10192 53475 10194 53531
rect 10194 53475 10246 53531
rect 10246 53475 10248 53531
rect 10192 53333 10248 53389
rect 10680 54043 10736 54099
rect 10680 53901 10682 53957
rect 10682 53901 10734 53957
rect 10734 53901 10736 53957
rect 10680 53759 10682 53815
rect 10682 53759 10734 53815
rect 10734 53759 10736 53815
rect 10680 53617 10682 53673
rect 10682 53617 10734 53673
rect 10734 53617 10736 53673
rect 10680 53475 10682 53531
rect 10682 53475 10734 53531
rect 10734 53475 10736 53531
rect 10680 53333 10736 53389
rect 11168 54043 11224 54099
rect 11168 53901 11170 53957
rect 11170 53901 11222 53957
rect 11222 53901 11224 53957
rect 11168 53759 11170 53815
rect 11170 53759 11222 53815
rect 11222 53759 11224 53815
rect 11168 53617 11170 53673
rect 11170 53617 11222 53673
rect 11222 53617 11224 53673
rect 11168 53475 11170 53531
rect 11170 53475 11222 53531
rect 11222 53475 11224 53531
rect 11168 53333 11224 53389
rect 11350 54104 11352 54160
rect 11352 54104 11404 54160
rect 11404 54104 11406 54160
rect 11350 53962 11352 54018
rect 11352 53962 11404 54018
rect 11404 53962 11406 54018
rect 11350 53820 11352 53876
rect 11352 53820 11404 53876
rect 11404 53820 11406 53876
rect 11350 53678 11352 53734
rect 11352 53678 11404 53734
rect 11404 53678 11406 53734
rect 11350 53536 11352 53592
rect 11352 53536 11404 53592
rect 11404 53536 11406 53592
rect 11350 53394 11352 53450
rect 11352 53394 11404 53450
rect 11404 53394 11406 53450
rect 10004 53252 10060 53308
rect 11532 54043 11588 54099
rect 11532 53901 11534 53957
rect 11534 53901 11586 53957
rect 11586 53901 11588 53957
rect 11532 53759 11534 53815
rect 11534 53759 11586 53815
rect 11586 53759 11588 53815
rect 11532 53617 11534 53673
rect 11534 53617 11586 53673
rect 11586 53617 11588 53673
rect 11532 53475 11534 53531
rect 11534 53475 11586 53531
rect 11586 53475 11588 53531
rect 11532 53333 11588 53389
rect 12020 54043 12076 54099
rect 12020 53901 12022 53957
rect 12022 53901 12074 53957
rect 12074 53901 12076 53957
rect 12020 53759 12022 53815
rect 12022 53759 12074 53815
rect 12074 53759 12076 53815
rect 12020 53617 12022 53673
rect 12022 53617 12074 53673
rect 12074 53617 12076 53673
rect 12020 53475 12022 53531
rect 12022 53475 12074 53531
rect 12074 53475 12076 53531
rect 12020 53333 12076 53389
rect 12508 54043 12564 54099
rect 12508 53901 12510 53957
rect 12510 53901 12562 53957
rect 12562 53901 12564 53957
rect 12508 53759 12510 53815
rect 12510 53759 12562 53815
rect 12562 53759 12564 53815
rect 12508 53617 12510 53673
rect 12510 53617 12562 53673
rect 12562 53617 12564 53673
rect 12508 53475 12510 53531
rect 12510 53475 12562 53531
rect 12562 53475 12564 53531
rect 12508 53333 12564 53389
rect 12696 54104 12698 54160
rect 12698 54104 12750 54160
rect 12750 54104 12752 54160
rect 12696 53962 12698 54018
rect 12698 53962 12750 54018
rect 12750 53962 12752 54018
rect 12696 53820 12698 53876
rect 12698 53820 12750 53876
rect 12750 53820 12752 53876
rect 12696 53678 12698 53734
rect 12698 53678 12750 53734
rect 12750 53678 12752 53734
rect 12696 53536 12698 53592
rect 12698 53536 12750 53592
rect 12750 53536 12752 53592
rect 12696 53394 12698 53450
rect 12698 53394 12750 53450
rect 12750 53394 12752 53450
rect 11350 53252 11406 53308
rect 12696 53252 12752 53308
rect 9179 53110 9235 53166
rect 9321 53110 9377 53166
rect 9463 53110 9519 53166
rect 9179 52968 9235 53024
rect 9321 52968 9377 53024
rect 9463 52968 9519 53024
rect 9179 52826 9235 52882
rect 9321 52826 9377 52882
rect 9463 52826 9519 52882
rect 3618 47704 3620 47760
rect 3620 47704 3672 47760
rect 3672 47704 3674 47760
rect 3618 47562 3620 47618
rect 3620 47562 3672 47618
rect 3672 47562 3674 47618
rect 3618 47420 3620 47476
rect 3620 47420 3672 47476
rect 3672 47420 3674 47476
rect 3618 47278 3620 47334
rect 3620 47278 3672 47334
rect 3672 47278 3674 47334
rect 3618 47136 3620 47192
rect 3620 47136 3672 47192
rect 3672 47136 3674 47192
rect 3618 46994 3620 47050
rect 3620 46994 3672 47050
rect 3672 46994 3674 47050
rect 3618 46852 3620 46908
rect 3620 46852 3672 46908
rect 3672 46852 3674 46908
rect 3618 46710 3620 46766
rect 3620 46710 3672 46766
rect 3672 46710 3674 46766
rect 11584 49846 11640 49902
rect 11696 49846 11752 49902
rect 11584 49734 11640 49790
rect 11696 49734 11752 49790
rect 11584 49622 11640 49678
rect 11696 49622 11752 49678
rect 10792 49304 10794 49360
rect 10794 49304 10846 49360
rect 10846 49304 10848 49360
rect 10792 49162 10794 49218
rect 10794 49162 10846 49218
rect 10846 49162 10848 49218
rect 10792 49020 10794 49076
rect 10794 49020 10846 49076
rect 10846 49020 10848 49076
rect 10792 48878 10794 48934
rect 10794 48878 10846 48934
rect 10846 48878 10848 48934
rect 10792 48736 10794 48792
rect 10794 48736 10846 48792
rect 10846 48736 10848 48792
rect 10792 48594 10794 48650
rect 10794 48594 10846 48650
rect 10846 48594 10848 48650
rect 10792 48452 10794 48508
rect 10794 48452 10846 48508
rect 10846 48452 10848 48508
rect 10792 48310 10848 48366
rect 10434 47980 10594 48036
rect 11011 47718 11067 47744
rect 11011 47688 11013 47718
rect 11013 47688 11065 47718
rect 11065 47688 11067 47718
rect 11011 47546 11013 47602
rect 11013 47546 11065 47602
rect 11065 47546 11067 47602
rect 11011 47404 11013 47460
rect 11013 47404 11065 47460
rect 11065 47404 11067 47460
rect 11011 47262 11013 47318
rect 11013 47262 11065 47318
rect 11065 47262 11067 47318
rect 11011 47146 11013 47176
rect 11013 47146 11065 47176
rect 11065 47146 11067 47176
rect 11011 47120 11067 47146
rect 10898 44822 10954 46126
rect 11027 44822 11083 46126
rect 3618 44543 3674 44560
rect 3618 44504 3620 44543
rect 3620 44504 3672 44543
rect 3672 44504 3674 44543
rect 3618 44362 3620 44418
rect 3620 44362 3672 44418
rect 3672 44362 3674 44418
rect 3618 44220 3620 44276
rect 3620 44220 3672 44276
rect 3672 44220 3674 44276
rect 3618 44078 3620 44134
rect 3620 44078 3672 44134
rect 3672 44078 3674 44134
rect 3618 43936 3620 43992
rect 3620 43936 3672 43992
rect 3672 43936 3674 43992
rect 3618 43794 3620 43850
rect 3620 43794 3672 43850
rect 3672 43794 3674 43850
rect 3618 43652 3620 43708
rect 3620 43652 3672 43708
rect 3672 43652 3674 43708
rect 3618 43510 3620 43566
rect 3620 43510 3672 43566
rect 3672 43510 3674 43566
rect 3618 43368 3620 43424
rect 3620 43368 3672 43424
rect 3672 43368 3674 43424
rect 3618 43243 3620 43282
rect 3620 43243 3672 43282
rect 3672 43243 3674 43282
rect 3618 43226 3674 43243
rect 3618 42943 3674 42960
rect 3618 42904 3620 42943
rect 3620 42904 3672 42943
rect 3672 42904 3674 42943
rect 3618 42762 3620 42818
rect 3620 42762 3672 42818
rect 3672 42762 3674 42818
rect 3618 42620 3620 42676
rect 3620 42620 3672 42676
rect 3672 42620 3674 42676
rect 3618 42478 3620 42534
rect 3620 42478 3672 42534
rect 3672 42478 3674 42534
rect 3618 42336 3620 42392
rect 3620 42336 3672 42392
rect 3672 42336 3674 42392
rect 3618 42194 3620 42250
rect 3620 42194 3672 42250
rect 3672 42194 3674 42250
rect 3618 42052 3620 42108
rect 3620 42052 3672 42108
rect 3672 42052 3674 42108
rect 3618 41910 3620 41966
rect 3620 41910 3672 41966
rect 3672 41910 3674 41966
rect 3618 41768 3620 41824
rect 3620 41768 3672 41824
rect 3672 41768 3674 41824
rect 3618 41643 3620 41682
rect 3620 41643 3672 41682
rect 3672 41643 3674 41682
rect 3618 41626 3674 41643
rect 1846 41070 1902 41072
rect 1988 41070 2044 41072
rect 2130 41070 2186 41072
rect 2272 41070 2328 41072
rect 2414 41070 2470 41072
rect 2556 41070 2612 41072
rect 2698 41070 2754 41072
rect 2840 41070 2896 41072
rect 2982 41070 3038 41072
rect 3124 41070 3180 41072
rect 3266 41070 3322 41072
rect 3408 41070 3464 41072
rect 3550 41070 3606 41072
rect 1846 41018 1848 41070
rect 1848 41018 1902 41070
rect 1988 41018 2044 41070
rect 2130 41018 2186 41070
rect 2272 41018 2328 41070
rect 2414 41018 2470 41070
rect 2556 41018 2612 41070
rect 2698 41018 2754 41070
rect 2840 41018 2896 41070
rect 2982 41018 3038 41070
rect 3124 41018 3180 41070
rect 3266 41018 3322 41070
rect 3408 41018 3464 41070
rect 3550 41018 3606 41070
rect 1846 41016 1902 41018
rect 1988 41016 2044 41018
rect 2130 41016 2186 41018
rect 2272 41016 2328 41018
rect 2414 41016 2470 41018
rect 2556 41016 2612 41018
rect 2698 41016 2754 41018
rect 2840 41016 2896 41018
rect 2982 41016 3038 41018
rect 3124 41016 3180 41018
rect 3266 41016 3322 41018
rect 3408 41016 3464 41018
rect 3550 41016 3606 41018
rect 3692 41016 3748 41072
rect 1781 39704 1783 39760
rect 1783 39704 1835 39760
rect 1835 39704 1837 39760
rect 1781 39562 1783 39618
rect 1783 39562 1835 39618
rect 1835 39562 1837 39618
rect 1781 39420 1783 39476
rect 1783 39420 1835 39476
rect 1835 39420 1837 39476
rect 1781 39278 1783 39334
rect 1783 39278 1835 39334
rect 1835 39278 1837 39334
rect 1781 39136 1837 39192
rect 2367 40260 2423 40316
rect 2509 40314 2565 40316
rect 2651 40314 2707 40316
rect 2793 40314 2849 40316
rect 2935 40314 2991 40316
rect 3077 40314 3133 40316
rect 3219 40314 3275 40316
rect 3361 40314 3417 40316
rect 3503 40314 3559 40316
rect 3645 40314 3701 40316
rect 3787 40314 3843 40316
rect 3929 40314 3985 40316
rect 4071 40314 4127 40316
rect 4213 40314 4269 40316
rect 4355 40314 4411 40316
rect 2509 40262 2565 40314
rect 2651 40262 2707 40314
rect 2793 40262 2849 40314
rect 2935 40262 2991 40314
rect 3077 40262 3133 40314
rect 3219 40262 3275 40314
rect 3361 40262 3417 40314
rect 3503 40262 3559 40314
rect 3645 40262 3701 40314
rect 3787 40262 3843 40314
rect 3929 40262 3985 40314
rect 4071 40262 4127 40314
rect 4213 40262 4269 40314
rect 4355 40262 4411 40314
rect 2509 40260 2565 40262
rect 2651 40260 2707 40262
rect 2793 40260 2849 40262
rect 2935 40260 2991 40262
rect 3077 40260 3133 40262
rect 3219 40260 3275 40262
rect 3361 40260 3417 40262
rect 3503 40260 3559 40262
rect 3645 40260 3701 40262
rect 3787 40260 3843 40262
rect 3929 40260 3985 40262
rect 4071 40260 4127 40262
rect 4213 40260 4269 40262
rect 4355 40260 4411 40262
rect 4497 40260 4553 40316
rect 5093 39758 5149 39760
rect 5093 39704 5095 39758
rect 5095 39704 5147 39758
rect 5147 39704 5149 39758
rect 5093 39562 5095 39618
rect 5095 39562 5147 39618
rect 5147 39562 5149 39618
rect 5093 39420 5095 39476
rect 5095 39420 5147 39476
rect 5147 39420 5149 39476
rect 5093 39278 5095 39334
rect 5095 39278 5147 39334
rect 5147 39278 5149 39334
rect 5093 39186 5095 39192
rect 5095 39186 5147 39192
rect 5147 39186 5149 39192
rect 5093 39136 5149 39186
rect 6059 39698 6061 39754
rect 6061 39698 6113 39754
rect 6113 39698 6115 39754
rect 6059 39556 6061 39612
rect 6061 39556 6113 39612
rect 6113 39556 6115 39612
rect 6059 39414 6061 39470
rect 6061 39414 6113 39470
rect 6113 39414 6115 39470
rect 6059 39272 6061 39328
rect 6061 39272 6113 39328
rect 6113 39272 6115 39328
rect 6059 39130 6061 39186
rect 6061 39130 6113 39186
rect 6113 39130 6115 39186
rect 7025 39758 7081 39760
rect 7025 39704 7027 39758
rect 7027 39704 7079 39758
rect 7079 39704 7081 39758
rect 7025 39562 7027 39618
rect 7027 39562 7079 39618
rect 7079 39562 7081 39618
rect 7025 39420 7027 39476
rect 7027 39420 7079 39476
rect 7079 39420 7081 39476
rect 7025 39278 7027 39334
rect 7027 39278 7079 39334
rect 7079 39278 7081 39334
rect 7025 39186 7027 39192
rect 7027 39186 7079 39192
rect 7079 39186 7081 39192
rect 7025 39136 7081 39186
rect 6059 38988 6061 39044
rect 6061 38988 6113 39044
rect 6113 38988 6115 39044
rect 6059 38846 6061 38902
rect 6061 38846 6113 38902
rect 6113 38846 6115 38902
rect 6059 38704 6115 38760
rect 56 38143 112 38167
rect 56 38111 58 38143
rect 58 38111 110 38143
rect 110 38111 112 38143
rect 56 37969 58 38025
rect 58 37969 110 38025
rect 110 37969 112 38025
rect 56 37827 58 37883
rect 58 37827 110 37883
rect 110 37827 112 37883
rect 56 37685 58 37741
rect 58 37685 110 37741
rect 110 37685 112 37741
rect 56 37543 58 37599
rect 58 37543 110 37599
rect 110 37543 112 37599
rect 56 37401 58 37457
rect 58 37401 110 37457
rect 110 37401 112 37457
rect 56 37259 58 37315
rect 58 37259 110 37315
rect 110 37259 112 37315
rect 56 37117 58 37173
rect 58 37117 110 37173
rect 110 37117 112 37173
rect 56 36975 58 37031
rect 58 36975 110 37031
rect 110 36975 112 37031
rect 56 36843 58 36889
rect 58 36843 110 36889
rect 110 36843 112 36889
rect 56 36833 112 36843
rect 734 38104 790 38160
rect 734 37962 790 38018
rect 734 37820 790 37876
rect 734 37678 790 37734
rect 734 37536 790 37592
rect 876 38104 932 38160
rect 1018 38104 1074 38160
rect 876 37962 932 38018
rect 1018 37962 1074 38018
rect 876 37820 932 37876
rect 1018 37820 1074 37876
rect 876 37678 932 37734
rect 1018 37678 1074 37734
rect 876 37536 932 37592
rect 1018 37536 1074 37592
rect 734 37394 790 37450
rect 876 37394 932 37450
rect 1018 37394 1074 37450
rect 734 37252 790 37308
rect 876 37252 932 37308
rect 1018 37252 1074 37308
rect 734 37110 790 37166
rect 876 37110 932 37166
rect 1018 37110 1074 37166
rect 734 36968 790 37024
rect 876 36968 932 37024
rect 1018 36968 1074 37024
rect 734 36826 790 36882
rect 876 36826 932 36882
rect 1018 36826 1074 36882
rect 175 36492 231 36548
rect 317 36492 373 36548
rect 175 36350 231 36406
rect 317 36350 373 36406
rect 175 36208 231 36264
rect 317 36208 373 36264
rect 175 36066 231 36122
rect 317 36066 373 36122
rect 175 35924 231 35980
rect 317 35924 373 35980
rect 175 35782 231 35838
rect 317 35782 373 35838
rect 175 35640 231 35696
rect 317 35640 373 35696
rect 175 35498 231 35554
rect 317 35498 373 35554
rect 175 35356 231 35412
rect 317 35356 373 35412
rect 175 35214 231 35270
rect 317 35214 373 35270
rect 175 35072 231 35128
rect 317 35072 373 35128
rect 175 34930 231 34986
rect 317 34930 373 34986
rect 175 34788 231 34844
rect 317 34788 373 34844
rect 175 34646 231 34702
rect 317 34646 373 34702
rect 175 34504 231 34560
rect 317 34504 373 34560
rect 175 34362 231 34418
rect 317 34362 373 34418
rect 175 34220 231 34276
rect 317 34220 373 34276
rect 175 34078 231 34134
rect 317 34078 373 34134
rect 496 35946 552 35987
rect 496 35931 498 35946
rect 498 35931 550 35946
rect 550 35931 552 35946
rect 496 35789 498 35845
rect 498 35789 550 35845
rect 550 35789 552 35845
rect 496 35647 498 35703
rect 498 35647 550 35703
rect 550 35647 552 35703
rect 496 35505 498 35561
rect 498 35505 550 35561
rect 550 35505 552 35561
rect 496 35363 498 35419
rect 498 35363 550 35419
rect 550 35363 552 35419
rect 496 35221 498 35277
rect 498 35221 550 35277
rect 550 35221 552 35277
rect 496 35079 498 35135
rect 498 35079 550 35135
rect 550 35079 552 35135
rect 496 34937 498 34993
rect 498 34937 550 34993
rect 550 34937 552 34993
rect 496 34795 498 34851
rect 498 34795 550 34851
rect 550 34795 552 34851
rect 496 34653 498 34709
rect 498 34653 550 34709
rect 550 34653 552 34709
rect 496 34511 498 34567
rect 498 34511 550 34567
rect 550 34511 552 34567
rect 734 35946 790 35982
rect 734 35926 736 35946
rect 736 35926 788 35946
rect 788 35926 790 35946
rect 734 35784 736 35840
rect 736 35784 788 35840
rect 788 35784 790 35840
rect 734 35642 736 35698
rect 736 35642 788 35698
rect 788 35642 790 35698
rect 734 35500 736 35556
rect 736 35500 788 35556
rect 788 35500 790 35556
rect 734 35358 736 35414
rect 736 35358 788 35414
rect 788 35358 790 35414
rect 734 35216 736 35272
rect 736 35216 788 35272
rect 788 35216 790 35272
rect 734 35074 736 35130
rect 736 35074 788 35130
rect 788 35074 790 35130
rect 734 34932 736 34988
rect 736 34932 788 34988
rect 788 34932 790 34988
rect 734 34790 736 34846
rect 736 34790 788 34846
rect 788 34790 790 34846
rect 734 34648 736 34704
rect 736 34648 788 34704
rect 788 34648 790 34704
rect 734 34542 736 34562
rect 736 34542 788 34562
rect 788 34542 790 34562
rect 734 34506 790 34542
rect 496 34369 498 34425
rect 498 34369 550 34425
rect 550 34369 552 34425
rect 496 34227 498 34283
rect 498 34227 550 34283
rect 550 34227 552 34283
rect 496 34126 498 34141
rect 498 34126 550 34141
rect 550 34126 552 34141
rect 496 34085 552 34126
rect 175 33936 231 33992
rect 317 33936 373 33992
rect 175 33794 231 33850
rect 317 33794 373 33850
rect 175 33652 231 33708
rect 317 33652 373 33708
rect 496 33292 498 33348
rect 498 33292 550 33348
rect 550 33292 552 33348
rect 496 33150 498 33206
rect 498 33150 550 33206
rect 550 33150 552 33206
rect 496 33008 498 33064
rect 498 33008 550 33064
rect 550 33008 552 33064
rect 496 32866 498 32922
rect 498 32866 550 32922
rect 550 32866 552 32922
rect 6059 38104 6061 38160
rect 6061 38104 6113 38160
rect 6113 38104 6115 38160
rect 6059 37962 6061 38018
rect 6061 37962 6113 38018
rect 6113 37962 6115 38018
rect 6059 37820 6061 37876
rect 6061 37820 6113 37876
rect 6113 37820 6115 37876
rect 6059 37678 6061 37734
rect 6061 37678 6113 37734
rect 6113 37678 6115 37734
rect 6059 37536 6061 37592
rect 6061 37536 6113 37592
rect 6113 37536 6115 37592
rect 6059 37394 6115 37450
rect 6059 37252 6115 37308
rect 6059 37110 6115 37166
rect 6059 36968 6115 37024
rect 6059 36826 6115 36882
rect 3102 35946 3158 35982
rect 3102 35926 3104 35946
rect 3104 35926 3156 35946
rect 3156 35926 3158 35946
rect 3102 35784 3104 35840
rect 3104 35784 3156 35840
rect 3156 35784 3158 35840
rect 3102 35642 3104 35698
rect 3104 35642 3156 35698
rect 3156 35642 3158 35698
rect 3102 35500 3104 35556
rect 3104 35500 3156 35556
rect 3156 35500 3158 35556
rect 3102 35358 3104 35414
rect 3104 35358 3156 35414
rect 3156 35358 3158 35414
rect 3102 35216 3104 35272
rect 3104 35216 3156 35272
rect 3156 35216 3158 35272
rect 3102 35074 3104 35130
rect 3104 35074 3156 35130
rect 3156 35074 3158 35130
rect 3102 34932 3104 34988
rect 3104 34932 3156 34988
rect 3156 34932 3158 34988
rect 3102 34790 3104 34846
rect 3104 34790 3156 34846
rect 3156 34790 3158 34846
rect 3102 34648 3104 34704
rect 3104 34648 3156 34704
rect 3156 34648 3158 34704
rect 3102 34542 3104 34562
rect 3104 34542 3156 34562
rect 3156 34542 3158 34562
rect 3102 34506 3158 34542
rect 4000 36030 4056 36086
rect 4000 35888 4002 35944
rect 4002 35888 4054 35944
rect 4054 35888 4056 35944
rect 4000 35746 4002 35802
rect 4002 35746 4054 35802
rect 4054 35746 4056 35802
rect 4000 35604 4002 35660
rect 4002 35604 4054 35660
rect 4054 35604 4056 35660
rect 4000 35462 4002 35518
rect 4002 35462 4054 35518
rect 4054 35462 4056 35518
rect 4000 35320 4002 35376
rect 4002 35320 4054 35376
rect 4054 35320 4056 35376
rect 4000 35178 4002 35234
rect 4002 35178 4054 35234
rect 4054 35178 4056 35234
rect 4000 35036 4002 35092
rect 4002 35036 4054 35092
rect 4054 35036 4056 35092
rect 4000 34894 4002 34950
rect 4002 34894 4054 34950
rect 4054 34894 4056 34950
rect 4000 34752 4002 34808
rect 4002 34752 4054 34808
rect 4054 34752 4056 34808
rect 4000 34610 4002 34666
rect 4002 34610 4054 34666
rect 4054 34610 4056 34666
rect 4000 34468 4002 34524
rect 4002 34468 4054 34524
rect 4054 34468 4056 34524
rect 4000 34326 4002 34382
rect 4002 34326 4054 34382
rect 4054 34326 4056 34382
rect 4898 35946 4954 35982
rect 4898 35926 4900 35946
rect 4900 35926 4952 35946
rect 4952 35926 4954 35946
rect 4898 35784 4900 35840
rect 4900 35784 4952 35840
rect 4952 35784 4954 35840
rect 4898 35642 4900 35698
rect 4900 35642 4952 35698
rect 4952 35642 4954 35698
rect 4898 35500 4900 35556
rect 4900 35500 4952 35556
rect 4952 35500 4954 35556
rect 4898 35358 4900 35414
rect 4900 35358 4952 35414
rect 4952 35358 4954 35414
rect 4898 35216 4900 35272
rect 4900 35216 4952 35272
rect 4952 35216 4954 35272
rect 4898 35074 4900 35130
rect 4900 35074 4952 35130
rect 4952 35074 4954 35130
rect 4898 34932 4900 34988
rect 4900 34932 4952 34988
rect 4952 34932 4954 34988
rect 4898 34790 4900 34846
rect 4900 34790 4952 34846
rect 4952 34790 4954 34846
rect 4898 34648 4900 34704
rect 4900 34648 4952 34704
rect 4952 34648 4954 34704
rect 4898 34542 4900 34562
rect 4900 34542 4952 34562
rect 4952 34542 4954 34562
rect 4898 34506 4954 34542
rect 4000 34184 4002 34240
rect 4002 34184 4054 34240
rect 4054 34184 4056 34240
rect 4000 34042 4002 34098
rect 4002 34042 4054 34098
rect 4054 34042 4056 34098
rect 4000 33900 4002 33956
rect 4002 33900 4054 33956
rect 4054 33900 4056 33956
rect 4000 33758 4002 33814
rect 4002 33758 4054 33814
rect 4054 33758 4056 33814
rect 4000 33616 4002 33672
rect 4002 33616 4054 33672
rect 4054 33616 4056 33672
rect 496 32724 498 32780
rect 498 32724 550 32780
rect 550 32724 552 32780
rect 4000 32849 4056 32905
rect 4000 32707 4002 32763
rect 4002 32707 4054 32763
rect 4054 32707 4056 32763
rect 496 32582 498 32638
rect 498 32582 550 32638
rect 550 32582 552 32638
rect 496 32440 498 32496
rect 498 32440 550 32496
rect 550 32440 552 32496
rect 496 32298 498 32354
rect 498 32298 550 32354
rect 550 32298 552 32354
rect 496 32156 498 32212
rect 498 32156 550 32212
rect 550 32156 552 32212
rect 496 32014 498 32070
rect 498 32014 550 32070
rect 550 32014 552 32070
rect 496 31872 498 31928
rect 498 31872 550 31928
rect 550 31872 552 31928
rect 496 31730 498 31786
rect 498 31730 550 31786
rect 550 31730 552 31786
rect 496 31588 498 31644
rect 498 31588 550 31644
rect 550 31588 552 31644
rect 496 31446 498 31502
rect 498 31446 550 31502
rect 550 31446 552 31502
rect 496 31304 498 31360
rect 498 31304 550 31360
rect 550 31304 552 31360
rect 496 31162 498 31218
rect 498 31162 550 31218
rect 550 31162 552 31218
rect 496 31020 498 31076
rect 498 31020 550 31076
rect 550 31020 552 31076
rect 496 30878 498 30934
rect 498 30878 550 30934
rect 550 30878 552 30934
rect 496 30736 498 30792
rect 498 30736 550 30792
rect 550 30736 552 30792
rect 496 30594 498 30650
rect 498 30594 550 30650
rect 550 30594 552 30650
rect 496 30452 498 30508
rect 498 30452 550 30508
rect 550 30452 552 30508
rect 978 32690 1034 32692
rect 978 32636 980 32690
rect 980 32636 1032 32690
rect 1032 32636 1034 32690
rect 978 32494 980 32550
rect 980 32494 1032 32550
rect 1032 32494 1034 32550
rect 978 32352 980 32408
rect 980 32352 1032 32408
rect 1032 32352 1034 32408
rect 978 32210 980 32266
rect 980 32210 1032 32266
rect 1032 32210 1034 32266
rect 978 32068 980 32124
rect 980 32068 1032 32124
rect 1032 32068 1034 32124
rect 978 31926 980 31982
rect 980 31926 1032 31982
rect 1032 31926 1034 31982
rect 978 31784 980 31840
rect 980 31784 1032 31840
rect 1032 31784 1034 31840
rect 978 31642 980 31698
rect 980 31642 1032 31698
rect 1032 31642 1034 31698
rect 978 31500 980 31556
rect 980 31500 1032 31556
rect 1032 31500 1034 31556
rect 978 31358 980 31414
rect 980 31358 1032 31414
rect 1032 31358 1034 31414
rect 978 31216 980 31272
rect 980 31216 1032 31272
rect 1032 31216 1034 31272
rect 978 31074 980 31130
rect 980 31074 1032 31130
rect 1032 31074 1034 31130
rect 978 30932 980 30988
rect 980 30932 1032 30988
rect 1032 30932 1034 30988
rect 978 30790 980 30846
rect 980 30790 1032 30846
rect 1032 30790 1034 30846
rect 978 30648 980 30704
rect 980 30648 1032 30704
rect 1032 30648 1034 30704
rect 2370 32690 2426 32692
rect 2370 32636 2372 32690
rect 2372 32636 2424 32690
rect 2424 32636 2426 32690
rect 2370 32494 2372 32550
rect 2372 32494 2424 32550
rect 2424 32494 2426 32550
rect 2370 32352 2372 32408
rect 2372 32352 2424 32408
rect 2424 32352 2426 32408
rect 2370 32210 2372 32266
rect 2372 32210 2424 32266
rect 2424 32210 2426 32266
rect 2370 32068 2372 32124
rect 2372 32068 2424 32124
rect 2424 32068 2426 32124
rect 2370 31926 2372 31982
rect 2372 31926 2424 31982
rect 2424 31926 2426 31982
rect 2370 31784 2372 31840
rect 2372 31784 2424 31840
rect 2424 31784 2426 31840
rect 2370 31642 2372 31698
rect 2372 31642 2424 31698
rect 2424 31642 2426 31698
rect 2370 31500 2372 31556
rect 2372 31500 2424 31556
rect 2424 31500 2426 31556
rect 2370 31358 2372 31414
rect 2372 31358 2424 31414
rect 2424 31358 2426 31414
rect 2370 31216 2372 31272
rect 2372 31216 2424 31272
rect 2424 31216 2426 31272
rect 2370 31074 2372 31130
rect 2372 31074 2424 31130
rect 2424 31074 2426 31130
rect 2370 30932 2372 30988
rect 2372 30932 2424 30988
rect 2424 30932 2426 30988
rect 2370 30790 2372 30846
rect 2372 30790 2424 30846
rect 2424 30790 2426 30846
rect 978 30506 980 30562
rect 980 30506 1032 30562
rect 1032 30506 1034 30562
rect 2370 30648 2372 30704
rect 2372 30648 2424 30704
rect 2424 30648 2426 30704
rect 2370 30506 2372 30562
rect 2372 30506 2424 30562
rect 2424 30506 2426 30562
rect 2786 32690 2842 32692
rect 2786 32636 2788 32690
rect 2788 32636 2840 32690
rect 2840 32636 2842 32690
rect 2786 32494 2788 32550
rect 2788 32494 2840 32550
rect 2840 32494 2842 32550
rect 2786 32352 2788 32408
rect 2788 32352 2840 32408
rect 2840 32352 2842 32408
rect 2786 32210 2788 32266
rect 2788 32210 2840 32266
rect 2840 32210 2842 32266
rect 2786 32068 2788 32124
rect 2788 32068 2840 32124
rect 2840 32068 2842 32124
rect 2786 31926 2788 31982
rect 2788 31926 2840 31982
rect 2840 31926 2842 31982
rect 2786 31784 2788 31840
rect 2788 31784 2840 31840
rect 2840 31784 2842 31840
rect 2786 31642 2788 31698
rect 2788 31642 2840 31698
rect 2840 31642 2842 31698
rect 2786 31500 2788 31556
rect 2788 31500 2840 31556
rect 2840 31500 2842 31556
rect 2786 31358 2788 31414
rect 2788 31358 2840 31414
rect 2840 31358 2842 31414
rect 2786 31216 2788 31272
rect 2788 31216 2840 31272
rect 2840 31216 2842 31272
rect 2786 31074 2788 31130
rect 2788 31074 2840 31130
rect 2840 31074 2842 31130
rect 3274 32690 3330 32693
rect 3274 32637 3276 32690
rect 3276 32637 3328 32690
rect 3328 32637 3330 32690
rect 3274 32495 3276 32551
rect 3276 32495 3328 32551
rect 3328 32495 3330 32551
rect 3274 32353 3276 32409
rect 3276 32353 3328 32409
rect 3328 32353 3330 32409
rect 3274 32211 3276 32267
rect 3276 32211 3328 32267
rect 3328 32211 3330 32267
rect 3274 32069 3276 32125
rect 3276 32069 3328 32125
rect 3328 32069 3330 32125
rect 3274 31927 3276 31983
rect 3276 31927 3328 31983
rect 3328 31927 3330 31983
rect 3274 31785 3276 31841
rect 3276 31785 3328 31841
rect 3328 31785 3330 31841
rect 3274 31643 3276 31699
rect 3276 31643 3328 31699
rect 3328 31643 3330 31699
rect 3274 31501 3276 31557
rect 3276 31501 3328 31557
rect 3328 31501 3330 31557
rect 3274 31359 3276 31415
rect 3276 31359 3328 31415
rect 3328 31359 3330 31415
rect 3274 31217 3276 31273
rect 3276 31217 3328 31273
rect 3328 31217 3330 31273
rect 3274 31078 3276 31131
rect 3276 31078 3328 31131
rect 3328 31078 3330 31131
rect 3274 31075 3330 31078
rect 3762 32640 3818 32642
rect 3762 32586 3764 32640
rect 3764 32586 3816 32640
rect 3816 32586 3818 32640
rect 3762 32444 3764 32500
rect 3764 32444 3816 32500
rect 3816 32444 3818 32500
rect 3762 32302 3764 32358
rect 3764 32302 3816 32358
rect 3816 32302 3818 32358
rect 3762 32160 3764 32216
rect 3764 32160 3816 32216
rect 3816 32160 3818 32216
rect 3762 32018 3764 32074
rect 3764 32018 3816 32074
rect 3816 32018 3818 32074
rect 3762 31876 3764 31932
rect 3764 31876 3816 31932
rect 3816 31876 3818 31932
rect 3762 31734 3764 31790
rect 3764 31734 3816 31790
rect 3816 31734 3818 31790
rect 3762 31592 3764 31648
rect 3764 31592 3816 31648
rect 3816 31592 3818 31648
rect 3762 31450 3764 31506
rect 3764 31450 3816 31506
rect 3816 31450 3818 31506
rect 3762 31308 3764 31364
rect 3764 31308 3816 31364
rect 3816 31308 3818 31364
rect 3762 31166 3764 31222
rect 3764 31166 3816 31222
rect 3816 31166 3818 31222
rect 3762 31028 3764 31080
rect 3764 31028 3816 31080
rect 3816 31028 3818 31080
rect 3762 31024 3818 31028
rect 4000 32565 4002 32621
rect 4002 32565 4054 32621
rect 4054 32565 4056 32621
rect 4000 32423 4002 32479
rect 4002 32423 4054 32479
rect 4054 32423 4056 32479
rect 4000 32281 4002 32337
rect 4002 32281 4054 32337
rect 4054 32281 4056 32337
rect 4000 32139 4002 32195
rect 4002 32139 4054 32195
rect 4054 32139 4056 32195
rect 4000 31997 4002 32053
rect 4002 31997 4054 32053
rect 4054 31997 4056 32053
rect 4000 31855 4002 31911
rect 4002 31855 4054 31911
rect 4054 31855 4056 31911
rect 4000 31713 4002 31769
rect 4002 31713 4054 31769
rect 4054 31713 4056 31769
rect 4000 31571 4002 31627
rect 4002 31571 4054 31627
rect 4054 31571 4056 31627
rect 4000 31429 4002 31485
rect 4002 31429 4054 31485
rect 4054 31429 4056 31485
rect 4000 31287 4002 31343
rect 4002 31287 4054 31343
rect 4054 31287 4056 31343
rect 4000 31145 4002 31201
rect 4002 31145 4054 31201
rect 4054 31145 4056 31201
rect 4000 31005 4002 31059
rect 4002 31005 4054 31059
rect 4054 31005 4056 31059
rect 4000 31003 4056 31005
rect 4238 32640 4294 32642
rect 4238 32586 4240 32640
rect 4240 32586 4292 32640
rect 4292 32586 4294 32640
rect 4238 32444 4240 32500
rect 4240 32444 4292 32500
rect 4292 32444 4294 32500
rect 4238 32302 4240 32358
rect 4240 32302 4292 32358
rect 4292 32302 4294 32358
rect 4238 32160 4240 32216
rect 4240 32160 4292 32216
rect 4292 32160 4294 32216
rect 4238 32018 4240 32074
rect 4240 32018 4292 32074
rect 4292 32018 4294 32074
rect 4238 31876 4240 31932
rect 4240 31876 4292 31932
rect 4292 31876 4294 31932
rect 4238 31734 4240 31790
rect 4240 31734 4292 31790
rect 4292 31734 4294 31790
rect 4238 31592 4240 31648
rect 4240 31592 4292 31648
rect 4292 31592 4294 31648
rect 4238 31450 4240 31506
rect 4240 31450 4292 31506
rect 4292 31450 4294 31506
rect 4238 31308 4240 31364
rect 4240 31308 4292 31364
rect 4292 31308 4294 31364
rect 4238 31166 4240 31222
rect 4240 31166 4292 31222
rect 4292 31166 4294 31222
rect 4238 31028 4240 31080
rect 4240 31028 4292 31080
rect 4292 31028 4294 31080
rect 4238 31024 4294 31028
rect 4726 32690 4782 32693
rect 4726 32637 4728 32690
rect 4728 32637 4780 32690
rect 4780 32637 4782 32690
rect 4726 32495 4728 32551
rect 4728 32495 4780 32551
rect 4780 32495 4782 32551
rect 4726 32353 4728 32409
rect 4728 32353 4780 32409
rect 4780 32353 4782 32409
rect 4726 32211 4728 32267
rect 4728 32211 4780 32267
rect 4780 32211 4782 32267
rect 4726 32069 4728 32125
rect 4728 32069 4780 32125
rect 4780 32069 4782 32125
rect 4726 31927 4728 31983
rect 4728 31927 4780 31983
rect 4780 31927 4782 31983
rect 4726 31785 4728 31841
rect 4728 31785 4780 31841
rect 4780 31785 4782 31841
rect 4726 31643 4728 31699
rect 4728 31643 4780 31699
rect 4780 31643 4782 31699
rect 4726 31501 4728 31557
rect 4728 31501 4780 31557
rect 4780 31501 4782 31557
rect 4726 31359 4728 31415
rect 4728 31359 4780 31415
rect 4780 31359 4782 31415
rect 4726 31217 4728 31273
rect 4728 31217 4780 31273
rect 4780 31217 4782 31273
rect 4726 31078 4728 31131
rect 4728 31078 4780 31131
rect 4780 31078 4782 31131
rect 4726 31075 4782 31078
rect 5214 32690 5270 32693
rect 5214 32637 5216 32690
rect 5216 32637 5268 32690
rect 5268 32637 5270 32690
rect 5214 32495 5216 32551
rect 5216 32495 5268 32551
rect 5268 32495 5270 32551
rect 5214 32353 5216 32409
rect 5216 32353 5268 32409
rect 5268 32353 5270 32409
rect 5214 32211 5216 32267
rect 5216 32211 5268 32267
rect 5268 32211 5270 32267
rect 5214 32069 5216 32125
rect 5216 32069 5268 32125
rect 5268 32069 5270 32125
rect 5214 31927 5216 31983
rect 5216 31927 5268 31983
rect 5268 31927 5270 31983
rect 5214 31785 5216 31841
rect 5216 31785 5268 31841
rect 5268 31785 5270 31841
rect 5214 31643 5216 31699
rect 5216 31643 5268 31699
rect 5268 31643 5270 31699
rect 5214 31501 5216 31557
rect 5216 31501 5268 31557
rect 5268 31501 5270 31557
rect 5214 31359 5216 31415
rect 5216 31359 5268 31415
rect 5268 31359 5270 31415
rect 5214 31217 5216 31273
rect 5216 31217 5268 31273
rect 5268 31217 5270 31273
rect 5214 31078 5216 31131
rect 5216 31078 5268 31131
rect 5268 31078 5270 31131
rect 5214 31075 5270 31078
rect 5630 32690 5686 32693
rect 5630 32637 5632 32690
rect 5632 32637 5684 32690
rect 5684 32637 5686 32690
rect 5630 32495 5632 32551
rect 5632 32495 5684 32551
rect 5684 32495 5686 32551
rect 5630 32353 5632 32409
rect 5632 32353 5684 32409
rect 5684 32353 5686 32409
rect 5630 32211 5632 32267
rect 5632 32211 5684 32267
rect 5684 32211 5686 32267
rect 5630 32069 5632 32125
rect 5632 32069 5684 32125
rect 5684 32069 5686 32125
rect 5630 31927 5632 31983
rect 5632 31927 5684 31983
rect 5684 31927 5686 31983
rect 5630 31785 5632 31841
rect 5632 31785 5684 31841
rect 5684 31785 5686 31841
rect 5630 31643 5632 31699
rect 5632 31643 5684 31699
rect 5684 31643 5686 31699
rect 5630 31501 5632 31557
rect 5632 31501 5684 31557
rect 5684 31501 5686 31557
rect 5630 31359 5632 31415
rect 5632 31359 5684 31415
rect 5684 31359 5686 31415
rect 5630 31217 5632 31273
rect 5632 31217 5684 31273
rect 5684 31217 5686 31273
rect 5630 31078 5632 31131
rect 5632 31078 5684 31131
rect 5684 31078 5686 31131
rect 5630 31075 5686 31078
rect 7022 32690 7078 32692
rect 7022 32636 7024 32690
rect 7024 32636 7076 32690
rect 7076 32636 7078 32690
rect 7022 32494 7024 32550
rect 7024 32494 7076 32550
rect 7076 32494 7078 32550
rect 7022 32352 7024 32408
rect 7024 32352 7076 32408
rect 7076 32352 7078 32408
rect 7022 32210 7024 32266
rect 7024 32210 7076 32266
rect 7076 32210 7078 32266
rect 7022 32068 7024 32124
rect 7024 32068 7076 32124
rect 7076 32068 7078 32124
rect 7022 31926 7024 31982
rect 7024 31926 7076 31982
rect 7076 31926 7078 31982
rect 7022 31784 7024 31840
rect 7024 31784 7076 31840
rect 7076 31784 7078 31840
rect 7022 31642 7024 31698
rect 7024 31642 7076 31698
rect 7076 31642 7078 31698
rect 7022 31500 7024 31556
rect 7024 31500 7076 31556
rect 7076 31500 7078 31556
rect 7022 31358 7024 31414
rect 7024 31358 7076 31414
rect 7076 31358 7078 31414
rect 7022 31216 7024 31272
rect 7024 31216 7076 31272
rect 7076 31216 7078 31272
rect 7022 31074 7024 31130
rect 7024 31074 7076 31130
rect 7076 31074 7078 31130
rect 2786 30932 2788 30988
rect 2788 30932 2840 30988
rect 2840 30932 2842 30988
rect 7022 30932 7024 30988
rect 7024 30932 7076 30988
rect 7076 30932 7078 30988
rect 2786 30790 2788 30846
rect 2788 30790 2840 30846
rect 2840 30790 2842 30846
rect 2786 30648 2788 30704
rect 2788 30648 2840 30704
rect 2840 30648 2842 30704
rect 2786 30506 2788 30562
rect 2788 30506 2840 30562
rect 2840 30506 2842 30562
rect 175 28511 231 28567
rect 317 28511 373 28567
rect 175 28369 231 28425
rect 317 28369 373 28425
rect 1995 30107 2051 30109
rect 2137 30107 2193 30109
rect 2279 30107 2335 30109
rect 2421 30107 2477 30109
rect 2563 30107 2619 30109
rect 2705 30107 2761 30109
rect 2847 30107 2903 30109
rect 2989 30107 3045 30109
rect 3131 30107 3187 30109
rect 3273 30107 3329 30109
rect 1995 30055 2012 30107
rect 2012 30055 2051 30107
rect 2137 30055 2193 30107
rect 2279 30055 2335 30107
rect 2421 30055 2477 30107
rect 2563 30055 2619 30107
rect 2705 30055 2761 30107
rect 2847 30055 2903 30107
rect 2989 30055 3045 30107
rect 3131 30055 3187 30107
rect 3273 30055 3312 30107
rect 3312 30055 3329 30107
rect 1995 30053 2051 30055
rect 2137 30053 2193 30055
rect 2279 30053 2335 30055
rect 2421 30053 2477 30055
rect 2563 30053 2619 30055
rect 2705 30053 2761 30055
rect 2847 30053 2903 30055
rect 2989 30053 3045 30055
rect 3131 30053 3187 30055
rect 3273 30053 3329 30055
rect 7022 30790 7024 30846
rect 7024 30790 7076 30846
rect 7076 30790 7078 30846
rect 7022 30648 7024 30704
rect 7024 30648 7076 30704
rect 7076 30648 7078 30704
rect 7022 30506 7024 30562
rect 7024 30506 7076 30562
rect 7076 30506 7078 30562
rect 175 28227 231 28283
rect 317 28227 373 28283
rect 175 28085 231 28141
rect 317 28085 373 28141
rect 7997 40314 8053 40316
rect 8139 40314 8195 40316
rect 8281 40314 8337 40316
rect 8423 40314 8479 40316
rect 8565 40314 8621 40316
rect 8707 40314 8763 40316
rect 8849 40314 8905 40316
rect 8991 40314 9047 40316
rect 9133 40314 9189 40316
rect 9275 40314 9331 40316
rect 9417 40314 9473 40316
rect 9559 40314 9615 40316
rect 9701 40314 9757 40316
rect 7997 40262 8053 40314
rect 8139 40262 8195 40314
rect 8281 40262 8337 40314
rect 8423 40262 8479 40314
rect 8565 40262 8621 40314
rect 8707 40262 8763 40314
rect 8849 40262 8905 40314
rect 8991 40262 9047 40314
rect 9133 40262 9189 40314
rect 9275 40262 9331 40314
rect 9417 40262 9473 40314
rect 9559 40262 9615 40314
rect 9701 40262 9720 40314
rect 9720 40262 9757 40314
rect 7997 40260 8053 40262
rect 8139 40260 8195 40262
rect 8281 40260 8337 40262
rect 8423 40260 8479 40262
rect 8565 40260 8621 40262
rect 8707 40260 8763 40262
rect 8849 40260 8905 40262
rect 8991 40260 9047 40262
rect 9133 40260 9189 40262
rect 9275 40260 9331 40262
rect 9417 40260 9473 40262
rect 9559 40260 9615 40262
rect 9701 40260 9757 40262
rect 10337 39704 10339 39760
rect 10339 39704 10391 39760
rect 10391 39704 10393 39760
rect 10337 39562 10339 39618
rect 10339 39562 10391 39618
rect 10391 39562 10393 39618
rect 10337 39420 10339 39476
rect 10339 39420 10391 39476
rect 10391 39420 10393 39476
rect 10337 39278 10339 39334
rect 10339 39278 10391 39334
rect 10391 39278 10393 39334
rect 10337 39136 10339 39192
rect 10339 39136 10391 39192
rect 10391 39136 10393 39192
rect 10337 38994 10339 39050
rect 10339 38994 10391 39050
rect 10391 38994 10393 39050
rect 10337 38852 10339 38908
rect 10339 38852 10391 38908
rect 10391 38852 10393 38908
rect 11210 39704 11212 39760
rect 11212 39704 11264 39760
rect 11264 39704 11266 39760
rect 11210 39562 11212 39618
rect 11212 39562 11264 39618
rect 11264 39562 11266 39618
rect 11210 39420 11212 39476
rect 11212 39420 11264 39476
rect 11264 39420 11266 39476
rect 11210 39278 11212 39334
rect 11212 39278 11264 39334
rect 11264 39278 11266 39334
rect 11210 39136 11212 39192
rect 11212 39136 11264 39192
rect 11264 39136 11266 39192
rect 11210 38994 11212 39050
rect 11212 38994 11264 39050
rect 11264 38994 11266 39050
rect 10337 38710 10393 38766
rect 11210 38852 11212 38908
rect 11212 38852 11264 38908
rect 11264 38852 11266 38908
rect 11210 38710 11266 38766
rect 8681 35946 8737 35982
rect 8681 35926 8735 35946
rect 8735 35926 8737 35946
rect 8681 35784 8737 35840
rect 8681 35642 8737 35698
rect 8681 35500 8737 35556
rect 8681 35358 8737 35414
rect 8681 35216 8737 35272
rect 8681 35074 8737 35130
rect 8681 34932 8737 34988
rect 8681 34790 8737 34846
rect 8681 34648 8737 34704
rect 8681 34506 8737 34562
rect 13191 42912 13247 42968
rect 13303 42912 13359 42968
rect 13415 42912 13471 42968
rect 13191 42800 13247 42856
rect 13303 42800 13359 42856
rect 13415 42800 13471 42856
rect 13191 42688 13247 42744
rect 13303 42688 13359 42744
rect 13415 42688 13471 42744
rect 13191 42576 13247 42632
rect 13303 42576 13359 42632
rect 13415 42576 13471 42632
rect 13191 42464 13247 42520
rect 13303 42464 13359 42520
rect 13415 42464 13471 42520
rect 13191 42352 13247 42408
rect 13303 42352 13359 42408
rect 13415 42352 13471 42408
rect 13191 42240 13247 42296
rect 13303 42240 13359 42296
rect 13415 42240 13471 42296
rect 13191 42128 13247 42184
rect 13303 42128 13359 42184
rect 13415 42128 13471 42184
rect 13191 42016 13247 42072
rect 13303 42016 13359 42072
rect 13415 42016 13471 42072
rect 13191 41904 13247 41960
rect 13303 41904 13359 41960
rect 13415 41904 13471 41960
rect 13191 41792 13247 41848
rect 13303 41792 13359 41848
rect 13415 41792 13471 41848
rect 14410 55711 14466 55767
rect 14552 55711 14608 55767
rect 14694 55711 14750 55767
rect 14410 55569 14466 55625
rect 14552 55569 14608 55625
rect 14694 55569 14750 55625
rect 14410 55427 14466 55483
rect 14552 55427 14608 55483
rect 14694 55427 14750 55483
rect 14410 55285 14466 55341
rect 14552 55285 14608 55341
rect 14694 55285 14750 55341
rect 14410 55143 14466 55199
rect 14552 55143 14608 55199
rect 14694 55143 14750 55199
rect 14410 55001 14466 55057
rect 14552 55001 14608 55057
rect 14694 55001 14750 55057
rect 14410 54859 14466 54915
rect 14552 54859 14608 54915
rect 14694 54859 14750 54915
rect 14410 54717 14466 54773
rect 14552 54717 14608 54773
rect 14694 54717 14750 54773
rect 14410 54575 14466 54631
rect 14552 54575 14608 54631
rect 14694 54575 14750 54631
rect 14410 54433 14466 54489
rect 14552 54433 14608 54489
rect 14694 54433 14750 54489
rect 14952 52433 14954 52489
rect 14954 52433 15006 52489
rect 15006 52433 15008 52489
rect 14952 52291 14954 52347
rect 14954 52291 15006 52347
rect 15006 52291 15008 52347
rect 14952 52149 14954 52205
rect 14954 52149 15006 52205
rect 15006 52149 15008 52205
rect 14952 52007 14954 52063
rect 14954 52007 15006 52063
rect 15006 52007 15008 52063
rect 14952 51865 14954 51921
rect 14954 51865 15006 51921
rect 15006 51865 15008 51921
rect 14952 51723 14954 51779
rect 14954 51723 15006 51779
rect 15006 51723 15008 51779
rect 14952 51581 14954 51637
rect 14954 51581 15006 51637
rect 15006 51581 15008 51637
rect 14952 51439 14954 51495
rect 14954 51439 15006 51495
rect 15006 51439 15008 51495
rect 14952 51297 14954 51353
rect 14954 51297 15006 51353
rect 15006 51297 15008 51353
rect 14410 47704 14466 47760
rect 14552 47704 14608 47760
rect 14694 47704 14750 47760
rect 14410 47562 14466 47618
rect 14552 47562 14608 47618
rect 14694 47562 14750 47618
rect 14410 47420 14466 47476
rect 14552 47420 14608 47476
rect 14694 47420 14750 47476
rect 14410 47278 14466 47334
rect 14552 47278 14608 47334
rect 14694 47278 14750 47334
rect 14410 47136 14466 47192
rect 14552 47136 14608 47192
rect 14694 47136 14750 47192
rect 14410 46994 14466 47050
rect 14552 46994 14608 47050
rect 14694 46994 14750 47050
rect 14410 46852 14466 46908
rect 14552 46852 14608 46908
rect 14694 46852 14750 46908
rect 14410 46710 14466 46766
rect 14552 46710 14608 46766
rect 14694 46710 14750 46766
rect 14410 46568 14466 46624
rect 14552 46568 14608 46624
rect 14694 46568 14750 46624
rect 14410 46426 14466 46482
rect 14552 46426 14608 46482
rect 14694 46426 14750 46482
rect 14410 41304 14466 41360
rect 14552 41304 14608 41360
rect 14694 41304 14750 41360
rect 14410 41162 14466 41218
rect 14552 41162 14608 41218
rect 14694 41162 14750 41218
rect 14410 41020 14466 41076
rect 14552 41020 14608 41076
rect 14694 41020 14750 41076
rect 14410 40878 14466 40934
rect 14552 40878 14608 40934
rect 14694 40878 14750 40934
rect 14410 40736 14466 40792
rect 14552 40736 14608 40792
rect 14694 40736 14750 40792
rect 14410 40594 14466 40650
rect 14552 40594 14608 40650
rect 14694 40594 14750 40650
rect 14410 40452 14466 40508
rect 14552 40452 14608 40508
rect 14694 40452 14750 40508
rect 12758 40314 12814 40316
rect 12900 40314 12956 40316
rect 13042 40314 13098 40316
rect 13184 40314 13240 40316
rect 13326 40314 13382 40316
rect 13468 40314 13524 40316
rect 13610 40314 13666 40316
rect 13752 40314 13808 40316
rect 12758 40262 12784 40314
rect 12784 40262 12814 40314
rect 12900 40262 12956 40314
rect 13042 40262 13098 40314
rect 13184 40262 13240 40314
rect 13326 40262 13382 40314
rect 13468 40262 13524 40314
rect 13610 40262 13666 40314
rect 13752 40262 13772 40314
rect 13772 40262 13808 40314
rect 12758 40260 12814 40262
rect 12900 40260 12956 40262
rect 13042 40260 13098 40262
rect 13184 40260 13240 40262
rect 13326 40260 13382 40262
rect 13468 40260 13524 40262
rect 13610 40260 13666 40262
rect 13752 40260 13808 40262
rect 14410 40310 14466 40366
rect 14552 40310 14608 40366
rect 14694 40310 14750 40366
rect 14410 40168 14466 40224
rect 14552 40168 14608 40224
rect 14694 40168 14750 40224
rect 14410 40026 14466 40082
rect 14552 40026 14608 40082
rect 14694 40026 14750 40082
rect 12416 38104 12472 38160
rect 12558 38104 12614 38160
rect 12416 37962 12472 38018
rect 12558 37962 12614 38018
rect 12416 37820 12472 37876
rect 12558 37820 12614 37876
rect 10435 37568 10491 37570
rect 10577 37568 10633 37570
rect 10719 37568 10775 37570
rect 10861 37568 10917 37570
rect 11003 37568 11059 37570
rect 11145 37568 11201 37570
rect 11287 37568 11343 37570
rect 11429 37568 11485 37570
rect 10435 37516 10491 37568
rect 10577 37516 10633 37568
rect 10719 37516 10775 37568
rect 10861 37516 10917 37568
rect 11003 37516 11059 37568
rect 11145 37516 11201 37568
rect 11287 37516 11343 37568
rect 11429 37516 11485 37568
rect 10435 37514 10491 37516
rect 10577 37514 10633 37516
rect 10719 37514 10775 37516
rect 10861 37514 10917 37516
rect 11003 37514 11059 37516
rect 11145 37514 11201 37516
rect 11287 37514 11343 37516
rect 11429 37514 11485 37516
rect 11008 36030 11064 36086
rect 10110 35946 10166 35982
rect 10110 35926 10112 35946
rect 10112 35926 10164 35946
rect 10164 35926 10166 35946
rect 10110 35784 10112 35840
rect 10112 35784 10164 35840
rect 10164 35784 10166 35840
rect 10110 35642 10112 35698
rect 10112 35642 10164 35698
rect 10164 35642 10166 35698
rect 10110 35500 10112 35556
rect 10112 35500 10164 35556
rect 10164 35500 10166 35556
rect 10110 35358 10112 35414
rect 10112 35358 10164 35414
rect 10164 35358 10166 35414
rect 10110 35216 10112 35272
rect 10112 35216 10164 35272
rect 10164 35216 10166 35272
rect 10110 35074 10112 35130
rect 10112 35074 10164 35130
rect 10164 35074 10166 35130
rect 10110 34932 10112 34988
rect 10112 34932 10164 34988
rect 10164 34932 10166 34988
rect 10110 34790 10112 34846
rect 10112 34790 10164 34846
rect 10164 34790 10166 34846
rect 10110 34648 10112 34704
rect 10112 34648 10164 34704
rect 10164 34648 10166 34704
rect 10110 34542 10112 34562
rect 10112 34542 10164 34562
rect 10164 34542 10166 34562
rect 10110 34506 10166 34542
rect 11008 35888 11010 35944
rect 11010 35888 11062 35944
rect 11062 35888 11064 35944
rect 11008 35746 11010 35802
rect 11010 35746 11062 35802
rect 11062 35746 11064 35802
rect 11008 35604 11010 35660
rect 11010 35604 11062 35660
rect 11062 35604 11064 35660
rect 11008 35462 11010 35518
rect 11010 35462 11062 35518
rect 11062 35462 11064 35518
rect 11008 35320 11010 35376
rect 11010 35320 11062 35376
rect 11062 35320 11064 35376
rect 11008 35178 11010 35234
rect 11010 35178 11062 35234
rect 11062 35178 11064 35234
rect 11008 35036 11010 35092
rect 11010 35036 11062 35092
rect 11062 35036 11064 35092
rect 11008 34894 11010 34950
rect 11010 34894 11062 34950
rect 11062 34894 11064 34950
rect 11008 34752 11010 34808
rect 11010 34752 11062 34808
rect 11062 34752 11064 34808
rect 11008 34610 11010 34666
rect 11010 34610 11062 34666
rect 11062 34610 11064 34666
rect 11008 34468 11010 34524
rect 11010 34468 11062 34524
rect 11062 34468 11064 34524
rect 11008 34326 11010 34382
rect 11010 34326 11062 34382
rect 11062 34326 11064 34382
rect 12416 37678 12472 37734
rect 12558 37678 12614 37734
rect 12416 37536 12472 37592
rect 12558 37536 12614 37592
rect 12416 37394 12472 37450
rect 12558 37394 12614 37450
rect 12416 37252 12472 37308
rect 12558 37252 12614 37308
rect 12416 37110 12472 37166
rect 12558 37110 12614 37166
rect 12416 36968 12472 37024
rect 12558 36968 12614 37024
rect 12416 36826 12472 36882
rect 12558 36826 12614 36882
rect 11906 35946 11962 35982
rect 11906 35926 11908 35946
rect 11908 35926 11960 35946
rect 11960 35926 11962 35946
rect 11906 35784 11908 35840
rect 11908 35784 11960 35840
rect 11960 35784 11962 35840
rect 11906 35642 11908 35698
rect 11908 35642 11960 35698
rect 11960 35642 11962 35698
rect 11906 35500 11908 35556
rect 11908 35500 11960 35556
rect 11960 35500 11962 35556
rect 11906 35358 11908 35414
rect 11908 35358 11960 35414
rect 11960 35358 11962 35414
rect 11906 35216 11908 35272
rect 11908 35216 11960 35272
rect 11960 35216 11962 35272
rect 11906 35074 11908 35130
rect 11908 35074 11960 35130
rect 11960 35074 11962 35130
rect 11906 34932 11908 34988
rect 11908 34932 11960 34988
rect 11960 34932 11962 34988
rect 11906 34790 11908 34846
rect 11908 34790 11960 34846
rect 11960 34790 11962 34846
rect 11906 34648 11908 34704
rect 11908 34648 11960 34704
rect 11960 34648 11962 34704
rect 11906 34542 11908 34562
rect 11908 34542 11960 34562
rect 11960 34542 11962 34562
rect 11906 34506 11962 34542
rect 11008 34184 11010 34240
rect 11010 34184 11062 34240
rect 11062 34184 11064 34240
rect 11008 34042 11010 34098
rect 11010 34042 11062 34098
rect 11062 34042 11064 34098
rect 11008 33900 11010 33956
rect 11010 33900 11062 33956
rect 11062 33900 11064 33956
rect 11008 33758 11010 33814
rect 11010 33758 11062 33814
rect 11062 33758 11064 33814
rect 11008 33616 11010 33672
rect 11010 33616 11062 33672
rect 11062 33616 11064 33672
rect 11008 32849 11064 32905
rect 14952 38143 15008 38160
rect 14952 38104 14954 38143
rect 14954 38104 15006 38143
rect 15006 38104 15008 38143
rect 14952 37962 14954 38018
rect 14954 37962 15006 38018
rect 15006 37962 15008 38018
rect 14952 37820 14954 37876
rect 14954 37820 15006 37876
rect 15006 37820 15008 37876
rect 14952 37678 14954 37734
rect 14954 37678 15006 37734
rect 15006 37678 15008 37734
rect 14952 37536 14954 37592
rect 14954 37536 15006 37592
rect 15006 37536 15008 37592
rect 14952 37394 14954 37450
rect 14954 37394 15006 37450
rect 15006 37394 15008 37450
rect 14952 37252 14954 37308
rect 14954 37252 15006 37308
rect 15006 37252 15008 37308
rect 14952 37110 14954 37166
rect 14954 37110 15006 37166
rect 15006 37110 15008 37166
rect 14952 36968 14954 37024
rect 14954 36968 15006 37024
rect 15006 36968 15008 37024
rect 14952 36843 14954 36882
rect 14954 36843 15006 36882
rect 15006 36843 15008 36882
rect 14952 36826 15008 36843
rect 14410 33292 14466 33348
rect 14552 33292 14566 33348
rect 14566 33292 14608 33348
rect 14694 33292 14750 33348
rect 14410 33150 14466 33206
rect 14552 33150 14566 33206
rect 14566 33150 14608 33206
rect 14694 33150 14750 33206
rect 14410 33008 14466 33064
rect 14552 33008 14566 33064
rect 14566 33008 14608 33064
rect 14694 33008 14750 33064
rect 11008 32707 11010 32763
rect 11010 32707 11062 32763
rect 11062 32707 11064 32763
rect 7986 32690 8042 32692
rect 7986 32636 7988 32690
rect 7988 32636 8040 32690
rect 8040 32636 8042 32690
rect 7986 32494 7988 32550
rect 7988 32494 8040 32550
rect 8040 32494 8042 32550
rect 7986 32352 7988 32408
rect 7988 32352 8040 32408
rect 8040 32352 8042 32408
rect 7986 32210 7988 32266
rect 7988 32210 8040 32266
rect 8040 32210 8042 32266
rect 7986 32068 7988 32124
rect 7988 32068 8040 32124
rect 8040 32068 8042 32124
rect 7986 31926 7988 31982
rect 7988 31926 8040 31982
rect 8040 31926 8042 31982
rect 7986 31784 7988 31840
rect 7988 31784 8040 31840
rect 8040 31784 8042 31840
rect 7986 31642 7988 31698
rect 7988 31642 8040 31698
rect 8040 31642 8042 31698
rect 7986 31500 7988 31556
rect 7988 31500 8040 31556
rect 8040 31500 8042 31556
rect 7986 31358 7988 31414
rect 7988 31358 8040 31414
rect 8040 31358 8042 31414
rect 7986 31216 7988 31272
rect 7988 31216 8040 31272
rect 8040 31216 8042 31272
rect 7986 31074 7988 31130
rect 7988 31074 8040 31130
rect 8040 31074 8042 31130
rect 9378 32690 9434 32693
rect 9378 32637 9380 32690
rect 9380 32637 9432 32690
rect 9432 32637 9434 32690
rect 9378 32495 9380 32551
rect 9380 32495 9432 32551
rect 9432 32495 9434 32551
rect 9378 32353 9380 32409
rect 9380 32353 9432 32409
rect 9432 32353 9434 32409
rect 9378 32211 9380 32267
rect 9380 32211 9432 32267
rect 9432 32211 9434 32267
rect 9378 32069 9380 32125
rect 9380 32069 9432 32125
rect 9432 32069 9434 32125
rect 9378 31927 9380 31983
rect 9380 31927 9432 31983
rect 9432 31927 9434 31983
rect 9378 31785 9380 31841
rect 9380 31785 9432 31841
rect 9432 31785 9434 31841
rect 9378 31643 9380 31699
rect 9380 31643 9432 31699
rect 9432 31643 9434 31699
rect 9378 31501 9380 31557
rect 9380 31501 9432 31557
rect 9432 31501 9434 31557
rect 9378 31359 9380 31415
rect 9380 31359 9432 31415
rect 9432 31359 9434 31415
rect 9378 31217 9380 31273
rect 9380 31217 9432 31273
rect 9432 31217 9434 31273
rect 9378 31078 9380 31131
rect 9380 31078 9432 31131
rect 9432 31078 9434 31131
rect 9378 31075 9434 31078
rect 9794 32690 9850 32693
rect 9794 32637 9796 32690
rect 9796 32637 9848 32690
rect 9848 32637 9850 32690
rect 9794 32495 9796 32551
rect 9796 32495 9848 32551
rect 9848 32495 9850 32551
rect 9794 32353 9796 32409
rect 9796 32353 9848 32409
rect 9848 32353 9850 32409
rect 9794 32211 9796 32267
rect 9796 32211 9848 32267
rect 9848 32211 9850 32267
rect 9794 32069 9796 32125
rect 9796 32069 9848 32125
rect 9848 32069 9850 32125
rect 9794 31927 9796 31983
rect 9796 31927 9848 31983
rect 9848 31927 9850 31983
rect 9794 31785 9796 31841
rect 9796 31785 9848 31841
rect 9848 31785 9850 31841
rect 9794 31643 9796 31699
rect 9796 31643 9848 31699
rect 9848 31643 9850 31699
rect 9794 31501 9796 31557
rect 9796 31501 9848 31557
rect 9848 31501 9850 31557
rect 9794 31359 9796 31415
rect 9796 31359 9848 31415
rect 9848 31359 9850 31415
rect 9794 31217 9796 31273
rect 9796 31217 9848 31273
rect 9848 31217 9850 31273
rect 9794 31078 9796 31131
rect 9796 31078 9848 31131
rect 9848 31078 9850 31131
rect 9794 31075 9850 31078
rect 10282 32690 10338 32693
rect 10282 32637 10284 32690
rect 10284 32637 10336 32690
rect 10336 32637 10338 32690
rect 10282 32495 10284 32551
rect 10284 32495 10336 32551
rect 10336 32495 10338 32551
rect 10282 32353 10284 32409
rect 10284 32353 10336 32409
rect 10336 32353 10338 32409
rect 10282 32211 10284 32267
rect 10284 32211 10336 32267
rect 10336 32211 10338 32267
rect 10282 32069 10284 32125
rect 10284 32069 10336 32125
rect 10336 32069 10338 32125
rect 10282 31927 10284 31983
rect 10284 31927 10336 31983
rect 10336 31927 10338 31983
rect 10282 31785 10284 31841
rect 10284 31785 10336 31841
rect 10336 31785 10338 31841
rect 10282 31643 10284 31699
rect 10284 31643 10336 31699
rect 10336 31643 10338 31699
rect 10282 31501 10284 31557
rect 10284 31501 10336 31557
rect 10336 31501 10338 31557
rect 10282 31359 10284 31415
rect 10284 31359 10336 31415
rect 10336 31359 10338 31415
rect 10282 31217 10284 31273
rect 10284 31217 10336 31273
rect 10336 31217 10338 31273
rect 10282 31078 10284 31131
rect 10284 31078 10336 31131
rect 10336 31078 10338 31131
rect 10282 31075 10338 31078
rect 10770 32640 10826 32642
rect 10770 32586 10772 32640
rect 10772 32586 10824 32640
rect 10824 32586 10826 32640
rect 10770 32444 10772 32500
rect 10772 32444 10824 32500
rect 10824 32444 10826 32500
rect 10770 32302 10772 32358
rect 10772 32302 10824 32358
rect 10824 32302 10826 32358
rect 10770 32160 10772 32216
rect 10772 32160 10824 32216
rect 10824 32160 10826 32216
rect 10770 32018 10772 32074
rect 10772 32018 10824 32074
rect 10824 32018 10826 32074
rect 10770 31876 10772 31932
rect 10772 31876 10824 31932
rect 10824 31876 10826 31932
rect 10770 31734 10772 31790
rect 10772 31734 10824 31790
rect 10824 31734 10826 31790
rect 10770 31592 10772 31648
rect 10772 31592 10824 31648
rect 10824 31592 10826 31648
rect 10770 31450 10772 31506
rect 10772 31450 10824 31506
rect 10824 31450 10826 31506
rect 10770 31308 10772 31364
rect 10772 31308 10824 31364
rect 10824 31308 10826 31364
rect 10770 31166 10772 31222
rect 10772 31166 10824 31222
rect 10824 31166 10826 31222
rect 10770 31028 10772 31080
rect 10772 31028 10824 31080
rect 10824 31028 10826 31080
rect 10770 31024 10826 31028
rect 14410 32866 14466 32922
rect 14552 32866 14566 32922
rect 14566 32866 14608 32922
rect 14694 32866 14750 32922
rect 14410 32724 14466 32780
rect 14552 32724 14566 32780
rect 14566 32724 14608 32780
rect 14694 32724 14750 32780
rect 11008 32565 11010 32621
rect 11010 32565 11062 32621
rect 11062 32565 11064 32621
rect 11008 32423 11010 32479
rect 11010 32423 11062 32479
rect 11062 32423 11064 32479
rect 11008 32281 11010 32337
rect 11010 32281 11062 32337
rect 11062 32281 11064 32337
rect 11008 32139 11010 32195
rect 11010 32139 11062 32195
rect 11062 32139 11064 32195
rect 11008 31997 11010 32053
rect 11010 31997 11062 32053
rect 11062 31997 11064 32053
rect 11008 31855 11010 31911
rect 11010 31855 11062 31911
rect 11062 31855 11064 31911
rect 11008 31713 11010 31769
rect 11010 31713 11062 31769
rect 11062 31713 11064 31769
rect 11008 31571 11010 31627
rect 11010 31571 11062 31627
rect 11062 31571 11064 31627
rect 11008 31429 11010 31485
rect 11010 31429 11062 31485
rect 11062 31429 11064 31485
rect 11008 31287 11010 31343
rect 11010 31287 11062 31343
rect 11062 31287 11064 31343
rect 11008 31145 11010 31201
rect 11010 31145 11062 31201
rect 11062 31145 11064 31201
rect 11008 31005 11010 31059
rect 11010 31005 11062 31059
rect 11062 31005 11064 31059
rect 11008 31003 11064 31005
rect 11246 32640 11302 32642
rect 11246 32586 11248 32640
rect 11248 32586 11300 32640
rect 11300 32586 11302 32640
rect 11246 32444 11248 32500
rect 11248 32444 11300 32500
rect 11300 32444 11302 32500
rect 11246 32302 11248 32358
rect 11248 32302 11300 32358
rect 11300 32302 11302 32358
rect 11246 32160 11248 32216
rect 11248 32160 11300 32216
rect 11300 32160 11302 32216
rect 11246 32018 11248 32074
rect 11248 32018 11300 32074
rect 11300 32018 11302 32074
rect 11246 31876 11248 31932
rect 11248 31876 11300 31932
rect 11300 31876 11302 31932
rect 11246 31734 11248 31790
rect 11248 31734 11300 31790
rect 11300 31734 11302 31790
rect 11246 31592 11248 31648
rect 11248 31592 11300 31648
rect 11300 31592 11302 31648
rect 11246 31450 11248 31506
rect 11248 31450 11300 31506
rect 11300 31450 11302 31506
rect 11246 31308 11248 31364
rect 11248 31308 11300 31364
rect 11300 31308 11302 31364
rect 11246 31166 11248 31222
rect 11248 31166 11300 31222
rect 11300 31166 11302 31222
rect 11246 31028 11248 31080
rect 11248 31028 11300 31080
rect 11300 31028 11302 31080
rect 11246 31024 11302 31028
rect 11734 32690 11790 32693
rect 11734 32637 11736 32690
rect 11736 32637 11788 32690
rect 11788 32637 11790 32690
rect 11734 32495 11736 32551
rect 11736 32495 11788 32551
rect 11788 32495 11790 32551
rect 11734 32353 11736 32409
rect 11736 32353 11788 32409
rect 11788 32353 11790 32409
rect 11734 32211 11736 32267
rect 11736 32211 11788 32267
rect 11788 32211 11790 32267
rect 11734 32069 11736 32125
rect 11736 32069 11788 32125
rect 11788 32069 11790 32125
rect 11734 31927 11736 31983
rect 11736 31927 11788 31983
rect 11788 31927 11790 31983
rect 11734 31785 11736 31841
rect 11736 31785 11788 31841
rect 11788 31785 11790 31841
rect 11734 31643 11736 31699
rect 11736 31643 11788 31699
rect 11788 31643 11790 31699
rect 11734 31501 11736 31557
rect 11736 31501 11788 31557
rect 11788 31501 11790 31557
rect 11734 31359 11736 31415
rect 11736 31359 11788 31415
rect 11788 31359 11790 31415
rect 11734 31217 11736 31273
rect 11736 31217 11788 31273
rect 11788 31217 11790 31273
rect 11734 31078 11736 31131
rect 11736 31078 11788 31131
rect 11788 31078 11790 31131
rect 11734 31075 11790 31078
rect 12222 32690 12278 32692
rect 12222 32636 12224 32690
rect 12224 32636 12276 32690
rect 12276 32636 12278 32690
rect 12222 32494 12224 32550
rect 12224 32494 12276 32550
rect 12276 32494 12278 32550
rect 12222 32352 12224 32408
rect 12224 32352 12276 32408
rect 12276 32352 12278 32408
rect 12222 32210 12224 32266
rect 12224 32210 12276 32266
rect 12276 32210 12278 32266
rect 12222 32068 12224 32124
rect 12224 32068 12276 32124
rect 12276 32068 12278 32124
rect 12222 31926 12224 31982
rect 12224 31926 12276 31982
rect 12276 31926 12278 31982
rect 12222 31784 12224 31840
rect 12224 31784 12276 31840
rect 12276 31784 12278 31840
rect 12222 31642 12224 31698
rect 12224 31642 12276 31698
rect 12276 31642 12278 31698
rect 12222 31500 12224 31556
rect 12224 31500 12276 31556
rect 12276 31500 12278 31556
rect 12222 31358 12224 31414
rect 12224 31358 12276 31414
rect 12276 31358 12278 31414
rect 12222 31216 12224 31272
rect 12224 31216 12276 31272
rect 12276 31216 12278 31272
rect 12222 31074 12224 31130
rect 12224 31074 12276 31130
rect 12276 31074 12278 31130
rect 7986 30932 7988 30988
rect 7988 30932 8040 30988
rect 8040 30932 8042 30988
rect 12222 30932 12224 30988
rect 12224 30932 12276 30988
rect 12276 30932 12278 30988
rect 7986 30790 7988 30846
rect 7988 30790 8040 30846
rect 8040 30790 8042 30846
rect 7986 30648 7988 30704
rect 7988 30648 8040 30704
rect 8040 30648 8042 30704
rect 7986 30506 7988 30562
rect 7988 30506 8040 30562
rect 8040 30506 8042 30562
rect 12222 30790 12224 30846
rect 12224 30790 12276 30846
rect 12276 30790 12278 30846
rect 12222 30648 12224 30704
rect 12224 30648 12276 30704
rect 12276 30648 12278 30704
rect 12222 30506 12224 30562
rect 12224 30506 12276 30562
rect 12276 30506 12278 30562
rect 12638 32690 12694 32692
rect 12638 32636 12640 32690
rect 12640 32636 12692 32690
rect 12692 32636 12694 32690
rect 12638 32494 12640 32550
rect 12640 32494 12692 32550
rect 12692 32494 12694 32550
rect 12638 32352 12640 32408
rect 12640 32352 12692 32408
rect 12692 32352 12694 32408
rect 12638 32210 12640 32266
rect 12640 32210 12692 32266
rect 12692 32210 12694 32266
rect 12638 32068 12640 32124
rect 12640 32068 12692 32124
rect 12692 32068 12694 32124
rect 12638 31926 12640 31982
rect 12640 31926 12692 31982
rect 12692 31926 12694 31982
rect 12638 31784 12640 31840
rect 12640 31784 12692 31840
rect 12692 31784 12694 31840
rect 12638 31642 12640 31698
rect 12640 31642 12692 31698
rect 12692 31642 12694 31698
rect 12638 31500 12640 31556
rect 12640 31500 12692 31556
rect 12692 31500 12694 31556
rect 12638 31358 12640 31414
rect 12640 31358 12692 31414
rect 12692 31358 12694 31414
rect 12638 31216 12640 31272
rect 12640 31216 12692 31272
rect 12692 31216 12694 31272
rect 12638 31074 12640 31130
rect 12640 31074 12692 31130
rect 12692 31074 12694 31130
rect 12638 30932 12640 30988
rect 12640 30932 12692 30988
rect 12692 30932 12694 30988
rect 12638 30790 12640 30846
rect 12640 30790 12692 30846
rect 12692 30790 12694 30846
rect 12638 30648 12640 30704
rect 12640 30648 12692 30704
rect 12692 30648 12694 30704
rect 14030 32690 14086 32692
rect 14030 32636 14032 32690
rect 14032 32636 14084 32690
rect 14084 32636 14086 32690
rect 14030 32494 14032 32550
rect 14032 32494 14084 32550
rect 14084 32494 14086 32550
rect 14030 32352 14032 32408
rect 14032 32352 14084 32408
rect 14084 32352 14086 32408
rect 14030 32210 14032 32266
rect 14032 32210 14084 32266
rect 14084 32210 14086 32266
rect 14030 32068 14032 32124
rect 14032 32068 14084 32124
rect 14084 32068 14086 32124
rect 14030 31926 14032 31982
rect 14032 31926 14084 31982
rect 14084 31926 14086 31982
rect 14030 31784 14032 31840
rect 14032 31784 14084 31840
rect 14084 31784 14086 31840
rect 14030 31642 14032 31698
rect 14032 31642 14084 31698
rect 14084 31642 14086 31698
rect 14030 31500 14032 31556
rect 14032 31500 14084 31556
rect 14084 31500 14086 31556
rect 14030 31358 14032 31414
rect 14032 31358 14084 31414
rect 14084 31358 14086 31414
rect 14030 31216 14032 31272
rect 14032 31216 14084 31272
rect 14084 31216 14086 31272
rect 14030 31074 14032 31130
rect 14032 31074 14084 31130
rect 14084 31074 14086 31130
rect 14030 30932 14032 30988
rect 14032 30932 14084 30988
rect 14084 30932 14086 30988
rect 14030 30790 14032 30846
rect 14032 30790 14084 30846
rect 14084 30790 14086 30846
rect 12638 30506 12640 30562
rect 12640 30506 12692 30562
rect 12692 30506 12694 30562
rect 11932 30107 11988 30109
rect 12074 30107 12130 30109
rect 12216 30107 12272 30109
rect 12358 30107 12414 30109
rect 12500 30107 12556 30109
rect 12642 30107 12698 30109
rect 12784 30107 12840 30109
rect 12926 30107 12982 30109
rect 13068 30107 13124 30109
rect 13210 30107 13266 30109
rect 11932 30055 11949 30107
rect 11949 30055 11988 30107
rect 12074 30055 12130 30107
rect 12216 30055 12272 30107
rect 12358 30055 12414 30107
rect 12500 30055 12556 30107
rect 12642 30055 12698 30107
rect 12784 30055 12840 30107
rect 12926 30055 12982 30107
rect 13068 30055 13124 30107
rect 13210 30055 13249 30107
rect 13249 30055 13266 30107
rect 11932 30053 11988 30055
rect 12074 30053 12130 30055
rect 12216 30053 12272 30055
rect 12358 30053 12414 30055
rect 12500 30053 12556 30055
rect 12642 30053 12698 30055
rect 12784 30053 12840 30055
rect 12926 30053 12982 30055
rect 13068 30053 13124 30055
rect 13210 30053 13266 30055
rect 14030 30648 14032 30704
rect 14032 30648 14084 30704
rect 14084 30648 14086 30704
rect 14030 30506 14032 30562
rect 14032 30506 14084 30562
rect 14084 30506 14086 30562
rect 14410 32582 14466 32638
rect 14552 32582 14566 32638
rect 14566 32582 14608 32638
rect 14694 32582 14750 32638
rect 14410 32440 14466 32496
rect 14552 32440 14566 32496
rect 14566 32440 14608 32496
rect 14694 32440 14750 32496
rect 14410 32298 14466 32354
rect 14552 32298 14566 32354
rect 14566 32298 14608 32354
rect 14694 32298 14750 32354
rect 14410 32156 14466 32212
rect 14552 32156 14566 32212
rect 14566 32156 14608 32212
rect 14694 32156 14750 32212
rect 14410 32014 14466 32070
rect 14552 32014 14566 32070
rect 14566 32014 14608 32070
rect 14694 32014 14750 32070
rect 14410 31872 14466 31928
rect 14552 31872 14566 31928
rect 14566 31872 14608 31928
rect 14694 31872 14750 31928
rect 14410 31730 14466 31786
rect 14552 31730 14566 31786
rect 14566 31730 14608 31786
rect 14694 31730 14750 31786
rect 14410 31588 14466 31644
rect 14552 31588 14566 31644
rect 14566 31588 14608 31644
rect 14694 31588 14750 31644
rect 14410 31446 14466 31502
rect 14552 31446 14566 31502
rect 14566 31446 14608 31502
rect 14694 31446 14750 31502
rect 14410 31304 14466 31360
rect 14552 31304 14566 31360
rect 14566 31304 14608 31360
rect 14694 31304 14750 31360
rect 14410 31162 14466 31218
rect 14552 31162 14566 31218
rect 14566 31162 14608 31218
rect 14694 31162 14750 31218
rect 14410 31020 14466 31076
rect 14552 31020 14566 31076
rect 14566 31020 14608 31076
rect 14694 31020 14750 31076
rect 14410 30878 14466 30934
rect 14552 30878 14566 30934
rect 14566 30878 14608 30934
rect 14694 30878 14750 30934
rect 14410 30736 14466 30792
rect 14552 30736 14566 30792
rect 14566 30736 14608 30792
rect 14694 30736 14750 30792
rect 14410 30594 14466 30650
rect 14552 30594 14566 30650
rect 14566 30594 14608 30650
rect 14694 30594 14750 30650
rect 14410 30452 14466 30508
rect 14552 30452 14566 30508
rect 14566 30452 14608 30508
rect 14694 30452 14750 30508
rect 14410 30111 14466 30167
rect 14552 30111 14566 30167
rect 14566 30111 14608 30167
rect 14694 30111 14750 30167
rect 14410 29969 14466 30025
rect 14552 29969 14608 30025
rect 14694 29969 14750 30025
rect 14410 29827 14466 29883
rect 14552 29827 14608 29883
rect 14694 29827 14750 29883
rect 14410 29685 14466 29741
rect 14552 29685 14608 29741
rect 14694 29685 14750 29741
rect 14410 29543 14466 29599
rect 14552 29543 14608 29599
rect 14694 29543 14750 29599
rect 14410 29401 14466 29457
rect 14552 29401 14608 29457
rect 14694 29401 14750 29457
rect 14410 29259 14466 29315
rect 14552 29259 14608 29315
rect 14694 29259 14750 29315
rect 14410 29117 14466 29173
rect 14552 29117 14608 29173
rect 14694 29117 14750 29173
rect 14410 28975 14466 29031
rect 14552 28975 14608 29031
rect 14694 28975 14750 29031
rect 14410 28833 14466 28889
rect 14552 28833 14608 28889
rect 14694 28833 14750 28889
rect 175 27943 231 27999
rect 317 27943 373 27999
rect 175 27801 231 27857
rect 317 27801 373 27857
rect 175 27659 231 27715
rect 317 27659 373 27715
rect 175 27517 231 27573
rect 317 27517 373 27573
rect 175 27375 231 27431
rect 317 27375 373 27431
rect 175 27233 231 27289
rect 317 27233 373 27289
rect 14410 26892 14466 26948
rect 14552 26892 14608 26948
rect 14694 26892 14750 26948
rect 14410 26750 14466 26806
rect 14552 26750 14608 26806
rect 14694 26750 14750 26806
rect 14410 26608 14466 26664
rect 14552 26608 14608 26664
rect 14694 26608 14750 26664
rect 14410 26466 14466 26522
rect 14552 26466 14608 26522
rect 14694 26466 14750 26522
rect 14410 26324 14466 26380
rect 14552 26324 14608 26380
rect 14694 26324 14750 26380
rect 14410 26182 14466 26238
rect 14552 26182 14608 26238
rect 14694 26182 14750 26238
rect 14410 26040 14466 26096
rect 14552 26040 14608 26096
rect 14694 26040 14750 26096
rect 14410 25898 14466 25954
rect 14552 25898 14608 25954
rect 14694 25898 14750 25954
rect 14410 25756 14466 25812
rect 14552 25756 14608 25812
rect 14694 25756 14750 25812
rect 14410 25614 14466 25670
rect 14552 25614 14608 25670
rect 14694 25614 14750 25670
rect 14410 25472 14466 25528
rect 14552 25472 14608 25528
rect 14694 25472 14750 25528
rect 14410 25330 14466 25386
rect 14552 25330 14608 25386
rect 14694 25330 14750 25386
rect 14410 25188 14466 25244
rect 14552 25188 14608 25244
rect 14694 25188 14750 25244
rect 14410 25046 14466 25102
rect 14552 25046 14608 25102
rect 14694 25046 14750 25102
rect 14410 24904 14466 24960
rect 14552 24904 14608 24960
rect 14694 24904 14750 24960
rect 14410 24762 14466 24818
rect 14552 24762 14608 24818
rect 14694 24762 14750 24818
rect 14410 24620 14466 24676
rect 14552 24620 14608 24676
rect 14694 24620 14750 24676
rect 14410 24478 14466 24534
rect 14552 24478 14608 24534
rect 14694 24478 14750 24534
rect 14410 24336 14466 24392
rect 14552 24336 14608 24392
rect 14694 24336 14750 24392
rect 14410 24194 14466 24250
rect 14552 24194 14608 24250
rect 14694 24194 14750 24250
rect 14410 24052 14466 24108
rect 14552 24052 14608 24108
rect 14694 24052 14750 24108
rect 14410 23692 14466 23748
rect 14552 23692 14608 23748
rect 14694 23692 14750 23748
rect 14410 23550 14466 23606
rect 14552 23550 14608 23606
rect 14694 23550 14750 23606
rect 14410 23408 14466 23464
rect 14552 23408 14608 23464
rect 14694 23408 14750 23464
rect 14410 23266 14466 23322
rect 14552 23266 14608 23322
rect 14694 23266 14750 23322
rect 14410 23124 14466 23180
rect 14552 23124 14608 23180
rect 14694 23124 14750 23180
rect 14410 22982 14466 23038
rect 14552 22982 14608 23038
rect 14694 22982 14750 23038
rect 14410 22840 14466 22896
rect 14552 22840 14608 22896
rect 14694 22840 14750 22896
rect 14410 22698 14466 22754
rect 14552 22698 14608 22754
rect 14694 22698 14750 22754
rect 14410 22556 14466 22612
rect 14552 22556 14608 22612
rect 14694 22556 14750 22612
rect 14410 22414 14466 22470
rect 14552 22414 14608 22470
rect 14694 22414 14750 22470
rect 14410 22272 14466 22328
rect 14552 22272 14608 22328
rect 14694 22272 14750 22328
rect 14410 22130 14466 22186
rect 14552 22130 14608 22186
rect 14694 22130 14750 22186
rect 14410 21988 14466 22044
rect 14552 21988 14608 22044
rect 14694 21988 14750 22044
rect 14410 21846 14466 21902
rect 14552 21846 14608 21902
rect 14694 21846 14750 21902
rect 14410 21704 14466 21760
rect 14552 21704 14608 21760
rect 14694 21704 14750 21760
rect 14410 21562 14466 21618
rect 14552 21562 14608 21618
rect 14694 21562 14750 21618
rect 14410 21420 14466 21476
rect 14552 21420 14608 21476
rect 14694 21420 14750 21476
rect 14410 21278 14466 21334
rect 14552 21278 14608 21334
rect 14694 21278 14750 21334
rect 14410 21136 14466 21192
rect 14552 21136 14608 21192
rect 14694 21136 14750 21192
rect 14410 20994 14466 21050
rect 14552 20994 14608 21050
rect 14694 20994 14750 21050
rect 14410 20852 14466 20908
rect 14552 20852 14608 20908
rect 14694 20852 14750 20908
rect 14410 20492 14466 20548
rect 14552 20492 14608 20548
rect 14694 20492 14750 20548
rect 14410 20350 14466 20406
rect 14552 20350 14608 20406
rect 14694 20350 14750 20406
rect 14410 20208 14466 20264
rect 14552 20208 14608 20264
rect 14694 20208 14750 20264
rect 14410 20066 14466 20122
rect 14552 20066 14608 20122
rect 14694 20066 14750 20122
rect 14410 19924 14466 19980
rect 14552 19924 14608 19980
rect 14694 19924 14750 19980
rect 14410 19782 14466 19838
rect 14552 19782 14608 19838
rect 14694 19782 14750 19838
rect 14410 19640 14466 19696
rect 14552 19640 14608 19696
rect 14694 19640 14750 19696
rect 14410 19498 14466 19554
rect 14552 19498 14608 19554
rect 14694 19498 14750 19554
rect 14410 19356 14466 19412
rect 14552 19356 14608 19412
rect 14694 19356 14750 19412
rect 14410 19214 14466 19270
rect 14552 19214 14608 19270
rect 14694 19214 14750 19270
rect 14410 19072 14466 19128
rect 14552 19072 14608 19128
rect 14694 19072 14750 19128
rect 14410 18930 14466 18986
rect 14552 18930 14608 18986
rect 14694 18930 14750 18986
rect 14410 18788 14466 18844
rect 14552 18788 14608 18844
rect 14694 18788 14750 18844
rect 14410 18646 14466 18702
rect 14552 18646 14608 18702
rect 14694 18646 14750 18702
rect 14410 18504 14466 18560
rect 14552 18504 14608 18560
rect 14694 18504 14750 18560
rect 14410 18362 14466 18418
rect 14552 18362 14608 18418
rect 14694 18362 14750 18418
rect 14410 18220 14466 18276
rect 14552 18220 14608 18276
rect 14694 18220 14750 18276
rect 14410 18078 14466 18134
rect 14552 18078 14608 18134
rect 14694 18078 14750 18134
rect 14410 17936 14466 17992
rect 14552 17936 14608 17992
rect 14694 17936 14750 17992
rect 14410 17794 14466 17850
rect 14552 17794 14608 17850
rect 14694 17794 14750 17850
rect 14410 17652 14466 17708
rect 14552 17652 14608 17708
rect 14694 17652 14750 17708
rect 14410 17292 14466 17348
rect 14552 17292 14608 17348
rect 14694 17292 14750 17348
rect 14410 17150 14466 17206
rect 14552 17150 14608 17206
rect 14694 17150 14750 17206
rect 14410 17008 14466 17064
rect 14552 17008 14608 17064
rect 14694 17008 14750 17064
rect 14410 16866 14466 16922
rect 14552 16866 14608 16922
rect 14694 16866 14750 16922
rect 14410 16724 14466 16780
rect 14552 16724 14608 16780
rect 14694 16724 14750 16780
rect 14410 16582 14466 16638
rect 14552 16582 14608 16638
rect 14694 16582 14750 16638
rect 14410 16440 14466 16496
rect 14552 16440 14608 16496
rect 14694 16440 14750 16496
rect 14410 16298 14466 16354
rect 14552 16298 14608 16354
rect 14694 16298 14750 16354
rect 14410 16156 14466 16212
rect 14552 16156 14608 16212
rect 14694 16156 14750 16212
rect 14410 16014 14466 16070
rect 14552 16014 14608 16070
rect 14694 16014 14750 16070
rect 14410 15872 14466 15928
rect 14552 15872 14608 15928
rect 14694 15872 14750 15928
rect 14410 15730 14466 15786
rect 14552 15730 14608 15786
rect 14694 15730 14750 15786
rect 14410 15588 14466 15644
rect 14552 15588 14608 15644
rect 14694 15588 14750 15644
rect 14410 15446 14466 15502
rect 14552 15446 14608 15502
rect 14694 15446 14750 15502
rect 14410 15304 14466 15360
rect 14552 15304 14608 15360
rect 14694 15304 14750 15360
rect 14410 15162 14466 15218
rect 14552 15162 14608 15218
rect 14694 15162 14750 15218
rect 14410 15020 14466 15076
rect 14552 15020 14608 15076
rect 14694 15020 14750 15076
rect 14410 14878 14466 14934
rect 14552 14878 14608 14934
rect 14694 14878 14750 14934
rect 14410 14736 14466 14792
rect 14552 14736 14608 14792
rect 14694 14736 14750 14792
rect 14410 14594 14466 14650
rect 14552 14594 14608 14650
rect 14694 14594 14750 14650
rect 14410 14452 14466 14508
rect 14552 14452 14608 14508
rect 14694 14452 14750 14508
rect 175 10892 231 10948
rect 317 10892 373 10948
rect 175 10750 231 10806
rect 317 10750 373 10806
rect 175 10608 231 10664
rect 317 10608 373 10664
rect 175 10466 231 10522
rect 317 10466 373 10522
rect 175 10324 231 10380
rect 317 10324 373 10380
rect 175 10182 231 10238
rect 317 10182 373 10238
rect 175 10040 231 10096
rect 317 10040 373 10096
rect 175 9898 231 9954
rect 317 9898 373 9954
rect 175 9756 231 9812
rect 317 9756 373 9812
rect 175 9614 231 9670
rect 317 9614 373 9670
rect 175 9472 231 9528
rect 317 9472 373 9528
rect 175 9330 231 9386
rect 317 9330 373 9386
rect 175 9188 231 9244
rect 317 9188 373 9244
rect 175 9046 231 9102
rect 317 9046 373 9102
rect 175 8904 231 8960
rect 317 8904 373 8960
rect 175 8762 231 8818
rect 317 8762 373 8818
rect 175 8620 231 8676
rect 317 8620 373 8676
rect 175 8478 231 8534
rect 317 8478 373 8534
rect 175 8336 231 8392
rect 317 8336 373 8392
rect 175 8194 231 8250
rect 317 8194 373 8250
rect 175 8052 231 8108
rect 317 8052 373 8108
rect 175 7692 231 7748
rect 317 7692 373 7748
rect 175 7550 231 7606
rect 317 7550 373 7606
rect 175 7408 231 7464
rect 317 7408 373 7464
rect 175 7266 231 7322
rect 317 7266 373 7322
rect 175 7124 231 7180
rect 317 7124 373 7180
rect 175 6982 231 7038
rect 317 6982 373 7038
rect 175 6840 231 6896
rect 317 6840 373 6896
rect 175 6698 231 6754
rect 317 6698 373 6754
rect 175 6556 231 6612
rect 317 6556 373 6612
rect 175 6414 231 6470
rect 317 6414 373 6470
rect 175 6272 231 6328
rect 317 6272 373 6328
rect 175 6130 231 6186
rect 317 6130 373 6186
rect 175 5988 231 6044
rect 317 5988 373 6044
rect 175 5846 231 5902
rect 317 5846 373 5902
rect 175 5704 231 5760
rect 317 5704 373 5760
rect 175 5562 231 5618
rect 317 5562 373 5618
rect 175 5420 231 5476
rect 317 5420 373 5476
rect 175 5278 231 5334
rect 317 5278 373 5334
rect 175 5136 231 5192
rect 317 5136 373 5192
rect 175 4994 231 5050
rect 317 4994 373 5050
rect 175 4852 231 4908
rect 317 4852 373 4908
rect 175 4492 231 4548
rect 317 4492 373 4548
rect 175 4350 231 4406
rect 317 4350 373 4406
rect 175 4208 231 4264
rect 317 4208 373 4264
rect 175 4066 231 4122
rect 317 4066 373 4122
rect 175 3924 231 3980
rect 317 3924 373 3980
rect 175 3782 231 3838
rect 317 3782 373 3838
rect 175 3640 231 3696
rect 317 3640 373 3696
rect 175 3498 231 3554
rect 317 3498 373 3554
rect 175 3356 231 3412
rect 317 3356 373 3412
rect 175 3214 231 3270
rect 317 3214 373 3270
rect 175 3072 231 3128
rect 317 3072 373 3128
rect 175 2930 231 2986
rect 317 2930 373 2986
rect 175 2788 231 2844
rect 317 2788 373 2844
rect 175 2646 231 2702
rect 317 2646 373 2702
rect 175 2504 231 2560
rect 317 2504 373 2560
rect 175 2362 231 2418
rect 317 2362 373 2418
rect 175 2220 231 2276
rect 317 2220 373 2276
rect 175 2078 231 2134
rect 317 2078 373 2134
rect 175 1936 231 1992
rect 317 1936 373 1992
rect 175 1794 231 1850
rect 317 1794 373 1850
rect 175 1652 231 1708
rect 317 1652 373 1708
<< metal3 >>
rect 1886 57235 1962 57245
rect 1886 57179 1896 57235
rect 1952 57179 1962 57235
rect 1886 57093 1962 57179
rect 1886 57037 1896 57093
rect 1952 57037 1962 57093
rect 1886 56951 1962 57037
rect 1886 56895 1896 56951
rect 1952 56895 1962 56951
rect 1886 56809 1962 56895
rect 2490 57180 13642 57190
rect 2490 57124 2500 57180
rect 2556 57124 2642 57180
rect 2698 57124 2784 57180
rect 2840 57124 2926 57180
rect 2982 57124 3068 57180
rect 3124 57124 3210 57180
rect 3266 57124 3352 57180
rect 3408 57124 3494 57180
rect 3550 57124 3636 57180
rect 3692 57124 3778 57180
rect 3834 57124 3920 57180
rect 3976 57124 4062 57180
rect 4118 57124 4204 57180
rect 4260 57124 4346 57180
rect 4402 57124 4488 57180
rect 4544 57124 4630 57180
rect 4686 57124 4772 57180
rect 4828 57124 4914 57180
rect 4970 57124 5056 57180
rect 5112 57124 5198 57180
rect 5254 57124 5340 57180
rect 5396 57124 5482 57180
rect 5538 57124 5624 57180
rect 5680 57124 5766 57180
rect 5822 57124 5908 57180
rect 5964 57124 6050 57180
rect 6106 57124 6192 57180
rect 6248 57124 6334 57180
rect 6390 57124 6476 57180
rect 6532 57124 6618 57180
rect 6674 57124 6760 57180
rect 6816 57124 6902 57180
rect 6958 57124 7044 57180
rect 7100 57124 7186 57180
rect 7242 57124 7328 57180
rect 7384 57124 7470 57180
rect 7526 57124 7612 57180
rect 7668 57124 7754 57180
rect 7810 57124 7896 57180
rect 7952 57124 8038 57180
rect 8094 57124 8180 57180
rect 8236 57124 8322 57180
rect 8378 57124 8464 57180
rect 8520 57124 8606 57180
rect 8662 57124 8748 57180
rect 8804 57124 8890 57180
rect 8946 57124 9032 57180
rect 9088 57124 9174 57180
rect 9230 57124 9316 57180
rect 9372 57124 9458 57180
rect 9514 57124 9600 57180
rect 9656 57124 9742 57180
rect 9798 57124 9884 57180
rect 9940 57124 10026 57180
rect 10082 57124 10168 57180
rect 10224 57124 10310 57180
rect 10366 57124 10452 57180
rect 10508 57124 10594 57180
rect 10650 57124 10736 57180
rect 10792 57124 10878 57180
rect 10934 57124 11020 57180
rect 11076 57124 11162 57180
rect 11218 57124 11304 57180
rect 11360 57124 11446 57180
rect 11502 57124 11588 57180
rect 11644 57124 11730 57180
rect 11786 57124 11872 57180
rect 11928 57124 12014 57180
rect 12070 57124 12156 57180
rect 12212 57124 12298 57180
rect 12354 57124 12440 57180
rect 12496 57124 12582 57180
rect 12638 57124 12724 57180
rect 12780 57124 12866 57180
rect 12922 57124 13008 57180
rect 13064 57124 13150 57180
rect 13206 57124 13292 57180
rect 13348 57124 13434 57180
rect 13490 57124 13576 57180
rect 13632 57124 13642 57180
rect 2490 57038 13642 57124
rect 2490 56982 2500 57038
rect 2556 56982 2642 57038
rect 2698 56982 2784 57038
rect 2840 56982 2926 57038
rect 2982 56982 3068 57038
rect 3124 56982 3210 57038
rect 3266 56982 3352 57038
rect 3408 56982 3494 57038
rect 3550 56982 3636 57038
rect 3692 56982 3778 57038
rect 3834 56982 3920 57038
rect 3976 56982 4062 57038
rect 4118 56982 4204 57038
rect 4260 56982 4346 57038
rect 4402 56982 4488 57038
rect 4544 56982 4630 57038
rect 4686 56982 4772 57038
rect 4828 56982 4914 57038
rect 4970 56982 5056 57038
rect 5112 56982 5198 57038
rect 5254 56982 5340 57038
rect 5396 56982 5482 57038
rect 5538 56982 5624 57038
rect 5680 56982 5766 57038
rect 5822 56982 5908 57038
rect 5964 56982 6050 57038
rect 6106 56982 6192 57038
rect 6248 56982 6334 57038
rect 6390 56982 6476 57038
rect 6532 56982 6618 57038
rect 6674 56982 6760 57038
rect 6816 56982 6902 57038
rect 6958 56982 7044 57038
rect 7100 56982 7186 57038
rect 7242 56982 7328 57038
rect 7384 56982 7470 57038
rect 7526 56982 7612 57038
rect 7668 56982 7754 57038
rect 7810 56982 7896 57038
rect 7952 56982 8038 57038
rect 8094 56982 8180 57038
rect 8236 56982 8322 57038
rect 8378 56982 8464 57038
rect 8520 56982 8606 57038
rect 8662 56982 8748 57038
rect 8804 56982 8890 57038
rect 8946 56982 9032 57038
rect 9088 56982 9174 57038
rect 9230 56982 9316 57038
rect 9372 56982 9458 57038
rect 9514 56982 9600 57038
rect 9656 56982 9742 57038
rect 9798 56982 9884 57038
rect 9940 56982 10026 57038
rect 10082 56982 10168 57038
rect 10224 56982 10310 57038
rect 10366 56982 10452 57038
rect 10508 56982 10594 57038
rect 10650 56982 10736 57038
rect 10792 56982 10878 57038
rect 10934 56982 11020 57038
rect 11076 56982 11162 57038
rect 11218 56982 11304 57038
rect 11360 56982 11446 57038
rect 11502 56982 11588 57038
rect 11644 56982 11730 57038
rect 11786 56982 11872 57038
rect 11928 56982 12014 57038
rect 12070 56982 12156 57038
rect 12212 56982 12298 57038
rect 12354 56982 12440 57038
rect 12496 56982 12582 57038
rect 12638 56982 12724 57038
rect 12780 56982 12866 57038
rect 12922 56982 13008 57038
rect 13064 56982 13150 57038
rect 13206 56982 13292 57038
rect 13348 56982 13434 57038
rect 13490 56982 13576 57038
rect 13632 56982 13642 57038
rect 2490 56896 13642 56982
rect 2490 56840 2500 56896
rect 2556 56840 2642 56896
rect 2698 56840 2784 56896
rect 2840 56840 2926 56896
rect 2982 56840 3068 56896
rect 3124 56840 3210 56896
rect 3266 56840 3352 56896
rect 3408 56840 3494 56896
rect 3550 56840 3636 56896
rect 3692 56840 3778 56896
rect 3834 56840 3920 56896
rect 3976 56840 4062 56896
rect 4118 56840 4204 56896
rect 4260 56840 4346 56896
rect 4402 56840 4488 56896
rect 4544 56840 4630 56896
rect 4686 56840 4772 56896
rect 4828 56840 4914 56896
rect 4970 56840 5056 56896
rect 5112 56840 5198 56896
rect 5254 56840 5340 56896
rect 5396 56840 5482 56896
rect 5538 56840 5624 56896
rect 5680 56840 5766 56896
rect 5822 56840 5908 56896
rect 5964 56840 6050 56896
rect 6106 56840 6192 56896
rect 6248 56840 6334 56896
rect 6390 56840 6476 56896
rect 6532 56840 6618 56896
rect 6674 56840 6760 56896
rect 6816 56840 6902 56896
rect 6958 56840 7044 56896
rect 7100 56840 7186 56896
rect 7242 56840 7328 56896
rect 7384 56840 7470 56896
rect 7526 56840 7612 56896
rect 7668 56840 7754 56896
rect 7810 56840 7896 56896
rect 7952 56840 8038 56896
rect 8094 56840 8180 56896
rect 8236 56840 8322 56896
rect 8378 56840 8464 56896
rect 8520 56840 8606 56896
rect 8662 56840 8748 56896
rect 8804 56840 8890 56896
rect 8946 56840 9032 56896
rect 9088 56840 9174 56896
rect 9230 56840 9316 56896
rect 9372 56840 9458 56896
rect 9514 56840 9600 56896
rect 9656 56840 9742 56896
rect 9798 56840 9884 56896
rect 9940 56840 10026 56896
rect 10082 56840 10168 56896
rect 10224 56840 10310 56896
rect 10366 56840 10452 56896
rect 10508 56840 10594 56896
rect 10650 56840 10736 56896
rect 10792 56840 10878 56896
rect 10934 56840 11020 56896
rect 11076 56840 11162 56896
rect 11218 56840 11304 56896
rect 11360 56840 11446 56896
rect 11502 56840 11588 56896
rect 11644 56840 11730 56896
rect 11786 56840 11872 56896
rect 11928 56840 12014 56896
rect 12070 56840 12156 56896
rect 12212 56840 12298 56896
rect 12354 56840 12440 56896
rect 12496 56840 12582 56896
rect 12638 56840 12724 56896
rect 12780 56840 12866 56896
rect 12922 56840 13008 56896
rect 13064 56840 13150 56896
rect 13206 56840 13292 56896
rect 13348 56840 13434 56896
rect 13490 56840 13576 56896
rect 13632 56840 13642 56896
rect 2490 56830 13642 56840
rect 1886 56753 1896 56809
rect 1952 56753 1962 56809
rect 1886 56667 1962 56753
rect 1886 56611 1896 56667
rect 1952 56611 1962 56667
rect 1886 56525 1962 56611
rect 1886 56469 1896 56525
rect 1952 56469 1962 56525
rect 1886 56383 1962 56469
rect 1886 56327 1896 56383
rect 1952 56327 1962 56383
rect 1886 56241 1962 56327
rect 1886 56185 1896 56241
rect 1952 56185 1962 56241
rect 1886 56099 1962 56185
rect 1886 56043 1896 56099
rect 1952 56043 1962 56099
rect 2490 56438 13642 56448
rect 2490 56382 2500 56438
rect 2556 56382 2642 56438
rect 2698 56382 2784 56438
rect 2840 56382 2926 56438
rect 2982 56382 3068 56438
rect 3124 56382 3210 56438
rect 3266 56382 3352 56438
rect 3408 56382 3494 56438
rect 3550 56382 3636 56438
rect 3692 56382 3778 56438
rect 3834 56382 3920 56438
rect 3976 56382 4062 56438
rect 4118 56382 4204 56438
rect 4260 56382 4346 56438
rect 4402 56382 4488 56438
rect 4544 56382 4630 56438
rect 4686 56382 4772 56438
rect 4828 56382 4914 56438
rect 4970 56382 5056 56438
rect 5112 56382 5198 56438
rect 5254 56382 5340 56438
rect 5396 56382 5482 56438
rect 5538 56382 5624 56438
rect 5680 56382 5766 56438
rect 5822 56382 5908 56438
rect 5964 56382 6050 56438
rect 6106 56382 6192 56438
rect 6248 56382 6334 56438
rect 6390 56382 6476 56438
rect 6532 56382 6618 56438
rect 6674 56382 6760 56438
rect 6816 56382 6902 56438
rect 6958 56382 7044 56438
rect 7100 56382 7186 56438
rect 7242 56382 7328 56438
rect 7384 56382 7470 56438
rect 7526 56382 7612 56438
rect 7668 56382 7754 56438
rect 7810 56382 7896 56438
rect 7952 56382 8038 56438
rect 8094 56382 8180 56438
rect 8236 56382 8322 56438
rect 8378 56382 8464 56438
rect 8520 56382 8606 56438
rect 8662 56382 8748 56438
rect 8804 56382 8890 56438
rect 8946 56382 9032 56438
rect 9088 56382 9174 56438
rect 9230 56382 9316 56438
rect 9372 56382 9458 56438
rect 9514 56382 9600 56438
rect 9656 56382 9742 56438
rect 9798 56382 9884 56438
rect 9940 56382 10026 56438
rect 10082 56382 10168 56438
rect 10224 56382 10310 56438
rect 10366 56382 10452 56438
rect 10508 56382 10594 56438
rect 10650 56382 10736 56438
rect 10792 56382 10878 56438
rect 10934 56382 11020 56438
rect 11076 56382 11162 56438
rect 11218 56382 11304 56438
rect 11360 56382 11446 56438
rect 11502 56382 11588 56438
rect 11644 56382 11730 56438
rect 11786 56382 11872 56438
rect 11928 56382 12014 56438
rect 12070 56382 12156 56438
rect 12212 56382 12298 56438
rect 12354 56382 12440 56438
rect 12496 56382 12582 56438
rect 12638 56382 12724 56438
rect 12780 56382 12866 56438
rect 12922 56382 13008 56438
rect 13064 56382 13150 56438
rect 13206 56382 13292 56438
rect 13348 56382 13434 56438
rect 13490 56382 13576 56438
rect 13632 56382 13642 56438
rect 2490 56296 13642 56382
rect 2490 56240 2500 56296
rect 2556 56240 2642 56296
rect 2698 56240 2784 56296
rect 2840 56240 2926 56296
rect 2982 56240 3068 56296
rect 3124 56240 3210 56296
rect 3266 56240 3352 56296
rect 3408 56240 3494 56296
rect 3550 56240 3636 56296
rect 3692 56240 3778 56296
rect 3834 56240 3920 56296
rect 3976 56240 4062 56296
rect 4118 56240 4204 56296
rect 4260 56240 4346 56296
rect 4402 56240 4488 56296
rect 4544 56240 4630 56296
rect 4686 56240 4772 56296
rect 4828 56240 4914 56296
rect 4970 56240 5056 56296
rect 5112 56240 5198 56296
rect 5254 56240 5340 56296
rect 5396 56240 5482 56296
rect 5538 56240 5624 56296
rect 5680 56240 5766 56296
rect 5822 56240 5908 56296
rect 5964 56240 6050 56296
rect 6106 56240 6192 56296
rect 6248 56240 6334 56296
rect 6390 56240 6476 56296
rect 6532 56240 6618 56296
rect 6674 56240 6760 56296
rect 6816 56240 6902 56296
rect 6958 56240 7044 56296
rect 7100 56240 7186 56296
rect 7242 56240 7328 56296
rect 7384 56240 7470 56296
rect 7526 56240 7612 56296
rect 7668 56240 7754 56296
rect 7810 56240 7896 56296
rect 7952 56240 8038 56296
rect 8094 56240 8180 56296
rect 8236 56240 8322 56296
rect 8378 56240 8464 56296
rect 8520 56240 8606 56296
rect 8662 56240 8748 56296
rect 8804 56240 8890 56296
rect 8946 56240 9032 56296
rect 9088 56240 9174 56296
rect 9230 56240 9316 56296
rect 9372 56240 9458 56296
rect 9514 56240 9600 56296
rect 9656 56240 9742 56296
rect 9798 56240 9884 56296
rect 9940 56240 10026 56296
rect 10082 56240 10168 56296
rect 10224 56240 10310 56296
rect 10366 56240 10452 56296
rect 10508 56240 10594 56296
rect 10650 56240 10736 56296
rect 10792 56240 10878 56296
rect 10934 56240 11020 56296
rect 11076 56240 11162 56296
rect 11218 56240 11304 56296
rect 11360 56240 11446 56296
rect 11502 56240 11588 56296
rect 11644 56240 11730 56296
rect 11786 56240 11872 56296
rect 11928 56240 12014 56296
rect 12070 56240 12156 56296
rect 12212 56240 12298 56296
rect 12354 56240 12440 56296
rect 12496 56240 12582 56296
rect 12638 56240 12724 56296
rect 12780 56240 12866 56296
rect 12922 56240 13008 56296
rect 13064 56240 13150 56296
rect 13206 56240 13292 56296
rect 13348 56240 13434 56296
rect 13490 56240 13576 56296
rect 13632 56240 13642 56296
rect 2490 56154 13642 56240
rect 2490 56098 2500 56154
rect 2556 56098 2642 56154
rect 2698 56098 2784 56154
rect 2840 56098 2926 56154
rect 2982 56098 3068 56154
rect 3124 56098 3210 56154
rect 3266 56098 3352 56154
rect 3408 56098 3494 56154
rect 3550 56098 3636 56154
rect 3692 56098 3778 56154
rect 3834 56098 3920 56154
rect 3976 56098 4062 56154
rect 4118 56098 4204 56154
rect 4260 56098 4346 56154
rect 4402 56098 4488 56154
rect 4544 56098 4630 56154
rect 4686 56098 4772 56154
rect 4828 56098 4914 56154
rect 4970 56098 5056 56154
rect 5112 56098 5198 56154
rect 5254 56098 5340 56154
rect 5396 56098 5482 56154
rect 5538 56098 5624 56154
rect 5680 56098 5766 56154
rect 5822 56098 5908 56154
rect 5964 56098 6050 56154
rect 6106 56098 6192 56154
rect 6248 56098 6334 56154
rect 6390 56098 6476 56154
rect 6532 56098 6618 56154
rect 6674 56098 6760 56154
rect 6816 56098 6902 56154
rect 6958 56098 7044 56154
rect 7100 56098 7186 56154
rect 7242 56098 7328 56154
rect 7384 56098 7470 56154
rect 7526 56098 7612 56154
rect 7668 56098 7754 56154
rect 7810 56098 7896 56154
rect 7952 56098 8038 56154
rect 8094 56098 8180 56154
rect 8236 56098 8322 56154
rect 8378 56098 8464 56154
rect 8520 56098 8606 56154
rect 8662 56098 8748 56154
rect 8804 56098 8890 56154
rect 8946 56098 9032 56154
rect 9088 56098 9174 56154
rect 9230 56098 9316 56154
rect 9372 56098 9458 56154
rect 9514 56098 9600 56154
rect 9656 56098 9742 56154
rect 9798 56098 9884 56154
rect 9940 56098 10026 56154
rect 10082 56098 10168 56154
rect 10224 56098 10310 56154
rect 10366 56098 10452 56154
rect 10508 56098 10594 56154
rect 10650 56098 10736 56154
rect 10792 56098 10878 56154
rect 10934 56098 11020 56154
rect 11076 56098 11162 56154
rect 11218 56098 11304 56154
rect 11360 56098 11446 56154
rect 11502 56098 11588 56154
rect 11644 56098 11730 56154
rect 11786 56098 11872 56154
rect 11928 56098 12014 56154
rect 12070 56098 12156 56154
rect 12212 56098 12298 56154
rect 12354 56098 12440 56154
rect 12496 56098 12582 56154
rect 12638 56098 12724 56154
rect 12780 56098 12866 56154
rect 12922 56098 13008 56154
rect 13064 56098 13150 56154
rect 13206 56098 13292 56154
rect 13348 56098 13434 56154
rect 13490 56098 13576 56154
rect 13632 56098 13642 56154
rect 2490 56088 13642 56098
rect 1886 56033 1962 56043
rect 4938 55751 5014 55761
rect 4750 55741 4826 55751
rect 4750 55685 4760 55741
rect 4816 55685 4826 55741
rect 4750 55599 4826 55685
rect 4750 55543 4760 55599
rect 4816 55543 4826 55599
rect 4750 55457 4826 55543
rect 4750 55401 4760 55457
rect 4816 55401 4826 55457
rect 4750 55315 4826 55401
rect 4750 55259 4760 55315
rect 4816 55259 4826 55315
rect 4750 55173 4826 55259
rect 4750 55117 4760 55173
rect 4816 55117 4826 55173
rect 4750 55031 4826 55117
rect 4750 54975 4760 55031
rect 4816 54975 4826 55031
rect 4938 55695 4948 55751
rect 5004 55695 5014 55751
rect 4938 55609 5014 55695
rect 4938 55553 4948 55609
rect 5004 55553 5014 55609
rect 4938 55467 5014 55553
rect 4938 55411 4948 55467
rect 5004 55411 5014 55467
rect 4938 55325 5014 55411
rect 4938 55269 4948 55325
rect 5004 55269 5014 55325
rect 4938 55183 5014 55269
rect 4938 55127 4948 55183
rect 5004 55127 5014 55183
rect 4938 55041 5014 55127
rect 4938 54985 4948 55041
rect 5004 54985 5014 55041
rect 4938 54975 5014 54985
rect 5426 55760 5502 55770
rect 5426 55704 5436 55760
rect 5492 55704 5502 55760
rect 5426 55618 5502 55704
rect 5426 55562 5436 55618
rect 5492 55562 5502 55618
rect 5426 55476 5502 55562
rect 5426 55420 5436 55476
rect 5492 55420 5502 55476
rect 5426 55334 5502 55420
rect 5426 55278 5436 55334
rect 5492 55278 5502 55334
rect 5426 55192 5502 55278
rect 5426 55136 5436 55192
rect 5492 55136 5502 55192
rect 5426 55050 5502 55136
rect 5426 54994 5436 55050
rect 5492 54994 5502 55050
rect 5426 54984 5502 54994
rect 5914 55760 5990 55770
rect 5914 55704 5924 55760
rect 5980 55704 5990 55760
rect 6278 55760 6354 55770
rect 5914 55618 5990 55704
rect 5914 55562 5924 55618
rect 5980 55562 5990 55618
rect 5914 55476 5990 55562
rect 5914 55420 5924 55476
rect 5980 55420 5990 55476
rect 5914 55334 5990 55420
rect 5914 55278 5924 55334
rect 5980 55278 5990 55334
rect 5914 55192 5990 55278
rect 5914 55136 5924 55192
rect 5980 55136 5990 55192
rect 5914 55050 5990 55136
rect 5914 54994 5924 55050
rect 5980 54994 5990 55050
rect 5914 54984 5990 54994
rect 6096 55741 6172 55751
rect 6096 55685 6106 55741
rect 6162 55685 6172 55741
rect 6096 55599 6172 55685
rect 6096 55543 6106 55599
rect 6162 55543 6172 55599
rect 6096 55457 6172 55543
rect 6096 55401 6106 55457
rect 6162 55401 6172 55457
rect 6096 55315 6172 55401
rect 6096 55259 6106 55315
rect 6162 55259 6172 55315
rect 6096 55173 6172 55259
rect 6096 55117 6106 55173
rect 6162 55117 6172 55173
rect 6096 55031 6172 55117
rect 6096 54975 6106 55031
rect 6162 54975 6172 55031
rect 6278 55704 6288 55760
rect 6344 55704 6354 55760
rect 6278 55618 6354 55704
rect 6278 55562 6288 55618
rect 6344 55562 6354 55618
rect 6278 55476 6354 55562
rect 6278 55420 6288 55476
rect 6344 55420 6354 55476
rect 6278 55334 6354 55420
rect 6278 55278 6288 55334
rect 6344 55278 6354 55334
rect 6278 55192 6354 55278
rect 6278 55136 6288 55192
rect 6344 55136 6354 55192
rect 6278 55050 6354 55136
rect 6278 54994 6288 55050
rect 6344 54994 6354 55050
rect 6278 54984 6354 54994
rect 6766 55760 6842 55770
rect 6766 55704 6776 55760
rect 6832 55704 6842 55760
rect 6766 55618 6842 55704
rect 6766 55562 6776 55618
rect 6832 55562 6842 55618
rect 6766 55476 6842 55562
rect 6766 55420 6776 55476
rect 6832 55420 6842 55476
rect 6766 55334 6842 55420
rect 6766 55278 6776 55334
rect 6832 55278 6842 55334
rect 6766 55192 6842 55278
rect 6766 55136 6776 55192
rect 6832 55136 6842 55192
rect 6766 55050 6842 55136
rect 6766 54994 6776 55050
rect 6832 54994 6842 55050
rect 6766 54984 6842 54994
rect 7254 55760 7330 55770
rect 7254 55704 7264 55760
rect 7320 55704 7330 55760
rect 10182 55760 10258 55770
rect 7254 55618 7330 55704
rect 7254 55562 7264 55618
rect 7320 55562 7330 55618
rect 7254 55476 7330 55562
rect 7254 55420 7264 55476
rect 7320 55420 7330 55476
rect 7254 55334 7330 55420
rect 7254 55278 7264 55334
rect 7320 55278 7330 55334
rect 7254 55192 7330 55278
rect 7254 55136 7264 55192
rect 7320 55136 7330 55192
rect 7254 55050 7330 55136
rect 7254 54994 7264 55050
rect 7320 54994 7330 55050
rect 7254 54984 7330 54994
rect 7442 55741 7518 55751
rect 7442 55685 7452 55741
rect 7508 55685 7518 55741
rect 7442 55599 7518 55685
rect 7442 55543 7452 55599
rect 7508 55543 7518 55599
rect 7442 55457 7518 55543
rect 7442 55401 7452 55457
rect 7508 55401 7518 55457
rect 7442 55315 7518 55401
rect 7442 55259 7452 55315
rect 7508 55259 7518 55315
rect 7442 55173 7518 55259
rect 7442 55117 7452 55173
rect 7508 55117 7518 55173
rect 7442 55031 7518 55117
rect 4750 54889 4826 54975
rect 4750 54833 4760 54889
rect 4816 54833 4826 54889
rect 4750 54823 4826 54833
rect 6096 54889 6172 54975
rect 6096 54833 6106 54889
rect 6162 54833 6172 54889
rect 6096 54823 6172 54833
rect 7442 54975 7452 55031
rect 7508 54975 7518 55031
rect 7442 54889 7518 54975
rect 7442 54833 7452 54889
rect 7508 54833 7518 54889
rect 7442 54823 7518 54833
rect 9994 55741 10070 55751
rect 9994 55685 10004 55741
rect 10060 55685 10070 55741
rect 9994 55599 10070 55685
rect 9994 55543 10004 55599
rect 10060 55543 10070 55599
rect 9994 55457 10070 55543
rect 9994 55401 10004 55457
rect 10060 55401 10070 55457
rect 9994 55315 10070 55401
rect 9994 55259 10004 55315
rect 10060 55259 10070 55315
rect 9994 55173 10070 55259
rect 9994 55117 10004 55173
rect 10060 55117 10070 55173
rect 9994 55031 10070 55117
rect 9994 54975 10004 55031
rect 10060 54975 10070 55031
rect 10182 55704 10192 55760
rect 10248 55704 10258 55760
rect 10182 55618 10258 55704
rect 10182 55562 10192 55618
rect 10248 55562 10258 55618
rect 10182 55476 10258 55562
rect 10182 55420 10192 55476
rect 10248 55420 10258 55476
rect 10182 55334 10258 55420
rect 10182 55278 10192 55334
rect 10248 55278 10258 55334
rect 10182 55192 10258 55278
rect 10182 55136 10192 55192
rect 10248 55136 10258 55192
rect 10182 55050 10258 55136
rect 10182 54994 10192 55050
rect 10248 54994 10258 55050
rect 10182 54984 10258 54994
rect 10670 55760 10746 55770
rect 10670 55704 10680 55760
rect 10736 55704 10746 55760
rect 10670 55618 10746 55704
rect 10670 55562 10680 55618
rect 10736 55562 10746 55618
rect 10670 55476 10746 55562
rect 10670 55420 10680 55476
rect 10736 55420 10746 55476
rect 10670 55334 10746 55420
rect 10670 55278 10680 55334
rect 10736 55278 10746 55334
rect 10670 55192 10746 55278
rect 10670 55136 10680 55192
rect 10736 55136 10746 55192
rect 10670 55050 10746 55136
rect 10670 54994 10680 55050
rect 10736 54994 10746 55050
rect 10670 54984 10746 54994
rect 11158 55760 11234 55770
rect 11158 55704 11168 55760
rect 11224 55704 11234 55760
rect 11522 55760 11598 55770
rect 11158 55618 11234 55704
rect 11158 55562 11168 55618
rect 11224 55562 11234 55618
rect 11158 55476 11234 55562
rect 11158 55420 11168 55476
rect 11224 55420 11234 55476
rect 11158 55334 11234 55420
rect 11158 55278 11168 55334
rect 11224 55278 11234 55334
rect 11158 55192 11234 55278
rect 11158 55136 11168 55192
rect 11224 55136 11234 55192
rect 11158 55050 11234 55136
rect 11158 54994 11168 55050
rect 11224 54994 11234 55050
rect 11158 54984 11234 54994
rect 11340 55741 11416 55751
rect 11340 55685 11350 55741
rect 11406 55685 11416 55741
rect 11340 55599 11416 55685
rect 11340 55543 11350 55599
rect 11406 55543 11416 55599
rect 11340 55457 11416 55543
rect 11340 55401 11350 55457
rect 11406 55401 11416 55457
rect 11340 55315 11416 55401
rect 11340 55259 11350 55315
rect 11406 55259 11416 55315
rect 11340 55173 11416 55259
rect 11340 55117 11350 55173
rect 11406 55117 11416 55173
rect 11340 55031 11416 55117
rect 9994 54889 10070 54975
rect 9994 54833 10004 54889
rect 10060 54833 10070 54889
rect 9994 54823 10070 54833
rect 11340 54975 11350 55031
rect 11406 54975 11416 55031
rect 11522 55704 11532 55760
rect 11588 55704 11598 55760
rect 11522 55618 11598 55704
rect 11522 55562 11532 55618
rect 11588 55562 11598 55618
rect 11522 55476 11598 55562
rect 11522 55420 11532 55476
rect 11588 55420 11598 55476
rect 11522 55334 11598 55420
rect 11522 55278 11532 55334
rect 11588 55278 11598 55334
rect 11522 55192 11598 55278
rect 11522 55136 11532 55192
rect 11588 55136 11598 55192
rect 11522 55050 11598 55136
rect 11522 54994 11532 55050
rect 11588 54994 11598 55050
rect 11522 54984 11598 54994
rect 12010 55760 12086 55770
rect 12010 55704 12020 55760
rect 12076 55704 12086 55760
rect 12010 55618 12086 55704
rect 12010 55562 12020 55618
rect 12076 55562 12086 55618
rect 12010 55476 12086 55562
rect 12010 55420 12020 55476
rect 12076 55420 12086 55476
rect 12010 55334 12086 55420
rect 12010 55278 12020 55334
rect 12076 55278 12086 55334
rect 12010 55192 12086 55278
rect 12010 55136 12020 55192
rect 12076 55136 12086 55192
rect 12010 55050 12086 55136
rect 12010 54994 12020 55050
rect 12076 54994 12086 55050
rect 12010 54984 12086 54994
rect 12498 55760 12574 55770
rect 12498 55704 12508 55760
rect 12564 55704 12574 55760
rect 14400 55767 14760 55777
rect 12498 55618 12574 55704
rect 12498 55562 12508 55618
rect 12564 55562 12574 55618
rect 12498 55476 12574 55562
rect 12498 55420 12508 55476
rect 12564 55420 12574 55476
rect 12498 55334 12574 55420
rect 12498 55278 12508 55334
rect 12564 55278 12574 55334
rect 12498 55192 12574 55278
rect 12498 55136 12508 55192
rect 12564 55136 12574 55192
rect 12498 55050 12574 55136
rect 12498 54994 12508 55050
rect 12564 54994 12574 55050
rect 12498 54984 12574 54994
rect 12686 55741 12762 55751
rect 12686 55685 12696 55741
rect 12752 55685 12762 55741
rect 12686 55599 12762 55685
rect 12686 55543 12696 55599
rect 12752 55543 12762 55599
rect 12686 55457 12762 55543
rect 12686 55401 12696 55457
rect 12752 55401 12762 55457
rect 12686 55315 12762 55401
rect 12686 55259 12696 55315
rect 12752 55259 12762 55315
rect 12686 55173 12762 55259
rect 12686 55117 12696 55173
rect 12752 55117 12762 55173
rect 12686 55031 12762 55117
rect 11340 54889 11416 54975
rect 11340 54833 11350 54889
rect 11406 54833 11416 54889
rect 11340 54823 11416 54833
rect 12686 54975 12696 55031
rect 12752 54975 12762 55031
rect 12686 54889 12762 54975
rect 12686 54833 12696 54889
rect 12752 54833 12762 54889
rect 12686 54823 12762 54833
rect 14400 55711 14410 55767
rect 14466 55711 14552 55767
rect 14608 55711 14694 55767
rect 14750 55711 14760 55767
rect 14400 55625 14760 55711
rect 14400 55569 14410 55625
rect 14466 55569 14552 55625
rect 14608 55569 14694 55625
rect 14750 55569 14760 55625
rect 14400 55483 14760 55569
rect 14400 55427 14410 55483
rect 14466 55427 14552 55483
rect 14608 55427 14694 55483
rect 14750 55427 14760 55483
rect 14400 55341 14760 55427
rect 14400 55285 14410 55341
rect 14466 55285 14552 55341
rect 14608 55285 14694 55341
rect 14750 55285 14760 55341
rect 14400 55199 14760 55285
rect 14400 55143 14410 55199
rect 14466 55143 14552 55199
rect 14608 55143 14694 55199
rect 14750 55143 14760 55199
rect 14400 55057 14760 55143
rect 14400 55001 14410 55057
rect 14466 55001 14552 55057
rect 14608 55001 14694 55057
rect 14750 55001 14760 55057
rect 14400 54915 14760 55001
rect 14400 54859 14410 54915
rect 14466 54859 14552 54915
rect 14608 54859 14694 54915
rect 14750 54859 14760 54915
rect 14400 54773 14760 54859
rect 14400 54717 14410 54773
rect 14466 54717 14552 54773
rect 14608 54717 14694 54773
rect 14750 54717 14760 54773
rect 14400 54631 14760 54717
rect 14400 54575 14410 54631
rect 14466 54575 14552 54631
rect 14608 54575 14694 54631
rect 14750 54575 14760 54631
rect 14400 54489 14760 54575
rect 14400 54433 14410 54489
rect 14466 54433 14552 54489
rect 14608 54433 14694 54489
rect 14750 54433 14760 54489
rect 14400 54423 14760 54433
rect 1886 54160 1962 54170
rect 1886 54104 1896 54160
rect 1952 54104 1962 54160
rect 1886 54018 1962 54104
rect 1886 53962 1896 54018
rect 1952 53962 1962 54018
rect 1886 53876 1962 53962
rect 1886 53820 1896 53876
rect 1952 53820 1962 53876
rect 1886 53734 1962 53820
rect 1886 53678 1896 53734
rect 1952 53678 1962 53734
rect 1886 53592 1962 53678
rect 1886 53536 1896 53592
rect 1952 53536 1962 53592
rect 1886 53450 1962 53536
rect 1886 53394 1896 53450
rect 1952 53394 1962 53450
rect 1886 53308 1962 53394
rect 1886 53252 1896 53308
rect 1952 53252 1962 53308
rect 1886 53166 1962 53252
rect 4750 54160 4826 54170
rect 4750 54104 4760 54160
rect 4816 54104 4826 54160
rect 6096 54160 6172 54170
rect 4750 54018 4826 54104
rect 4750 53962 4760 54018
rect 4816 53962 4826 54018
rect 4750 53876 4826 53962
rect 4750 53820 4760 53876
rect 4816 53820 4826 53876
rect 4750 53734 4826 53820
rect 4750 53678 4760 53734
rect 4816 53678 4826 53734
rect 4750 53592 4826 53678
rect 4750 53536 4760 53592
rect 4816 53536 4826 53592
rect 4750 53450 4826 53536
rect 4750 53394 4760 53450
rect 4816 53394 4826 53450
rect 4750 53308 4826 53394
rect 4938 54099 5014 54109
rect 4938 54043 4948 54099
rect 5004 54043 5014 54099
rect 4938 53957 5014 54043
rect 4938 53901 4948 53957
rect 5004 53901 5014 53957
rect 4938 53815 5014 53901
rect 4938 53759 4948 53815
rect 5004 53759 5014 53815
rect 4938 53673 5014 53759
rect 4938 53617 4948 53673
rect 5004 53617 5014 53673
rect 4938 53531 5014 53617
rect 4938 53475 4948 53531
rect 5004 53475 5014 53531
rect 4938 53389 5014 53475
rect 4938 53333 4948 53389
rect 5004 53333 5014 53389
rect 4938 53323 5014 53333
rect 5426 54099 5502 54109
rect 5426 54043 5436 54099
rect 5492 54043 5502 54099
rect 5426 53957 5502 54043
rect 5426 53901 5436 53957
rect 5492 53901 5502 53957
rect 5426 53815 5502 53901
rect 5426 53759 5436 53815
rect 5492 53759 5502 53815
rect 5426 53673 5502 53759
rect 5426 53617 5436 53673
rect 5492 53617 5502 53673
rect 5426 53531 5502 53617
rect 5426 53475 5436 53531
rect 5492 53475 5502 53531
rect 5426 53389 5502 53475
rect 5426 53333 5436 53389
rect 5492 53333 5502 53389
rect 5426 53323 5502 53333
rect 5914 54099 5990 54109
rect 5914 54043 5924 54099
rect 5980 54043 5990 54099
rect 5914 53957 5990 54043
rect 5914 53901 5924 53957
rect 5980 53901 5990 53957
rect 5914 53815 5990 53901
rect 5914 53759 5924 53815
rect 5980 53759 5990 53815
rect 5914 53673 5990 53759
rect 5914 53617 5924 53673
rect 5980 53617 5990 53673
rect 5914 53531 5990 53617
rect 5914 53475 5924 53531
rect 5980 53475 5990 53531
rect 5914 53389 5990 53475
rect 5914 53333 5924 53389
rect 5980 53333 5990 53389
rect 5914 53323 5990 53333
rect 6096 54104 6106 54160
rect 6162 54104 6172 54160
rect 7442 54160 7518 54170
rect 6096 54018 6172 54104
rect 6096 53962 6106 54018
rect 6162 53962 6172 54018
rect 6096 53876 6172 53962
rect 6096 53820 6106 53876
rect 6162 53820 6172 53876
rect 6096 53734 6172 53820
rect 6096 53678 6106 53734
rect 6162 53678 6172 53734
rect 6096 53592 6172 53678
rect 6096 53536 6106 53592
rect 6162 53536 6172 53592
rect 6096 53450 6172 53536
rect 6096 53394 6106 53450
rect 6162 53394 6172 53450
rect 4750 53252 4760 53308
rect 4816 53252 4826 53308
rect 4750 53242 4826 53252
rect 6096 53308 6172 53394
rect 6278 54099 6354 54109
rect 6278 54043 6288 54099
rect 6344 54043 6354 54099
rect 6278 53957 6354 54043
rect 6278 53901 6288 53957
rect 6344 53901 6354 53957
rect 6278 53815 6354 53901
rect 6278 53759 6288 53815
rect 6344 53759 6354 53815
rect 6278 53673 6354 53759
rect 6278 53617 6288 53673
rect 6344 53617 6354 53673
rect 6278 53531 6354 53617
rect 6278 53475 6288 53531
rect 6344 53475 6354 53531
rect 6278 53389 6354 53475
rect 6278 53333 6288 53389
rect 6344 53333 6354 53389
rect 6278 53323 6354 53333
rect 6766 54099 6842 54109
rect 6766 54043 6776 54099
rect 6832 54043 6842 54099
rect 6766 53957 6842 54043
rect 6766 53901 6776 53957
rect 6832 53901 6842 53957
rect 6766 53815 6842 53901
rect 6766 53759 6776 53815
rect 6832 53759 6842 53815
rect 6766 53673 6842 53759
rect 6766 53617 6776 53673
rect 6832 53617 6842 53673
rect 6766 53531 6842 53617
rect 6766 53475 6776 53531
rect 6832 53475 6842 53531
rect 6766 53389 6842 53475
rect 6766 53333 6776 53389
rect 6832 53333 6842 53389
rect 6766 53323 6842 53333
rect 7254 54099 7330 54109
rect 7254 54043 7264 54099
rect 7320 54043 7330 54099
rect 7254 53957 7330 54043
rect 7254 53901 7264 53957
rect 7320 53901 7330 53957
rect 7254 53815 7330 53901
rect 7254 53759 7264 53815
rect 7320 53759 7330 53815
rect 7254 53673 7330 53759
rect 7254 53617 7264 53673
rect 7320 53617 7330 53673
rect 7254 53531 7330 53617
rect 7254 53475 7264 53531
rect 7320 53475 7330 53531
rect 7254 53389 7330 53475
rect 7254 53333 7264 53389
rect 7320 53333 7330 53389
rect 7254 53323 7330 53333
rect 7442 54104 7452 54160
rect 7508 54104 7518 54160
rect 7442 54018 7518 54104
rect 7442 53962 7452 54018
rect 7508 53962 7518 54018
rect 7442 53876 7518 53962
rect 7442 53820 7452 53876
rect 7508 53820 7518 53876
rect 7442 53734 7518 53820
rect 7442 53678 7452 53734
rect 7508 53678 7518 53734
rect 7442 53592 7518 53678
rect 7442 53536 7452 53592
rect 7508 53536 7518 53592
rect 7442 53450 7518 53536
rect 7442 53394 7452 53450
rect 7508 53394 7518 53450
rect 6096 53252 6106 53308
rect 6162 53252 6172 53308
rect 6096 53242 6172 53252
rect 7442 53308 7518 53394
rect 7442 53252 7452 53308
rect 7508 53252 7518 53308
rect 7442 53242 7518 53252
rect 9169 54160 9529 54170
rect 9169 54104 9179 54160
rect 9235 54104 9321 54160
rect 9377 54104 9463 54160
rect 9519 54104 9529 54160
rect 9169 54018 9529 54104
rect 9169 53962 9179 54018
rect 9235 53962 9321 54018
rect 9377 53962 9463 54018
rect 9519 53962 9529 54018
rect 9169 53876 9529 53962
rect 9169 53820 9179 53876
rect 9235 53820 9321 53876
rect 9377 53820 9463 53876
rect 9519 53820 9529 53876
rect 9169 53734 9529 53820
rect 9169 53678 9179 53734
rect 9235 53678 9321 53734
rect 9377 53678 9463 53734
rect 9519 53678 9529 53734
rect 9169 53592 9529 53678
rect 9169 53536 9179 53592
rect 9235 53536 9321 53592
rect 9377 53536 9463 53592
rect 9519 53536 9529 53592
rect 9169 53450 9529 53536
rect 9169 53394 9179 53450
rect 9235 53394 9321 53450
rect 9377 53394 9463 53450
rect 9519 53394 9529 53450
rect 9169 53308 9529 53394
rect 9169 53252 9179 53308
rect 9235 53252 9321 53308
rect 9377 53252 9463 53308
rect 9519 53252 9529 53308
rect 1886 53110 1896 53166
rect 1952 53110 1962 53166
rect 1886 53024 1962 53110
rect 1886 52968 1896 53024
rect 1952 52968 1962 53024
rect 1886 52882 1962 52968
rect 1886 52826 1896 52882
rect 1952 52826 1962 52882
rect 1886 52816 1962 52826
rect 9169 53166 9529 53252
rect 9994 54160 10070 54170
rect 9994 54104 10004 54160
rect 10060 54104 10070 54160
rect 11340 54160 11416 54170
rect 9994 54018 10070 54104
rect 9994 53962 10004 54018
rect 10060 53962 10070 54018
rect 9994 53876 10070 53962
rect 9994 53820 10004 53876
rect 10060 53820 10070 53876
rect 9994 53734 10070 53820
rect 9994 53678 10004 53734
rect 10060 53678 10070 53734
rect 9994 53592 10070 53678
rect 9994 53536 10004 53592
rect 10060 53536 10070 53592
rect 9994 53450 10070 53536
rect 9994 53394 10004 53450
rect 10060 53394 10070 53450
rect 9994 53308 10070 53394
rect 10182 54099 10258 54109
rect 10182 54043 10192 54099
rect 10248 54043 10258 54099
rect 10182 53957 10258 54043
rect 10182 53901 10192 53957
rect 10248 53901 10258 53957
rect 10182 53815 10258 53901
rect 10182 53759 10192 53815
rect 10248 53759 10258 53815
rect 10182 53673 10258 53759
rect 10182 53617 10192 53673
rect 10248 53617 10258 53673
rect 10182 53531 10258 53617
rect 10182 53475 10192 53531
rect 10248 53475 10258 53531
rect 10182 53389 10258 53475
rect 10182 53333 10192 53389
rect 10248 53333 10258 53389
rect 10182 53323 10258 53333
rect 10670 54099 10746 54109
rect 10670 54043 10680 54099
rect 10736 54043 10746 54099
rect 10670 53957 10746 54043
rect 10670 53901 10680 53957
rect 10736 53901 10746 53957
rect 10670 53815 10746 53901
rect 10670 53759 10680 53815
rect 10736 53759 10746 53815
rect 10670 53673 10746 53759
rect 10670 53617 10680 53673
rect 10736 53617 10746 53673
rect 10670 53531 10746 53617
rect 10670 53475 10680 53531
rect 10736 53475 10746 53531
rect 10670 53389 10746 53475
rect 10670 53333 10680 53389
rect 10736 53333 10746 53389
rect 10670 53323 10746 53333
rect 11158 54099 11234 54109
rect 11158 54043 11168 54099
rect 11224 54043 11234 54099
rect 11158 53957 11234 54043
rect 11158 53901 11168 53957
rect 11224 53901 11234 53957
rect 11158 53815 11234 53901
rect 11158 53759 11168 53815
rect 11224 53759 11234 53815
rect 11158 53673 11234 53759
rect 11158 53617 11168 53673
rect 11224 53617 11234 53673
rect 11158 53531 11234 53617
rect 11158 53475 11168 53531
rect 11224 53475 11234 53531
rect 11158 53389 11234 53475
rect 11158 53333 11168 53389
rect 11224 53333 11234 53389
rect 11158 53323 11234 53333
rect 11340 54104 11350 54160
rect 11406 54104 11416 54160
rect 12686 54160 12762 54170
rect 11340 54018 11416 54104
rect 11340 53962 11350 54018
rect 11406 53962 11416 54018
rect 11340 53876 11416 53962
rect 11340 53820 11350 53876
rect 11406 53820 11416 53876
rect 11340 53734 11416 53820
rect 11340 53678 11350 53734
rect 11406 53678 11416 53734
rect 11340 53592 11416 53678
rect 11340 53536 11350 53592
rect 11406 53536 11416 53592
rect 11340 53450 11416 53536
rect 11340 53394 11350 53450
rect 11406 53394 11416 53450
rect 9994 53252 10004 53308
rect 10060 53252 10070 53308
rect 9994 53242 10070 53252
rect 11340 53308 11416 53394
rect 11522 54099 11598 54109
rect 11522 54043 11532 54099
rect 11588 54043 11598 54099
rect 11522 53957 11598 54043
rect 11522 53901 11532 53957
rect 11588 53901 11598 53957
rect 11522 53815 11598 53901
rect 11522 53759 11532 53815
rect 11588 53759 11598 53815
rect 11522 53673 11598 53759
rect 11522 53617 11532 53673
rect 11588 53617 11598 53673
rect 11522 53531 11598 53617
rect 11522 53475 11532 53531
rect 11588 53475 11598 53531
rect 11522 53389 11598 53475
rect 11522 53333 11532 53389
rect 11588 53333 11598 53389
rect 11522 53323 11598 53333
rect 12010 54099 12086 54109
rect 12010 54043 12020 54099
rect 12076 54043 12086 54099
rect 12010 53957 12086 54043
rect 12010 53901 12020 53957
rect 12076 53901 12086 53957
rect 12010 53815 12086 53901
rect 12010 53759 12020 53815
rect 12076 53759 12086 53815
rect 12010 53673 12086 53759
rect 12010 53617 12020 53673
rect 12076 53617 12086 53673
rect 12010 53531 12086 53617
rect 12010 53475 12020 53531
rect 12076 53475 12086 53531
rect 12010 53389 12086 53475
rect 12010 53333 12020 53389
rect 12076 53333 12086 53389
rect 12010 53323 12086 53333
rect 12498 54099 12574 54109
rect 12498 54043 12508 54099
rect 12564 54043 12574 54099
rect 12498 53957 12574 54043
rect 12498 53901 12508 53957
rect 12564 53901 12574 53957
rect 12498 53815 12574 53901
rect 12498 53759 12508 53815
rect 12564 53759 12574 53815
rect 12498 53673 12574 53759
rect 12498 53617 12508 53673
rect 12564 53617 12574 53673
rect 12498 53531 12574 53617
rect 12498 53475 12508 53531
rect 12564 53475 12574 53531
rect 12498 53389 12574 53475
rect 12498 53333 12508 53389
rect 12564 53333 12574 53389
rect 12498 53323 12574 53333
rect 12686 54104 12696 54160
rect 12752 54104 12762 54160
rect 12686 54018 12762 54104
rect 12686 53962 12696 54018
rect 12752 53962 12762 54018
rect 12686 53876 12762 53962
rect 12686 53820 12696 53876
rect 12752 53820 12762 53876
rect 12686 53734 12762 53820
rect 12686 53678 12696 53734
rect 12752 53678 12762 53734
rect 12686 53592 12762 53678
rect 12686 53536 12696 53592
rect 12752 53536 12762 53592
rect 12686 53450 12762 53536
rect 12686 53394 12696 53450
rect 12752 53394 12762 53450
rect 11340 53252 11350 53308
rect 11406 53252 11416 53308
rect 11340 53242 11416 53252
rect 12686 53308 12762 53394
rect 12686 53252 12696 53308
rect 12752 53252 12762 53308
rect 12686 53242 12762 53252
rect 9169 53110 9179 53166
rect 9235 53110 9321 53166
rect 9377 53110 9463 53166
rect 9519 53110 9529 53166
rect 9169 53024 9529 53110
rect 9169 52968 9179 53024
rect 9235 52968 9321 53024
rect 9377 52968 9463 53024
rect 9519 52968 9529 53024
rect 9169 52882 9529 52968
rect 9169 52826 9179 52882
rect 9235 52826 9321 52882
rect 9377 52826 9463 52882
rect 9519 52826 9529 52882
rect 9169 52816 9529 52826
rect 46 52567 122 52577
rect 46 52511 56 52567
rect 112 52511 122 52567
rect 46 52425 122 52511
rect 46 52369 56 52425
rect 112 52369 122 52425
rect 46 52283 122 52369
rect 46 52227 56 52283
rect 112 52227 122 52283
rect 46 52141 122 52227
rect 46 52085 56 52141
rect 112 52085 122 52141
rect 46 51999 122 52085
rect 46 51943 56 51999
rect 112 51943 122 51999
rect 46 51857 122 51943
rect 46 51801 56 51857
rect 112 51801 122 51857
rect 46 51715 122 51801
rect 46 51659 56 51715
rect 112 51659 122 51715
rect 46 51573 122 51659
rect 46 51517 56 51573
rect 112 51517 122 51573
rect 46 51431 122 51517
rect 46 51375 56 51431
rect 112 51375 122 51431
rect 46 51289 122 51375
rect 46 51233 56 51289
rect 112 51233 122 51289
rect 46 51223 122 51233
rect 724 52560 1084 52570
rect 724 52504 734 52560
rect 790 52504 876 52560
rect 932 52504 1018 52560
rect 1074 52504 1084 52560
rect 724 52418 1084 52504
rect 724 52362 734 52418
rect 790 52362 876 52418
rect 932 52362 1018 52418
rect 1074 52362 1084 52418
rect 724 52276 1084 52362
rect 724 52220 734 52276
rect 790 52220 876 52276
rect 932 52220 1018 52276
rect 1074 52220 1084 52276
rect 724 52134 1084 52220
rect 724 52078 734 52134
rect 790 52078 876 52134
rect 932 52078 1018 52134
rect 1074 52078 1084 52134
rect 724 51992 1084 52078
rect 724 51936 734 51992
rect 790 51936 876 51992
rect 932 51936 1018 51992
rect 1074 51936 1084 51992
rect 724 51850 1084 51936
rect 724 51794 734 51850
rect 790 51794 876 51850
rect 932 51794 1018 51850
rect 1074 51794 1084 51850
rect 724 51708 1084 51794
rect 724 51652 734 51708
rect 790 51652 876 51708
rect 932 51652 1018 51708
rect 1074 51652 1084 51708
rect 724 51566 1084 51652
rect 724 51510 734 51566
rect 790 51510 876 51566
rect 932 51510 1018 51566
rect 1074 51510 1084 51566
rect 724 51424 1084 51510
rect 724 51368 734 51424
rect 790 51368 876 51424
rect 932 51368 1018 51424
rect 1074 51368 1084 51424
rect 724 51282 1084 51368
rect 14942 52489 15018 52499
rect 14942 52433 14952 52489
rect 15008 52433 15018 52489
rect 14942 52347 15018 52433
rect 14942 52291 14952 52347
rect 15008 52291 15018 52347
rect 14942 52205 15018 52291
rect 14942 52149 14952 52205
rect 15008 52149 15018 52205
rect 14942 52063 15018 52149
rect 14942 52007 14952 52063
rect 15008 52007 15018 52063
rect 14942 51921 15018 52007
rect 14942 51865 14952 51921
rect 15008 51865 15018 51921
rect 14942 51779 15018 51865
rect 14942 51723 14952 51779
rect 15008 51723 15018 51779
rect 14942 51637 15018 51723
rect 14942 51581 14952 51637
rect 15008 51581 15018 51637
rect 14942 51495 15018 51581
rect 14942 51439 14952 51495
rect 15008 51439 15018 51495
rect 14942 51353 15018 51439
rect 14942 51297 14952 51353
rect 15008 51297 15018 51353
rect 14942 51287 15018 51297
rect 724 51226 734 51282
rect 790 51226 876 51282
rect 932 51226 1018 51282
rect 1074 51226 1084 51282
rect 724 51216 1084 51226
rect 204 50960 564 50970
rect 204 50904 214 50960
rect 270 50904 356 50960
rect 412 50904 498 50960
rect 554 50904 564 50960
rect 204 50818 564 50904
rect 204 50762 214 50818
rect 270 50762 356 50818
rect 412 50762 498 50818
rect 554 50762 564 50818
rect 204 50676 564 50762
rect 204 50620 214 50676
rect 270 50620 356 50676
rect 412 50620 498 50676
rect 554 50620 564 50676
rect 204 50534 564 50620
rect 204 50478 214 50534
rect 270 50478 356 50534
rect 412 50478 498 50534
rect 554 50478 564 50534
rect 204 50392 564 50478
rect 204 50336 214 50392
rect 270 50336 356 50392
rect 412 50336 498 50392
rect 554 50336 564 50392
rect 204 50250 564 50336
rect 204 50194 214 50250
rect 270 50194 356 50250
rect 412 50194 498 50250
rect 554 50194 564 50250
rect 204 50108 564 50194
rect 204 50052 214 50108
rect 270 50052 356 50108
rect 412 50052 498 50108
rect 554 50052 564 50108
rect 204 49966 564 50052
rect 204 49910 214 49966
rect 270 49910 356 49966
rect 412 49910 498 49966
rect 554 49910 564 49966
rect 204 49824 564 49910
rect 204 49768 214 49824
rect 270 49768 356 49824
rect 412 49768 498 49824
rect 554 49768 564 49824
rect 204 49682 564 49768
rect 204 49626 214 49682
rect 270 49626 356 49682
rect 412 49626 498 49682
rect 554 49626 564 49682
rect 204 49616 564 49626
rect 11574 49902 11762 49912
rect 11574 49846 11584 49902
rect 11640 49846 11696 49902
rect 11752 49846 11762 49902
rect 11574 49790 11762 49846
rect 11574 49734 11584 49790
rect 11640 49734 11696 49790
rect 11752 49734 11762 49790
rect 11574 49678 11762 49734
rect 11574 49622 11584 49678
rect 11640 49622 11696 49678
rect 11752 49622 11762 49678
rect 11574 49612 11762 49622
rect 10782 49360 10858 49370
rect 10782 49304 10792 49360
rect 10848 49304 10858 49360
rect 10782 49218 10858 49304
rect 10782 49162 10792 49218
rect 10848 49162 10858 49218
rect 10782 49076 10858 49162
rect 10782 49020 10792 49076
rect 10848 49020 10858 49076
rect 10782 48934 10858 49020
rect 10782 48878 10792 48934
rect 10848 48878 10858 48934
rect 10782 48792 10858 48878
rect 10782 48736 10792 48792
rect 10848 48736 10858 48792
rect 10782 48650 10858 48736
rect 10782 48594 10792 48650
rect 10848 48594 10858 48650
rect 10782 48508 10858 48594
rect 10782 48452 10792 48508
rect 10848 48452 10858 48508
rect 10782 48366 10858 48452
rect 10782 48310 10792 48366
rect 10848 48310 10858 48366
rect 10782 48300 10858 48310
rect 10424 48036 10604 48046
rect 10424 47980 10434 48036
rect 10594 47980 10604 48036
rect 10424 47970 10604 47980
rect 3608 47760 3684 47770
rect 3608 47704 3618 47760
rect 3674 47704 3684 47760
rect 14400 47760 14760 47770
rect 3608 47618 3684 47704
rect 3608 47562 3618 47618
rect 3674 47562 3684 47618
rect 3608 47476 3684 47562
rect 3608 47420 3618 47476
rect 3674 47420 3684 47476
rect 3608 47334 3684 47420
rect 3608 47278 3618 47334
rect 3674 47278 3684 47334
rect 3608 47192 3684 47278
rect 3608 47136 3618 47192
rect 3674 47136 3684 47192
rect 3608 47050 3684 47136
rect 11001 47744 11077 47754
rect 11001 47688 11011 47744
rect 11067 47688 11077 47744
rect 11001 47602 11077 47688
rect 11001 47546 11011 47602
rect 11067 47546 11077 47602
rect 11001 47460 11077 47546
rect 11001 47404 11011 47460
rect 11067 47404 11077 47460
rect 11001 47318 11077 47404
rect 11001 47262 11011 47318
rect 11067 47262 11077 47318
rect 11001 47176 11077 47262
rect 11001 47120 11011 47176
rect 11067 47120 11077 47176
rect 11001 47110 11077 47120
rect 14400 47704 14410 47760
rect 14466 47704 14552 47760
rect 14608 47704 14694 47760
rect 14750 47704 14760 47760
rect 14400 47618 14760 47704
rect 14400 47562 14410 47618
rect 14466 47562 14552 47618
rect 14608 47562 14694 47618
rect 14750 47562 14760 47618
rect 14400 47476 14760 47562
rect 14400 47420 14410 47476
rect 14466 47420 14552 47476
rect 14608 47420 14694 47476
rect 14750 47420 14760 47476
rect 14400 47334 14760 47420
rect 14400 47278 14410 47334
rect 14466 47278 14552 47334
rect 14608 47278 14694 47334
rect 14750 47278 14760 47334
rect 14400 47192 14760 47278
rect 14400 47136 14410 47192
rect 14466 47136 14552 47192
rect 14608 47136 14694 47192
rect 14750 47136 14760 47192
rect 3608 46994 3618 47050
rect 3674 46994 3684 47050
rect 3608 46908 3684 46994
rect 3608 46852 3618 46908
rect 3674 46852 3684 46908
rect 3608 46766 3684 46852
rect 3608 46710 3618 46766
rect 3674 46710 3684 46766
rect 3608 46700 3684 46710
rect 14400 47050 14760 47136
rect 14400 46994 14410 47050
rect 14466 46994 14552 47050
rect 14608 46994 14694 47050
rect 14750 46994 14760 47050
rect 14400 46908 14760 46994
rect 14400 46852 14410 46908
rect 14466 46852 14552 46908
rect 14608 46852 14694 46908
rect 14750 46852 14760 46908
rect 14400 46766 14760 46852
rect 14400 46710 14410 46766
rect 14466 46710 14552 46766
rect 14608 46710 14694 46766
rect 14750 46710 14760 46766
rect 14400 46624 14760 46710
rect 14400 46568 14410 46624
rect 14466 46568 14552 46624
rect 14608 46568 14694 46624
rect 14750 46568 14760 46624
rect 14400 46482 14760 46568
rect 14400 46426 14410 46482
rect 14466 46426 14552 46482
rect 14608 46426 14694 46482
rect 14750 46426 14760 46482
rect 14400 46416 14760 46426
rect 10888 46126 10964 46136
rect 10888 44822 10898 46126
rect 10954 44822 10964 46126
rect 10888 44812 10964 44822
rect 11017 46126 11093 46136
rect 11017 44822 11027 46126
rect 11083 44822 11093 46126
rect 11017 44812 11093 44822
rect 3608 44560 3684 44570
rect 3608 44504 3618 44560
rect 3674 44504 3684 44560
rect 3608 44418 3684 44504
rect 3608 44362 3618 44418
rect 3674 44362 3684 44418
rect 3608 44276 3684 44362
rect 3608 44220 3618 44276
rect 3674 44220 3684 44276
rect 3608 44134 3684 44220
rect 3608 44078 3618 44134
rect 3674 44078 3684 44134
rect 3608 43992 3684 44078
rect 3608 43936 3618 43992
rect 3674 43936 3684 43992
rect 3608 43850 3684 43936
rect 3608 43794 3618 43850
rect 3674 43794 3684 43850
rect 3608 43708 3684 43794
rect 3608 43652 3618 43708
rect 3674 43652 3684 43708
rect 3608 43566 3684 43652
rect 3608 43510 3618 43566
rect 3674 43510 3684 43566
rect 3608 43424 3684 43510
rect 3608 43368 3618 43424
rect 3674 43368 3684 43424
rect 3608 43282 3684 43368
rect 3608 43226 3618 43282
rect 3674 43226 3684 43282
rect 3608 43216 3684 43226
rect 3608 42960 3684 42970
rect 3608 42904 3618 42960
rect 3674 42904 3684 42960
rect 3608 42818 3684 42904
rect 3608 42762 3618 42818
rect 3674 42762 3684 42818
rect 3608 42676 3684 42762
rect 3608 42620 3618 42676
rect 3674 42620 3684 42676
rect 3608 42534 3684 42620
rect 3608 42478 3618 42534
rect 3674 42478 3684 42534
rect 3608 42392 3684 42478
rect 3608 42336 3618 42392
rect 3674 42336 3684 42392
rect 3608 42250 3684 42336
rect 3608 42194 3618 42250
rect 3674 42194 3684 42250
rect 3608 42108 3684 42194
rect 3608 42052 3618 42108
rect 3674 42052 3684 42108
rect 3608 41966 3684 42052
rect 3608 41910 3618 41966
rect 3674 41910 3684 41966
rect 3608 41824 3684 41910
rect 3608 41768 3618 41824
rect 3674 41768 3684 41824
rect 13181 42968 13481 42978
rect 13181 42912 13191 42968
rect 13247 42912 13303 42968
rect 13359 42912 13415 42968
rect 13471 42912 13481 42968
rect 13181 42856 13481 42912
rect 13181 42800 13191 42856
rect 13247 42800 13303 42856
rect 13359 42800 13415 42856
rect 13471 42800 13481 42856
rect 13181 42744 13481 42800
rect 13181 42688 13191 42744
rect 13247 42688 13303 42744
rect 13359 42688 13415 42744
rect 13471 42688 13481 42744
rect 13181 42632 13481 42688
rect 13181 42576 13191 42632
rect 13247 42576 13303 42632
rect 13359 42576 13415 42632
rect 13471 42576 13481 42632
rect 13181 42520 13481 42576
rect 13181 42464 13191 42520
rect 13247 42464 13303 42520
rect 13359 42464 13415 42520
rect 13471 42464 13481 42520
rect 13181 42408 13481 42464
rect 13181 42352 13191 42408
rect 13247 42352 13303 42408
rect 13359 42352 13415 42408
rect 13471 42352 13481 42408
rect 13181 42296 13481 42352
rect 13181 42240 13191 42296
rect 13247 42240 13303 42296
rect 13359 42240 13415 42296
rect 13471 42240 13481 42296
rect 13181 42184 13481 42240
rect 13181 42128 13191 42184
rect 13247 42128 13303 42184
rect 13359 42128 13415 42184
rect 13471 42128 13481 42184
rect 13181 42072 13481 42128
rect 13181 42016 13191 42072
rect 13247 42016 13303 42072
rect 13359 42016 13415 42072
rect 13471 42016 13481 42072
rect 13181 41960 13481 42016
rect 13181 41904 13191 41960
rect 13247 41904 13303 41960
rect 13359 41904 13415 41960
rect 13471 41904 13481 41960
rect 13181 41848 13481 41904
rect 13181 41792 13191 41848
rect 13247 41792 13303 41848
rect 13359 41792 13415 41848
rect 13471 41792 13481 41848
rect 13181 41782 13481 41792
rect 3608 41682 3684 41768
rect 3608 41626 3618 41682
rect 3674 41626 3684 41682
rect 3608 41616 3684 41626
rect 14400 41360 14760 41370
rect 14400 41304 14410 41360
rect 14466 41304 14552 41360
rect 14608 41304 14694 41360
rect 14750 41304 14760 41360
rect 14400 41218 14760 41304
rect 14400 41162 14410 41218
rect 14466 41162 14552 41218
rect 14608 41162 14694 41218
rect 14750 41162 14760 41218
rect 1836 41072 3758 41082
rect 1836 41016 1846 41072
rect 1902 41016 1988 41072
rect 2044 41016 2130 41072
rect 2186 41016 2272 41072
rect 2328 41016 2414 41072
rect 2470 41016 2556 41072
rect 2612 41016 2698 41072
rect 2754 41016 2840 41072
rect 2896 41016 2982 41072
rect 3038 41016 3124 41072
rect 3180 41016 3266 41072
rect 3322 41016 3408 41072
rect 3464 41016 3550 41072
rect 3606 41016 3692 41072
rect 3748 41016 3758 41072
rect 1836 41006 3758 41016
rect 14400 41076 14760 41162
rect 14400 41020 14410 41076
rect 14466 41020 14552 41076
rect 14608 41020 14694 41076
rect 14750 41020 14760 41076
rect 14400 40934 14760 41020
rect 14400 40878 14410 40934
rect 14466 40878 14552 40934
rect 14608 40878 14694 40934
rect 14750 40878 14760 40934
rect 14400 40792 14760 40878
rect 14400 40736 14410 40792
rect 14466 40736 14552 40792
rect 14608 40736 14694 40792
rect 14750 40736 14760 40792
rect 14400 40650 14760 40736
rect 14400 40594 14410 40650
rect 14466 40594 14552 40650
rect 14608 40594 14694 40650
rect 14750 40594 14760 40650
rect 14400 40508 14760 40594
rect 14400 40452 14410 40508
rect 14466 40452 14552 40508
rect 14608 40452 14694 40508
rect 14750 40452 14760 40508
rect 14400 40366 14760 40452
rect 2357 40316 4563 40326
rect 2357 40260 2367 40316
rect 2423 40260 2509 40316
rect 2565 40260 2651 40316
rect 2707 40260 2793 40316
rect 2849 40260 2935 40316
rect 2991 40260 3077 40316
rect 3133 40260 3219 40316
rect 3275 40260 3361 40316
rect 3417 40260 3503 40316
rect 3559 40260 3645 40316
rect 3701 40260 3787 40316
rect 3843 40260 3929 40316
rect 3985 40260 4071 40316
rect 4127 40260 4213 40316
rect 4269 40260 4355 40316
rect 4411 40260 4497 40316
rect 4553 40260 4563 40316
rect 2357 40250 4563 40260
rect 7987 40316 9767 40326
rect 7987 40260 7997 40316
rect 8053 40260 8139 40316
rect 8195 40260 8281 40316
rect 8337 40260 8423 40316
rect 8479 40260 8565 40316
rect 8621 40260 8707 40316
rect 8763 40260 8849 40316
rect 8905 40260 8991 40316
rect 9047 40260 9133 40316
rect 9189 40260 9275 40316
rect 9331 40260 9417 40316
rect 9473 40260 9559 40316
rect 9615 40260 9701 40316
rect 9757 40260 9767 40316
rect 7987 40250 9767 40260
rect 12748 40316 13818 40326
rect 12748 40260 12758 40316
rect 12814 40260 12900 40316
rect 12956 40260 13042 40316
rect 13098 40260 13184 40316
rect 13240 40260 13326 40316
rect 13382 40260 13468 40316
rect 13524 40260 13610 40316
rect 13666 40260 13752 40316
rect 13808 40260 13818 40316
rect 12748 40250 13818 40260
rect 14400 40310 14410 40366
rect 14466 40310 14552 40366
rect 14608 40310 14694 40366
rect 14750 40310 14760 40366
rect 14400 40224 14760 40310
rect 14400 40168 14410 40224
rect 14466 40168 14552 40224
rect 14608 40168 14694 40224
rect 14750 40168 14760 40224
rect 14400 40082 14760 40168
rect 14400 40026 14410 40082
rect 14466 40026 14552 40082
rect 14608 40026 14694 40082
rect 14750 40026 14760 40082
rect 14400 40016 14760 40026
rect 204 39760 564 39770
rect 204 39704 214 39760
rect 270 39704 356 39760
rect 412 39704 498 39760
rect 554 39704 564 39760
rect 204 39618 564 39704
rect 204 39562 214 39618
rect 270 39562 356 39618
rect 412 39562 498 39618
rect 554 39562 564 39618
rect 204 39476 564 39562
rect 204 39420 214 39476
rect 270 39420 356 39476
rect 412 39420 498 39476
rect 554 39420 564 39476
rect 204 39334 564 39420
rect 204 39278 214 39334
rect 270 39278 356 39334
rect 412 39278 498 39334
rect 554 39278 564 39334
rect 204 39192 564 39278
rect 204 39136 214 39192
rect 270 39136 356 39192
rect 412 39136 498 39192
rect 554 39136 564 39192
rect 204 39050 564 39136
rect 1771 39760 1847 39770
rect 1771 39704 1781 39760
rect 1837 39704 1847 39760
rect 1771 39618 1847 39704
rect 1771 39562 1781 39618
rect 1837 39562 1847 39618
rect 1771 39476 1847 39562
rect 1771 39420 1781 39476
rect 1837 39420 1847 39476
rect 1771 39334 1847 39420
rect 1771 39278 1781 39334
rect 1837 39278 1847 39334
rect 1771 39192 1847 39278
rect 1771 39136 1781 39192
rect 1837 39136 1847 39192
rect 1771 39126 1847 39136
rect 5083 39760 5159 39770
rect 5083 39704 5093 39760
rect 5149 39704 5159 39760
rect 5083 39618 5159 39704
rect 5083 39562 5093 39618
rect 5149 39562 5159 39618
rect 5083 39476 5159 39562
rect 5083 39420 5093 39476
rect 5149 39420 5159 39476
rect 5083 39334 5159 39420
rect 5083 39278 5093 39334
rect 5149 39278 5159 39334
rect 5083 39192 5159 39278
rect 5083 39136 5093 39192
rect 5149 39136 5159 39192
rect 5083 39126 5159 39136
rect 6049 39754 6125 39764
rect 6049 39698 6059 39754
rect 6115 39698 6125 39754
rect 6049 39612 6125 39698
rect 6049 39556 6059 39612
rect 6115 39556 6125 39612
rect 6049 39470 6125 39556
rect 6049 39414 6059 39470
rect 6115 39414 6125 39470
rect 6049 39328 6125 39414
rect 6049 39272 6059 39328
rect 6115 39272 6125 39328
rect 6049 39186 6125 39272
rect 6049 39130 6059 39186
rect 6115 39130 6125 39186
rect 204 38994 214 39050
rect 270 38994 356 39050
rect 412 38994 498 39050
rect 554 38994 564 39050
rect 204 38908 564 38994
rect 204 38852 214 38908
rect 270 38852 356 38908
rect 412 38852 498 38908
rect 554 38852 564 38908
rect 204 38766 564 38852
rect 204 38710 214 38766
rect 270 38710 356 38766
rect 412 38710 498 38766
rect 554 38710 564 38766
rect 204 38624 564 38710
rect 6049 39044 6125 39130
rect 7015 39760 7091 39770
rect 7015 39704 7025 39760
rect 7081 39704 7091 39760
rect 7015 39618 7091 39704
rect 7015 39562 7025 39618
rect 7081 39562 7091 39618
rect 7015 39476 7091 39562
rect 7015 39420 7025 39476
rect 7081 39420 7091 39476
rect 7015 39334 7091 39420
rect 7015 39278 7025 39334
rect 7081 39278 7091 39334
rect 7015 39192 7091 39278
rect 7015 39136 7025 39192
rect 7081 39136 7091 39192
rect 7015 39126 7091 39136
rect 10327 39760 10403 39770
rect 10327 39704 10337 39760
rect 10393 39704 10403 39760
rect 10327 39618 10403 39704
rect 10327 39562 10337 39618
rect 10393 39562 10403 39618
rect 10327 39476 10403 39562
rect 10327 39420 10337 39476
rect 10393 39420 10403 39476
rect 10327 39334 10403 39420
rect 10327 39278 10337 39334
rect 10393 39278 10403 39334
rect 10327 39192 10403 39278
rect 10327 39136 10337 39192
rect 10393 39136 10403 39192
rect 6049 38988 6059 39044
rect 6115 38988 6125 39044
rect 6049 38902 6125 38988
rect 6049 38846 6059 38902
rect 6115 38846 6125 38902
rect 6049 38760 6125 38846
rect 6049 38704 6059 38760
rect 6115 38704 6125 38760
rect 6049 38694 6125 38704
rect 10327 39050 10403 39136
rect 10327 38994 10337 39050
rect 10393 38994 10403 39050
rect 10327 38908 10403 38994
rect 10327 38852 10337 38908
rect 10393 38852 10403 38908
rect 10327 38766 10403 38852
rect 10327 38710 10337 38766
rect 10393 38710 10403 38766
rect 10327 38700 10403 38710
rect 11200 39760 11276 39770
rect 11200 39704 11210 39760
rect 11266 39704 11276 39760
rect 11200 39618 11276 39704
rect 11200 39562 11210 39618
rect 11266 39562 11276 39618
rect 11200 39476 11276 39562
rect 11200 39420 11210 39476
rect 11266 39420 11276 39476
rect 11200 39334 11276 39420
rect 11200 39278 11210 39334
rect 11266 39278 11276 39334
rect 11200 39192 11276 39278
rect 11200 39136 11210 39192
rect 11266 39136 11276 39192
rect 11200 39050 11276 39136
rect 11200 38994 11210 39050
rect 11266 38994 11276 39050
rect 11200 38908 11276 38994
rect 11200 38852 11210 38908
rect 11266 38852 11276 38908
rect 11200 38766 11276 38852
rect 11200 38710 11210 38766
rect 11266 38710 11276 38766
rect 11200 38700 11276 38710
rect 204 38568 214 38624
rect 270 38568 356 38624
rect 412 38568 498 38624
rect 554 38568 564 38624
rect 204 38482 564 38568
rect 204 38426 214 38482
rect 270 38426 356 38482
rect 412 38426 498 38482
rect 554 38426 564 38482
rect 204 38416 564 38426
rect 46 38167 122 38177
rect 46 38111 56 38167
rect 112 38111 122 38167
rect 46 38025 122 38111
rect 46 37969 56 38025
rect 112 37969 122 38025
rect 46 37883 122 37969
rect 46 37827 56 37883
rect 112 37827 122 37883
rect 46 37741 122 37827
rect 46 37685 56 37741
rect 112 37685 122 37741
rect 46 37599 122 37685
rect 46 37543 56 37599
rect 112 37543 122 37599
rect 46 37457 122 37543
rect 46 37401 56 37457
rect 112 37401 122 37457
rect 46 37315 122 37401
rect 46 37259 56 37315
rect 112 37259 122 37315
rect 46 37173 122 37259
rect 46 37117 56 37173
rect 112 37117 122 37173
rect 46 37031 122 37117
rect 46 36975 56 37031
rect 112 36975 122 37031
rect 46 36889 122 36975
rect 46 36833 56 36889
rect 112 36833 122 36889
rect 46 36823 122 36833
rect 724 38160 1084 38170
rect 724 38104 734 38160
rect 790 38104 876 38160
rect 932 38104 1018 38160
rect 1074 38104 1084 38160
rect 724 38018 1084 38104
rect 724 37962 734 38018
rect 790 37962 876 38018
rect 932 37962 1018 38018
rect 1074 37962 1084 38018
rect 724 37876 1084 37962
rect 724 37820 734 37876
rect 790 37820 876 37876
rect 932 37820 1018 37876
rect 1074 37820 1084 37876
rect 724 37734 1084 37820
rect 724 37678 734 37734
rect 790 37678 876 37734
rect 932 37678 1018 37734
rect 1074 37678 1084 37734
rect 724 37592 1084 37678
rect 724 37536 734 37592
rect 790 37536 876 37592
rect 932 37536 1018 37592
rect 1074 37536 1084 37592
rect 724 37450 1084 37536
rect 724 37394 734 37450
rect 790 37394 876 37450
rect 932 37394 1018 37450
rect 1074 37394 1084 37450
rect 724 37308 1084 37394
rect 724 37252 734 37308
rect 790 37252 876 37308
rect 932 37252 1018 37308
rect 1074 37252 1084 37308
rect 724 37166 1084 37252
rect 724 37110 734 37166
rect 790 37110 876 37166
rect 932 37110 1018 37166
rect 1074 37110 1084 37166
rect 724 37024 1084 37110
rect 724 36968 734 37024
rect 790 36968 876 37024
rect 932 36968 1018 37024
rect 1074 36968 1084 37024
rect 724 36882 1084 36968
rect 724 36826 734 36882
rect 790 36826 876 36882
rect 932 36826 1018 36882
rect 1074 36826 1084 36882
rect 724 36816 1084 36826
rect 6049 38160 6125 38170
rect 6049 38104 6059 38160
rect 6115 38104 6125 38160
rect 6049 38018 6125 38104
rect 6049 37962 6059 38018
rect 6115 37962 6125 38018
rect 6049 37876 6125 37962
rect 6049 37820 6059 37876
rect 6115 37820 6125 37876
rect 6049 37734 6125 37820
rect 6049 37678 6059 37734
rect 6115 37678 6125 37734
rect 6049 37592 6125 37678
rect 6049 37536 6059 37592
rect 6115 37536 6125 37592
rect 12406 38160 12624 38170
rect 12406 38104 12416 38160
rect 12472 38104 12558 38160
rect 12614 38104 12624 38160
rect 12406 38018 12624 38104
rect 12406 37962 12416 38018
rect 12472 37962 12558 38018
rect 12614 37962 12624 38018
rect 12406 37876 12624 37962
rect 12406 37820 12416 37876
rect 12472 37820 12558 37876
rect 12614 37820 12624 37876
rect 12406 37734 12624 37820
rect 12406 37678 12416 37734
rect 12472 37678 12558 37734
rect 12614 37678 12624 37734
rect 12406 37592 12624 37678
rect 6049 37450 6125 37536
rect 10425 37570 11495 37580
rect 10425 37514 10435 37570
rect 10491 37514 10577 37570
rect 10633 37514 10719 37570
rect 10775 37514 10861 37570
rect 10917 37514 11003 37570
rect 11059 37514 11145 37570
rect 11201 37514 11287 37570
rect 11343 37514 11429 37570
rect 11485 37514 11495 37570
rect 10425 37504 11495 37514
rect 12406 37536 12416 37592
rect 12472 37536 12558 37592
rect 12614 37536 12624 37592
rect 6049 37394 6059 37450
rect 6115 37394 6125 37450
rect 6049 37308 6125 37394
rect 6049 37252 6059 37308
rect 6115 37252 6125 37308
rect 6049 37166 6125 37252
rect 6049 37110 6059 37166
rect 6115 37110 6125 37166
rect 6049 37024 6125 37110
rect 6049 36968 6059 37024
rect 6115 36968 6125 37024
rect 6049 36882 6125 36968
rect 6049 36826 6059 36882
rect 6115 36826 6125 36882
rect 6049 36816 6125 36826
rect 12406 37450 12624 37536
rect 12406 37394 12416 37450
rect 12472 37394 12558 37450
rect 12614 37394 12624 37450
rect 12406 37308 12624 37394
rect 12406 37252 12416 37308
rect 12472 37252 12558 37308
rect 12614 37252 12624 37308
rect 12406 37166 12624 37252
rect 12406 37110 12416 37166
rect 12472 37110 12558 37166
rect 12614 37110 12624 37166
rect 12406 37024 12624 37110
rect 12406 36968 12416 37024
rect 12472 36968 12558 37024
rect 12614 36968 12624 37024
rect 12406 36882 12624 36968
rect 12406 36826 12416 36882
rect 12472 36826 12558 36882
rect 12614 36826 12624 36882
rect 12406 36816 12624 36826
rect 14942 38160 15018 38170
rect 14942 38104 14952 38160
rect 15008 38104 15018 38160
rect 14942 38018 15018 38104
rect 14942 37962 14952 38018
rect 15008 37962 15018 38018
rect 14942 37876 15018 37962
rect 14942 37820 14952 37876
rect 15008 37820 15018 37876
rect 14942 37734 15018 37820
rect 14942 37678 14952 37734
rect 15008 37678 15018 37734
rect 14942 37592 15018 37678
rect 14942 37536 14952 37592
rect 15008 37536 15018 37592
rect 14942 37450 15018 37536
rect 14942 37394 14952 37450
rect 15008 37394 15018 37450
rect 14942 37308 15018 37394
rect 14942 37252 14952 37308
rect 15008 37252 15018 37308
rect 14942 37166 15018 37252
rect 14942 37110 14952 37166
rect 15008 37110 15018 37166
rect 14942 37024 15018 37110
rect 14942 36968 14952 37024
rect 15008 36968 15018 37024
rect 14942 36882 15018 36968
rect 14942 36826 14952 36882
rect 15008 36826 15018 36882
rect 14942 36816 15018 36826
rect 165 36548 383 36558
rect 165 36492 175 36548
rect 231 36492 317 36548
rect 373 36492 383 36548
rect 165 36406 383 36492
rect 165 36350 175 36406
rect 231 36350 317 36406
rect 373 36350 383 36406
rect 165 36264 383 36350
rect 165 36208 175 36264
rect 231 36208 317 36264
rect 373 36208 383 36264
rect 165 36122 383 36208
rect 165 36066 175 36122
rect 231 36066 317 36122
rect 373 36066 383 36122
rect 165 35980 383 36066
rect 3990 36086 4066 36096
rect 3990 36030 4000 36086
rect 4056 36030 4066 36086
rect 165 35924 175 35980
rect 231 35924 317 35980
rect 373 35924 383 35980
rect 165 35838 383 35924
rect 165 35782 175 35838
rect 231 35782 317 35838
rect 373 35782 383 35838
rect 165 35696 383 35782
rect 165 35640 175 35696
rect 231 35640 317 35696
rect 373 35640 383 35696
rect 165 35554 383 35640
rect 165 35498 175 35554
rect 231 35498 317 35554
rect 373 35498 383 35554
rect 165 35412 383 35498
rect 165 35356 175 35412
rect 231 35356 317 35412
rect 373 35356 383 35412
rect 165 35270 383 35356
rect 165 35214 175 35270
rect 231 35214 317 35270
rect 373 35214 383 35270
rect 165 35128 383 35214
rect 165 35072 175 35128
rect 231 35072 317 35128
rect 373 35072 383 35128
rect 165 34986 383 35072
rect 165 34930 175 34986
rect 231 34930 317 34986
rect 373 34930 383 34986
rect 165 34844 383 34930
rect 165 34788 175 34844
rect 231 34788 317 34844
rect 373 34788 383 34844
rect 165 34702 383 34788
rect 165 34646 175 34702
rect 231 34646 317 34702
rect 373 34646 383 34702
rect 165 34560 383 34646
rect 165 34504 175 34560
rect 231 34504 317 34560
rect 373 34504 383 34560
rect 165 34418 383 34504
rect 165 34362 175 34418
rect 231 34362 317 34418
rect 373 34362 383 34418
rect 165 34276 383 34362
rect 165 34220 175 34276
rect 231 34220 317 34276
rect 373 34220 383 34276
rect 165 34134 383 34220
rect 165 34078 175 34134
rect 231 34078 317 34134
rect 373 34078 383 34134
rect 165 33992 383 34078
rect 486 35987 562 35997
rect 486 35931 496 35987
rect 552 35931 562 35987
rect 486 35845 562 35931
rect 486 35789 496 35845
rect 552 35789 562 35845
rect 486 35703 562 35789
rect 486 35647 496 35703
rect 552 35647 562 35703
rect 486 35561 562 35647
rect 486 35505 496 35561
rect 552 35505 562 35561
rect 486 35419 562 35505
rect 486 35363 496 35419
rect 552 35363 562 35419
rect 486 35277 562 35363
rect 486 35221 496 35277
rect 552 35221 562 35277
rect 486 35135 562 35221
rect 486 35079 496 35135
rect 552 35079 562 35135
rect 486 34993 562 35079
rect 486 34937 496 34993
rect 552 34937 562 34993
rect 486 34851 562 34937
rect 486 34795 496 34851
rect 552 34795 562 34851
rect 486 34709 562 34795
rect 486 34653 496 34709
rect 552 34653 562 34709
rect 486 34567 562 34653
rect 486 34511 496 34567
rect 552 34511 562 34567
rect 486 34425 562 34511
rect 724 35982 800 35992
rect 724 35926 734 35982
rect 790 35926 800 35982
rect 724 35840 800 35926
rect 724 35784 734 35840
rect 790 35784 800 35840
rect 724 35698 800 35784
rect 724 35642 734 35698
rect 790 35642 800 35698
rect 724 35556 800 35642
rect 724 35500 734 35556
rect 790 35500 800 35556
rect 724 35414 800 35500
rect 724 35358 734 35414
rect 790 35358 800 35414
rect 724 35272 800 35358
rect 724 35216 734 35272
rect 790 35216 800 35272
rect 724 35130 800 35216
rect 724 35074 734 35130
rect 790 35074 800 35130
rect 724 34988 800 35074
rect 724 34932 734 34988
rect 790 34932 800 34988
rect 724 34846 800 34932
rect 724 34790 734 34846
rect 790 34790 800 34846
rect 724 34704 800 34790
rect 724 34648 734 34704
rect 790 34648 800 34704
rect 724 34562 800 34648
rect 724 34506 734 34562
rect 790 34506 800 34562
rect 724 34496 800 34506
rect 3092 35982 3168 35992
rect 3092 35926 3102 35982
rect 3158 35926 3168 35982
rect 3092 35840 3168 35926
rect 3092 35784 3102 35840
rect 3158 35784 3168 35840
rect 3092 35698 3168 35784
rect 3092 35642 3102 35698
rect 3158 35642 3168 35698
rect 3092 35556 3168 35642
rect 3092 35500 3102 35556
rect 3158 35500 3168 35556
rect 3092 35414 3168 35500
rect 3092 35358 3102 35414
rect 3158 35358 3168 35414
rect 3092 35272 3168 35358
rect 3092 35216 3102 35272
rect 3158 35216 3168 35272
rect 3092 35130 3168 35216
rect 3092 35074 3102 35130
rect 3158 35074 3168 35130
rect 3092 34988 3168 35074
rect 3092 34932 3102 34988
rect 3158 34932 3168 34988
rect 3092 34846 3168 34932
rect 3092 34790 3102 34846
rect 3158 34790 3168 34846
rect 3092 34704 3168 34790
rect 3092 34648 3102 34704
rect 3158 34648 3168 34704
rect 3092 34562 3168 34648
rect 3092 34506 3102 34562
rect 3158 34506 3168 34562
rect 3092 34496 3168 34506
rect 3990 35944 4066 36030
rect 10998 36086 11074 36096
rect 10998 36030 11008 36086
rect 11064 36030 11074 36086
rect 3990 35888 4000 35944
rect 4056 35888 4066 35944
rect 3990 35802 4066 35888
rect 3990 35746 4000 35802
rect 4056 35746 4066 35802
rect 3990 35660 4066 35746
rect 3990 35604 4000 35660
rect 4056 35604 4066 35660
rect 3990 35518 4066 35604
rect 3990 35462 4000 35518
rect 4056 35462 4066 35518
rect 3990 35376 4066 35462
rect 3990 35320 4000 35376
rect 4056 35320 4066 35376
rect 3990 35234 4066 35320
rect 3990 35178 4000 35234
rect 4056 35178 4066 35234
rect 3990 35092 4066 35178
rect 3990 35036 4000 35092
rect 4056 35036 4066 35092
rect 3990 34950 4066 35036
rect 3990 34894 4000 34950
rect 4056 34894 4066 34950
rect 3990 34808 4066 34894
rect 3990 34752 4000 34808
rect 4056 34752 4066 34808
rect 3990 34666 4066 34752
rect 3990 34610 4000 34666
rect 4056 34610 4066 34666
rect 3990 34524 4066 34610
rect 486 34369 496 34425
rect 552 34369 562 34425
rect 486 34283 562 34369
rect 486 34227 496 34283
rect 552 34227 562 34283
rect 486 34141 562 34227
rect 486 34085 496 34141
rect 552 34085 562 34141
rect 486 34075 562 34085
rect 3990 34468 4000 34524
rect 4056 34468 4066 34524
rect 4888 35982 4964 35992
rect 4888 35926 4898 35982
rect 4954 35926 4964 35982
rect 4888 35840 4964 35926
rect 4888 35784 4898 35840
rect 4954 35784 4964 35840
rect 4888 35698 4964 35784
rect 4888 35642 4898 35698
rect 4954 35642 4964 35698
rect 4888 35556 4964 35642
rect 4888 35500 4898 35556
rect 4954 35500 4964 35556
rect 4888 35414 4964 35500
rect 4888 35358 4898 35414
rect 4954 35358 4964 35414
rect 4888 35272 4964 35358
rect 4888 35216 4898 35272
rect 4954 35216 4964 35272
rect 4888 35130 4964 35216
rect 4888 35074 4898 35130
rect 4954 35074 4964 35130
rect 4888 34988 4964 35074
rect 4888 34932 4898 34988
rect 4954 34932 4964 34988
rect 4888 34846 4964 34932
rect 4888 34790 4898 34846
rect 4954 34790 4964 34846
rect 4888 34704 4964 34790
rect 4888 34648 4898 34704
rect 4954 34648 4964 34704
rect 4888 34562 4964 34648
rect 4888 34506 4898 34562
rect 4954 34506 4964 34562
rect 4888 34496 4964 34506
rect 8671 35982 8747 35992
rect 8671 35926 8681 35982
rect 8737 35926 8747 35982
rect 8671 35840 8747 35926
rect 8671 35784 8681 35840
rect 8737 35784 8747 35840
rect 8671 35698 8747 35784
rect 8671 35642 8681 35698
rect 8737 35642 8747 35698
rect 8671 35556 8747 35642
rect 8671 35500 8681 35556
rect 8737 35500 8747 35556
rect 8671 35414 8747 35500
rect 8671 35358 8681 35414
rect 8737 35358 8747 35414
rect 8671 35272 8747 35358
rect 8671 35216 8681 35272
rect 8737 35216 8747 35272
rect 8671 35130 8747 35216
rect 8671 35074 8681 35130
rect 8737 35074 8747 35130
rect 8671 34988 8747 35074
rect 8671 34932 8681 34988
rect 8737 34932 8747 34988
rect 8671 34846 8747 34932
rect 8671 34790 8681 34846
rect 8737 34790 8747 34846
rect 8671 34704 8747 34790
rect 8671 34648 8681 34704
rect 8737 34648 8747 34704
rect 8671 34562 8747 34648
rect 8671 34506 8681 34562
rect 8737 34506 8747 34562
rect 8671 34496 8747 34506
rect 10100 35982 10176 35992
rect 10100 35926 10110 35982
rect 10166 35926 10176 35982
rect 10100 35840 10176 35926
rect 10100 35784 10110 35840
rect 10166 35784 10176 35840
rect 10100 35698 10176 35784
rect 10100 35642 10110 35698
rect 10166 35642 10176 35698
rect 10100 35556 10176 35642
rect 10100 35500 10110 35556
rect 10166 35500 10176 35556
rect 10100 35414 10176 35500
rect 10100 35358 10110 35414
rect 10166 35358 10176 35414
rect 10100 35272 10176 35358
rect 10100 35216 10110 35272
rect 10166 35216 10176 35272
rect 10100 35130 10176 35216
rect 10100 35074 10110 35130
rect 10166 35074 10176 35130
rect 10100 34988 10176 35074
rect 10100 34932 10110 34988
rect 10166 34932 10176 34988
rect 10100 34846 10176 34932
rect 10100 34790 10110 34846
rect 10166 34790 10176 34846
rect 10100 34704 10176 34790
rect 10100 34648 10110 34704
rect 10166 34648 10176 34704
rect 10100 34562 10176 34648
rect 10100 34506 10110 34562
rect 10166 34506 10176 34562
rect 10100 34496 10176 34506
rect 10998 35944 11074 36030
rect 10998 35888 11008 35944
rect 11064 35888 11074 35944
rect 10998 35802 11074 35888
rect 10998 35746 11008 35802
rect 11064 35746 11074 35802
rect 10998 35660 11074 35746
rect 10998 35604 11008 35660
rect 11064 35604 11074 35660
rect 10998 35518 11074 35604
rect 10998 35462 11008 35518
rect 11064 35462 11074 35518
rect 10998 35376 11074 35462
rect 10998 35320 11008 35376
rect 11064 35320 11074 35376
rect 10998 35234 11074 35320
rect 10998 35178 11008 35234
rect 11064 35178 11074 35234
rect 10998 35092 11074 35178
rect 10998 35036 11008 35092
rect 11064 35036 11074 35092
rect 10998 34950 11074 35036
rect 10998 34894 11008 34950
rect 11064 34894 11074 34950
rect 10998 34808 11074 34894
rect 10998 34752 11008 34808
rect 11064 34752 11074 34808
rect 10998 34666 11074 34752
rect 10998 34610 11008 34666
rect 11064 34610 11074 34666
rect 10998 34524 11074 34610
rect 3990 34382 4066 34468
rect 3990 34326 4000 34382
rect 4056 34326 4066 34382
rect 3990 34240 4066 34326
rect 3990 34184 4000 34240
rect 4056 34184 4066 34240
rect 3990 34098 4066 34184
rect 165 33936 175 33992
rect 231 33936 317 33992
rect 373 33936 383 33992
rect 165 33850 383 33936
rect 165 33794 175 33850
rect 231 33794 317 33850
rect 373 33794 383 33850
rect 165 33708 383 33794
rect 165 33652 175 33708
rect 231 33652 317 33708
rect 373 33652 383 33708
rect 165 33642 383 33652
rect 3990 34042 4000 34098
rect 4056 34042 4066 34098
rect 3990 33956 4066 34042
rect 3990 33900 4000 33956
rect 4056 33900 4066 33956
rect 3990 33814 4066 33900
rect 3990 33758 4000 33814
rect 4056 33758 4066 33814
rect 3990 33672 4066 33758
rect 3990 33616 4000 33672
rect 4056 33616 4066 33672
rect 3990 33606 4066 33616
rect 10998 34468 11008 34524
rect 11064 34468 11074 34524
rect 11896 35982 11972 35992
rect 11896 35926 11906 35982
rect 11962 35926 11972 35982
rect 11896 35840 11972 35926
rect 11896 35784 11906 35840
rect 11962 35784 11972 35840
rect 11896 35698 11972 35784
rect 11896 35642 11906 35698
rect 11962 35642 11972 35698
rect 11896 35556 11972 35642
rect 11896 35500 11906 35556
rect 11962 35500 11972 35556
rect 11896 35414 11972 35500
rect 11896 35358 11906 35414
rect 11962 35358 11972 35414
rect 11896 35272 11972 35358
rect 11896 35216 11906 35272
rect 11962 35216 11972 35272
rect 11896 35130 11972 35216
rect 11896 35074 11906 35130
rect 11962 35074 11972 35130
rect 11896 34988 11972 35074
rect 11896 34932 11906 34988
rect 11962 34932 11972 34988
rect 11896 34846 11972 34932
rect 11896 34790 11906 34846
rect 11962 34790 11972 34846
rect 11896 34704 11972 34790
rect 11896 34648 11906 34704
rect 11962 34648 11972 34704
rect 11896 34562 11972 34648
rect 11896 34506 11906 34562
rect 11962 34506 11972 34562
rect 11896 34496 11972 34506
rect 10998 34382 11074 34468
rect 10998 34326 11008 34382
rect 11064 34326 11074 34382
rect 10998 34240 11074 34326
rect 10998 34184 11008 34240
rect 11064 34184 11074 34240
rect 10998 34098 11074 34184
rect 10998 34042 11008 34098
rect 11064 34042 11074 34098
rect 10998 33956 11074 34042
rect 10998 33900 11008 33956
rect 11064 33900 11074 33956
rect 10998 33814 11074 33900
rect 10998 33758 11008 33814
rect 11064 33758 11074 33814
rect 10998 33672 11074 33758
rect 10998 33616 11008 33672
rect 11064 33616 11074 33672
rect 10998 33606 11074 33616
rect 486 33348 562 33358
rect 486 33292 496 33348
rect 552 33292 562 33348
rect 486 33206 562 33292
rect 486 33150 496 33206
rect 552 33150 562 33206
rect 486 33064 562 33150
rect 486 33008 496 33064
rect 552 33008 562 33064
rect 486 32922 562 33008
rect 486 32866 496 32922
rect 552 32866 562 32922
rect 14400 33348 14760 33358
rect 14400 33292 14410 33348
rect 14466 33292 14552 33348
rect 14608 33292 14694 33348
rect 14750 33292 14760 33348
rect 14400 33206 14760 33292
rect 14400 33150 14410 33206
rect 14466 33150 14552 33206
rect 14608 33150 14694 33206
rect 14750 33150 14760 33206
rect 14400 33064 14760 33150
rect 14400 33008 14410 33064
rect 14466 33008 14552 33064
rect 14608 33008 14694 33064
rect 14750 33008 14760 33064
rect 14400 32922 14760 33008
rect 486 32780 562 32866
rect 486 32724 496 32780
rect 552 32724 562 32780
rect 486 32638 562 32724
rect 3990 32905 4066 32915
rect 3990 32849 4000 32905
rect 4056 32849 4066 32905
rect 3990 32763 4066 32849
rect 3990 32707 4000 32763
rect 4056 32707 4066 32763
rect 486 32582 496 32638
rect 552 32582 562 32638
rect 486 32496 562 32582
rect 486 32440 496 32496
rect 552 32440 562 32496
rect 486 32354 562 32440
rect 486 32298 496 32354
rect 552 32298 562 32354
rect 486 32212 562 32298
rect 486 32156 496 32212
rect 552 32156 562 32212
rect 486 32070 562 32156
rect 486 32014 496 32070
rect 552 32014 562 32070
rect 486 31928 562 32014
rect 486 31872 496 31928
rect 552 31872 562 31928
rect 486 31786 562 31872
rect 486 31730 496 31786
rect 552 31730 562 31786
rect 486 31644 562 31730
rect 486 31588 496 31644
rect 552 31588 562 31644
rect 486 31502 562 31588
rect 486 31446 496 31502
rect 552 31446 562 31502
rect 486 31360 562 31446
rect 486 31304 496 31360
rect 552 31304 562 31360
rect 486 31218 562 31304
rect 486 31162 496 31218
rect 552 31162 562 31218
rect 486 31076 562 31162
rect 486 31020 496 31076
rect 552 31020 562 31076
rect 486 30934 562 31020
rect 486 30878 496 30934
rect 552 30878 562 30934
rect 486 30792 562 30878
rect 486 30736 496 30792
rect 552 30736 562 30792
rect 486 30650 562 30736
rect 486 30594 496 30650
rect 552 30594 562 30650
rect 486 30508 562 30594
rect 486 30452 496 30508
rect 552 30452 562 30508
rect 968 32692 1044 32702
rect 968 32636 978 32692
rect 1034 32636 1044 32692
rect 968 32550 1044 32636
rect 968 32494 978 32550
rect 1034 32494 1044 32550
rect 968 32408 1044 32494
rect 968 32352 978 32408
rect 1034 32352 1044 32408
rect 968 32266 1044 32352
rect 968 32210 978 32266
rect 1034 32210 1044 32266
rect 968 32124 1044 32210
rect 968 32068 978 32124
rect 1034 32068 1044 32124
rect 968 31982 1044 32068
rect 968 31926 978 31982
rect 1034 31926 1044 31982
rect 968 31840 1044 31926
rect 968 31784 978 31840
rect 1034 31784 1044 31840
rect 968 31698 1044 31784
rect 968 31642 978 31698
rect 1034 31642 1044 31698
rect 968 31556 1044 31642
rect 968 31500 978 31556
rect 1034 31500 1044 31556
rect 968 31414 1044 31500
rect 968 31358 978 31414
rect 1034 31358 1044 31414
rect 968 31272 1044 31358
rect 968 31216 978 31272
rect 1034 31216 1044 31272
rect 968 31130 1044 31216
rect 968 31074 978 31130
rect 1034 31074 1044 31130
rect 968 30988 1044 31074
rect 968 30932 978 30988
rect 1034 30932 1044 30988
rect 968 30846 1044 30932
rect 968 30790 978 30846
rect 1034 30790 1044 30846
rect 968 30704 1044 30790
rect 968 30648 978 30704
rect 1034 30648 1044 30704
rect 968 30562 1044 30648
rect 968 30506 978 30562
rect 1034 30506 1044 30562
rect 968 30496 1044 30506
rect 2360 32692 2436 32702
rect 2360 32636 2370 32692
rect 2426 32636 2436 32692
rect 2360 32550 2436 32636
rect 2360 32494 2370 32550
rect 2426 32494 2436 32550
rect 2360 32408 2436 32494
rect 2360 32352 2370 32408
rect 2426 32352 2436 32408
rect 2360 32266 2436 32352
rect 2360 32210 2370 32266
rect 2426 32210 2436 32266
rect 2360 32124 2436 32210
rect 2360 32068 2370 32124
rect 2426 32068 2436 32124
rect 2360 31982 2436 32068
rect 2360 31926 2370 31982
rect 2426 31926 2436 31982
rect 2360 31840 2436 31926
rect 2360 31784 2370 31840
rect 2426 31784 2436 31840
rect 2360 31698 2436 31784
rect 2360 31642 2370 31698
rect 2426 31642 2436 31698
rect 2360 31556 2436 31642
rect 2360 31500 2370 31556
rect 2426 31500 2436 31556
rect 2360 31414 2436 31500
rect 2360 31358 2370 31414
rect 2426 31358 2436 31414
rect 2360 31272 2436 31358
rect 2360 31216 2370 31272
rect 2426 31216 2436 31272
rect 2360 31130 2436 31216
rect 2360 31074 2370 31130
rect 2426 31074 2436 31130
rect 2360 30988 2436 31074
rect 2360 30932 2370 30988
rect 2426 30932 2436 30988
rect 2360 30846 2436 30932
rect 2360 30790 2370 30846
rect 2426 30790 2436 30846
rect 2360 30704 2436 30790
rect 2360 30648 2370 30704
rect 2426 30648 2436 30704
rect 2360 30562 2436 30648
rect 2360 30506 2370 30562
rect 2426 30506 2436 30562
rect 2360 30496 2436 30506
rect 2776 32692 2852 32702
rect 2776 32636 2786 32692
rect 2842 32636 2852 32692
rect 2776 32550 2852 32636
rect 2776 32494 2786 32550
rect 2842 32494 2852 32550
rect 2776 32408 2852 32494
rect 2776 32352 2786 32408
rect 2842 32352 2852 32408
rect 2776 32266 2852 32352
rect 2776 32210 2786 32266
rect 2842 32210 2852 32266
rect 2776 32124 2852 32210
rect 2776 32068 2786 32124
rect 2842 32068 2852 32124
rect 2776 31982 2852 32068
rect 2776 31926 2786 31982
rect 2842 31926 2852 31982
rect 2776 31840 2852 31926
rect 2776 31784 2786 31840
rect 2842 31784 2852 31840
rect 2776 31698 2852 31784
rect 2776 31642 2786 31698
rect 2842 31642 2852 31698
rect 2776 31556 2852 31642
rect 2776 31500 2786 31556
rect 2842 31500 2852 31556
rect 2776 31414 2852 31500
rect 2776 31358 2786 31414
rect 2842 31358 2852 31414
rect 2776 31272 2852 31358
rect 2776 31216 2786 31272
rect 2842 31216 2852 31272
rect 2776 31130 2852 31216
rect 2776 31074 2786 31130
rect 2842 31074 2852 31130
rect 2776 30988 2852 31074
rect 3264 32693 3340 32703
rect 3264 32637 3274 32693
rect 3330 32637 3340 32693
rect 3264 32551 3340 32637
rect 3264 32495 3274 32551
rect 3330 32495 3340 32551
rect 3264 32409 3340 32495
rect 3264 32353 3274 32409
rect 3330 32353 3340 32409
rect 3264 32267 3340 32353
rect 3264 32211 3274 32267
rect 3330 32211 3340 32267
rect 3264 32125 3340 32211
rect 3264 32069 3274 32125
rect 3330 32069 3340 32125
rect 3264 31983 3340 32069
rect 3264 31927 3274 31983
rect 3330 31927 3340 31983
rect 3264 31841 3340 31927
rect 3264 31785 3274 31841
rect 3330 31785 3340 31841
rect 3264 31699 3340 31785
rect 3264 31643 3274 31699
rect 3330 31643 3340 31699
rect 3264 31557 3340 31643
rect 3264 31501 3274 31557
rect 3330 31501 3340 31557
rect 3264 31415 3340 31501
rect 3264 31359 3274 31415
rect 3330 31359 3340 31415
rect 3264 31273 3340 31359
rect 3264 31217 3274 31273
rect 3330 31217 3340 31273
rect 3264 31131 3340 31217
rect 3264 31075 3274 31131
rect 3330 31075 3340 31131
rect 3264 31065 3340 31075
rect 3752 32642 3828 32652
rect 3752 32586 3762 32642
rect 3818 32586 3828 32642
rect 3752 32500 3828 32586
rect 3752 32444 3762 32500
rect 3818 32444 3828 32500
rect 3752 32358 3828 32444
rect 3752 32302 3762 32358
rect 3818 32302 3828 32358
rect 3752 32216 3828 32302
rect 3752 32160 3762 32216
rect 3818 32160 3828 32216
rect 3752 32074 3828 32160
rect 3752 32018 3762 32074
rect 3818 32018 3828 32074
rect 3752 31932 3828 32018
rect 3752 31876 3762 31932
rect 3818 31876 3828 31932
rect 3752 31790 3828 31876
rect 3752 31734 3762 31790
rect 3818 31734 3828 31790
rect 3752 31648 3828 31734
rect 3752 31592 3762 31648
rect 3818 31592 3828 31648
rect 3752 31506 3828 31592
rect 3752 31450 3762 31506
rect 3818 31450 3828 31506
rect 3752 31364 3828 31450
rect 3752 31308 3762 31364
rect 3818 31308 3828 31364
rect 3752 31222 3828 31308
rect 3752 31166 3762 31222
rect 3818 31166 3828 31222
rect 3752 31080 3828 31166
rect 3752 31024 3762 31080
rect 3818 31024 3828 31080
rect 3752 31014 3828 31024
rect 3990 32621 4066 32707
rect 10998 32905 11074 32915
rect 10998 32849 11008 32905
rect 11064 32849 11074 32905
rect 10998 32763 11074 32849
rect 10998 32707 11008 32763
rect 11064 32707 11074 32763
rect 4716 32693 4792 32703
rect 3990 32565 4000 32621
rect 4056 32565 4066 32621
rect 3990 32479 4066 32565
rect 3990 32423 4000 32479
rect 4056 32423 4066 32479
rect 3990 32337 4066 32423
rect 3990 32281 4000 32337
rect 4056 32281 4066 32337
rect 3990 32195 4066 32281
rect 3990 32139 4000 32195
rect 4056 32139 4066 32195
rect 3990 32053 4066 32139
rect 3990 31997 4000 32053
rect 4056 31997 4066 32053
rect 3990 31911 4066 31997
rect 3990 31855 4000 31911
rect 4056 31855 4066 31911
rect 3990 31769 4066 31855
rect 3990 31713 4000 31769
rect 4056 31713 4066 31769
rect 3990 31627 4066 31713
rect 3990 31571 4000 31627
rect 4056 31571 4066 31627
rect 3990 31485 4066 31571
rect 3990 31429 4000 31485
rect 4056 31429 4066 31485
rect 3990 31343 4066 31429
rect 3990 31287 4000 31343
rect 4056 31287 4066 31343
rect 3990 31201 4066 31287
rect 3990 31145 4000 31201
rect 4056 31145 4066 31201
rect 3990 31059 4066 31145
rect 3990 31003 4000 31059
rect 4056 31003 4066 31059
rect 4228 32642 4304 32652
rect 4228 32586 4238 32642
rect 4294 32586 4304 32642
rect 4228 32500 4304 32586
rect 4228 32444 4238 32500
rect 4294 32444 4304 32500
rect 4228 32358 4304 32444
rect 4228 32302 4238 32358
rect 4294 32302 4304 32358
rect 4228 32216 4304 32302
rect 4228 32160 4238 32216
rect 4294 32160 4304 32216
rect 4228 32074 4304 32160
rect 4228 32018 4238 32074
rect 4294 32018 4304 32074
rect 4228 31932 4304 32018
rect 4228 31876 4238 31932
rect 4294 31876 4304 31932
rect 4228 31790 4304 31876
rect 4228 31734 4238 31790
rect 4294 31734 4304 31790
rect 4228 31648 4304 31734
rect 4228 31592 4238 31648
rect 4294 31592 4304 31648
rect 4228 31506 4304 31592
rect 4228 31450 4238 31506
rect 4294 31450 4304 31506
rect 4228 31364 4304 31450
rect 4228 31308 4238 31364
rect 4294 31308 4304 31364
rect 4228 31222 4304 31308
rect 4228 31166 4238 31222
rect 4294 31166 4304 31222
rect 4228 31080 4304 31166
rect 4228 31024 4238 31080
rect 4294 31024 4304 31080
rect 4716 32637 4726 32693
rect 4782 32637 4792 32693
rect 4716 32551 4792 32637
rect 4716 32495 4726 32551
rect 4782 32495 4792 32551
rect 4716 32409 4792 32495
rect 4716 32353 4726 32409
rect 4782 32353 4792 32409
rect 4716 32267 4792 32353
rect 4716 32211 4726 32267
rect 4782 32211 4792 32267
rect 4716 32125 4792 32211
rect 4716 32069 4726 32125
rect 4782 32069 4792 32125
rect 4716 31983 4792 32069
rect 4716 31927 4726 31983
rect 4782 31927 4792 31983
rect 4716 31841 4792 31927
rect 4716 31785 4726 31841
rect 4782 31785 4792 31841
rect 4716 31699 4792 31785
rect 4716 31643 4726 31699
rect 4782 31643 4792 31699
rect 4716 31557 4792 31643
rect 4716 31501 4726 31557
rect 4782 31501 4792 31557
rect 4716 31415 4792 31501
rect 4716 31359 4726 31415
rect 4782 31359 4792 31415
rect 4716 31273 4792 31359
rect 4716 31217 4726 31273
rect 4782 31217 4792 31273
rect 4716 31131 4792 31217
rect 4716 31075 4726 31131
rect 4782 31075 4792 31131
rect 4716 31065 4792 31075
rect 5204 32693 5280 32703
rect 5204 32637 5214 32693
rect 5270 32637 5280 32693
rect 5204 32551 5280 32637
rect 5204 32495 5214 32551
rect 5270 32495 5280 32551
rect 5204 32409 5280 32495
rect 5204 32353 5214 32409
rect 5270 32353 5280 32409
rect 5204 32267 5280 32353
rect 5204 32211 5214 32267
rect 5270 32211 5280 32267
rect 5204 32125 5280 32211
rect 5204 32069 5214 32125
rect 5270 32069 5280 32125
rect 5204 31983 5280 32069
rect 5204 31927 5214 31983
rect 5270 31927 5280 31983
rect 5204 31841 5280 31927
rect 5204 31785 5214 31841
rect 5270 31785 5280 31841
rect 5204 31699 5280 31785
rect 5204 31643 5214 31699
rect 5270 31643 5280 31699
rect 5204 31557 5280 31643
rect 5204 31501 5214 31557
rect 5270 31501 5280 31557
rect 5204 31415 5280 31501
rect 5204 31359 5214 31415
rect 5270 31359 5280 31415
rect 5204 31273 5280 31359
rect 5204 31217 5214 31273
rect 5270 31217 5280 31273
rect 5204 31131 5280 31217
rect 5204 31075 5214 31131
rect 5270 31075 5280 31131
rect 5204 31065 5280 31075
rect 5620 32693 5696 32703
rect 5620 32637 5630 32693
rect 5686 32637 5696 32693
rect 5620 32551 5696 32637
rect 5620 32495 5630 32551
rect 5686 32495 5696 32551
rect 5620 32409 5696 32495
rect 5620 32353 5630 32409
rect 5686 32353 5696 32409
rect 5620 32267 5696 32353
rect 5620 32211 5630 32267
rect 5686 32211 5696 32267
rect 5620 32125 5696 32211
rect 5620 32069 5630 32125
rect 5686 32069 5696 32125
rect 5620 31983 5696 32069
rect 5620 31927 5630 31983
rect 5686 31927 5696 31983
rect 5620 31841 5696 31927
rect 5620 31785 5630 31841
rect 5686 31785 5696 31841
rect 5620 31699 5696 31785
rect 5620 31643 5630 31699
rect 5686 31643 5696 31699
rect 5620 31557 5696 31643
rect 5620 31501 5630 31557
rect 5686 31501 5696 31557
rect 5620 31415 5696 31501
rect 5620 31359 5630 31415
rect 5686 31359 5696 31415
rect 5620 31273 5696 31359
rect 5620 31217 5630 31273
rect 5686 31217 5696 31273
rect 5620 31131 5696 31217
rect 5620 31075 5630 31131
rect 5686 31075 5696 31131
rect 5620 31065 5696 31075
rect 7012 32692 7088 32702
rect 7012 32636 7022 32692
rect 7078 32636 7088 32692
rect 7012 32550 7088 32636
rect 7012 32494 7022 32550
rect 7078 32494 7088 32550
rect 7012 32408 7088 32494
rect 7012 32352 7022 32408
rect 7078 32352 7088 32408
rect 7012 32266 7088 32352
rect 7012 32210 7022 32266
rect 7078 32210 7088 32266
rect 7012 32124 7088 32210
rect 7012 32068 7022 32124
rect 7078 32068 7088 32124
rect 7012 31982 7088 32068
rect 7012 31926 7022 31982
rect 7078 31926 7088 31982
rect 7012 31840 7088 31926
rect 7012 31784 7022 31840
rect 7078 31784 7088 31840
rect 7012 31698 7088 31784
rect 7012 31642 7022 31698
rect 7078 31642 7088 31698
rect 7012 31556 7088 31642
rect 7012 31500 7022 31556
rect 7078 31500 7088 31556
rect 7012 31414 7088 31500
rect 7012 31358 7022 31414
rect 7078 31358 7088 31414
rect 7012 31272 7088 31358
rect 7012 31216 7022 31272
rect 7078 31216 7088 31272
rect 7012 31130 7088 31216
rect 7012 31074 7022 31130
rect 7078 31074 7088 31130
rect 4228 31014 4304 31024
rect 3990 30993 4066 31003
rect 2776 30932 2786 30988
rect 2842 30932 2852 30988
rect 2776 30846 2852 30932
rect 2776 30790 2786 30846
rect 2842 30790 2852 30846
rect 2776 30704 2852 30790
rect 2776 30648 2786 30704
rect 2842 30648 2852 30704
rect 2776 30562 2852 30648
rect 2776 30506 2786 30562
rect 2842 30506 2852 30562
rect 2776 30496 2852 30506
rect 7012 30988 7088 31074
rect 7012 30932 7022 30988
rect 7078 30932 7088 30988
rect 7012 30846 7088 30932
rect 7012 30790 7022 30846
rect 7078 30790 7088 30846
rect 7012 30704 7088 30790
rect 7012 30648 7022 30704
rect 7078 30648 7088 30704
rect 7012 30562 7088 30648
rect 7012 30506 7022 30562
rect 7078 30506 7088 30562
rect 7012 30496 7088 30506
rect 7976 32692 8052 32702
rect 7976 32636 7986 32692
rect 8042 32636 8052 32692
rect 7976 32550 8052 32636
rect 7976 32494 7986 32550
rect 8042 32494 8052 32550
rect 7976 32408 8052 32494
rect 7976 32352 7986 32408
rect 8042 32352 8052 32408
rect 7976 32266 8052 32352
rect 7976 32210 7986 32266
rect 8042 32210 8052 32266
rect 7976 32124 8052 32210
rect 7976 32068 7986 32124
rect 8042 32068 8052 32124
rect 7976 31982 8052 32068
rect 7976 31926 7986 31982
rect 8042 31926 8052 31982
rect 7976 31840 8052 31926
rect 7976 31784 7986 31840
rect 8042 31784 8052 31840
rect 7976 31698 8052 31784
rect 7976 31642 7986 31698
rect 8042 31642 8052 31698
rect 7976 31556 8052 31642
rect 7976 31500 7986 31556
rect 8042 31500 8052 31556
rect 7976 31414 8052 31500
rect 7976 31358 7986 31414
rect 8042 31358 8052 31414
rect 7976 31272 8052 31358
rect 7976 31216 7986 31272
rect 8042 31216 8052 31272
rect 7976 31130 8052 31216
rect 7976 31074 7986 31130
rect 8042 31074 8052 31130
rect 7976 30988 8052 31074
rect 9368 32693 9444 32703
rect 9368 32637 9378 32693
rect 9434 32637 9444 32693
rect 9368 32551 9444 32637
rect 9368 32495 9378 32551
rect 9434 32495 9444 32551
rect 9368 32409 9444 32495
rect 9368 32353 9378 32409
rect 9434 32353 9444 32409
rect 9368 32267 9444 32353
rect 9368 32211 9378 32267
rect 9434 32211 9444 32267
rect 9368 32125 9444 32211
rect 9368 32069 9378 32125
rect 9434 32069 9444 32125
rect 9368 31983 9444 32069
rect 9368 31927 9378 31983
rect 9434 31927 9444 31983
rect 9368 31841 9444 31927
rect 9368 31785 9378 31841
rect 9434 31785 9444 31841
rect 9368 31699 9444 31785
rect 9368 31643 9378 31699
rect 9434 31643 9444 31699
rect 9368 31557 9444 31643
rect 9368 31501 9378 31557
rect 9434 31501 9444 31557
rect 9368 31415 9444 31501
rect 9368 31359 9378 31415
rect 9434 31359 9444 31415
rect 9368 31273 9444 31359
rect 9368 31217 9378 31273
rect 9434 31217 9444 31273
rect 9368 31131 9444 31217
rect 9368 31075 9378 31131
rect 9434 31075 9444 31131
rect 9368 31065 9444 31075
rect 9784 32693 9860 32703
rect 9784 32637 9794 32693
rect 9850 32637 9860 32693
rect 9784 32551 9860 32637
rect 9784 32495 9794 32551
rect 9850 32495 9860 32551
rect 9784 32409 9860 32495
rect 9784 32353 9794 32409
rect 9850 32353 9860 32409
rect 9784 32267 9860 32353
rect 9784 32211 9794 32267
rect 9850 32211 9860 32267
rect 9784 32125 9860 32211
rect 9784 32069 9794 32125
rect 9850 32069 9860 32125
rect 9784 31983 9860 32069
rect 9784 31927 9794 31983
rect 9850 31927 9860 31983
rect 9784 31841 9860 31927
rect 9784 31785 9794 31841
rect 9850 31785 9860 31841
rect 9784 31699 9860 31785
rect 9784 31643 9794 31699
rect 9850 31643 9860 31699
rect 9784 31557 9860 31643
rect 9784 31501 9794 31557
rect 9850 31501 9860 31557
rect 9784 31415 9860 31501
rect 9784 31359 9794 31415
rect 9850 31359 9860 31415
rect 9784 31273 9860 31359
rect 9784 31217 9794 31273
rect 9850 31217 9860 31273
rect 9784 31131 9860 31217
rect 9784 31075 9794 31131
rect 9850 31075 9860 31131
rect 9784 31065 9860 31075
rect 10272 32693 10348 32703
rect 10272 32637 10282 32693
rect 10338 32637 10348 32693
rect 10272 32551 10348 32637
rect 10272 32495 10282 32551
rect 10338 32495 10348 32551
rect 10272 32409 10348 32495
rect 10272 32353 10282 32409
rect 10338 32353 10348 32409
rect 10272 32267 10348 32353
rect 10272 32211 10282 32267
rect 10338 32211 10348 32267
rect 10272 32125 10348 32211
rect 10272 32069 10282 32125
rect 10338 32069 10348 32125
rect 10272 31983 10348 32069
rect 10272 31927 10282 31983
rect 10338 31927 10348 31983
rect 10272 31841 10348 31927
rect 10272 31785 10282 31841
rect 10338 31785 10348 31841
rect 10272 31699 10348 31785
rect 10272 31643 10282 31699
rect 10338 31643 10348 31699
rect 10272 31557 10348 31643
rect 10272 31501 10282 31557
rect 10338 31501 10348 31557
rect 10272 31415 10348 31501
rect 10272 31359 10282 31415
rect 10338 31359 10348 31415
rect 10272 31273 10348 31359
rect 10272 31217 10282 31273
rect 10338 31217 10348 31273
rect 10272 31131 10348 31217
rect 10272 31075 10282 31131
rect 10338 31075 10348 31131
rect 10272 31065 10348 31075
rect 10760 32642 10836 32652
rect 10760 32586 10770 32642
rect 10826 32586 10836 32642
rect 10760 32500 10836 32586
rect 10760 32444 10770 32500
rect 10826 32444 10836 32500
rect 10760 32358 10836 32444
rect 10760 32302 10770 32358
rect 10826 32302 10836 32358
rect 10760 32216 10836 32302
rect 10760 32160 10770 32216
rect 10826 32160 10836 32216
rect 10760 32074 10836 32160
rect 10760 32018 10770 32074
rect 10826 32018 10836 32074
rect 10760 31932 10836 32018
rect 10760 31876 10770 31932
rect 10826 31876 10836 31932
rect 10760 31790 10836 31876
rect 10760 31734 10770 31790
rect 10826 31734 10836 31790
rect 10760 31648 10836 31734
rect 10760 31592 10770 31648
rect 10826 31592 10836 31648
rect 10760 31506 10836 31592
rect 10760 31450 10770 31506
rect 10826 31450 10836 31506
rect 10760 31364 10836 31450
rect 10760 31308 10770 31364
rect 10826 31308 10836 31364
rect 10760 31222 10836 31308
rect 10760 31166 10770 31222
rect 10826 31166 10836 31222
rect 10760 31080 10836 31166
rect 10760 31024 10770 31080
rect 10826 31024 10836 31080
rect 10760 31014 10836 31024
rect 10998 32621 11074 32707
rect 14400 32866 14410 32922
rect 14466 32866 14552 32922
rect 14608 32866 14694 32922
rect 14750 32866 14760 32922
rect 14400 32780 14760 32866
rect 14400 32724 14410 32780
rect 14466 32724 14552 32780
rect 14608 32724 14694 32780
rect 14750 32724 14760 32780
rect 11724 32693 11800 32703
rect 10998 32565 11008 32621
rect 11064 32565 11074 32621
rect 10998 32479 11074 32565
rect 10998 32423 11008 32479
rect 11064 32423 11074 32479
rect 10998 32337 11074 32423
rect 10998 32281 11008 32337
rect 11064 32281 11074 32337
rect 10998 32195 11074 32281
rect 10998 32139 11008 32195
rect 11064 32139 11074 32195
rect 10998 32053 11074 32139
rect 10998 31997 11008 32053
rect 11064 31997 11074 32053
rect 10998 31911 11074 31997
rect 10998 31855 11008 31911
rect 11064 31855 11074 31911
rect 10998 31769 11074 31855
rect 10998 31713 11008 31769
rect 11064 31713 11074 31769
rect 10998 31627 11074 31713
rect 10998 31571 11008 31627
rect 11064 31571 11074 31627
rect 10998 31485 11074 31571
rect 10998 31429 11008 31485
rect 11064 31429 11074 31485
rect 10998 31343 11074 31429
rect 10998 31287 11008 31343
rect 11064 31287 11074 31343
rect 10998 31201 11074 31287
rect 10998 31145 11008 31201
rect 11064 31145 11074 31201
rect 10998 31059 11074 31145
rect 10998 31003 11008 31059
rect 11064 31003 11074 31059
rect 11236 32642 11312 32652
rect 11236 32586 11246 32642
rect 11302 32586 11312 32642
rect 11236 32500 11312 32586
rect 11236 32444 11246 32500
rect 11302 32444 11312 32500
rect 11236 32358 11312 32444
rect 11236 32302 11246 32358
rect 11302 32302 11312 32358
rect 11236 32216 11312 32302
rect 11236 32160 11246 32216
rect 11302 32160 11312 32216
rect 11236 32074 11312 32160
rect 11236 32018 11246 32074
rect 11302 32018 11312 32074
rect 11236 31932 11312 32018
rect 11236 31876 11246 31932
rect 11302 31876 11312 31932
rect 11236 31790 11312 31876
rect 11236 31734 11246 31790
rect 11302 31734 11312 31790
rect 11236 31648 11312 31734
rect 11236 31592 11246 31648
rect 11302 31592 11312 31648
rect 11236 31506 11312 31592
rect 11236 31450 11246 31506
rect 11302 31450 11312 31506
rect 11236 31364 11312 31450
rect 11236 31308 11246 31364
rect 11302 31308 11312 31364
rect 11236 31222 11312 31308
rect 11236 31166 11246 31222
rect 11302 31166 11312 31222
rect 11236 31080 11312 31166
rect 11236 31024 11246 31080
rect 11302 31024 11312 31080
rect 11724 32637 11734 32693
rect 11790 32637 11800 32693
rect 11724 32551 11800 32637
rect 11724 32495 11734 32551
rect 11790 32495 11800 32551
rect 11724 32409 11800 32495
rect 11724 32353 11734 32409
rect 11790 32353 11800 32409
rect 11724 32267 11800 32353
rect 11724 32211 11734 32267
rect 11790 32211 11800 32267
rect 11724 32125 11800 32211
rect 11724 32069 11734 32125
rect 11790 32069 11800 32125
rect 11724 31983 11800 32069
rect 11724 31927 11734 31983
rect 11790 31927 11800 31983
rect 11724 31841 11800 31927
rect 11724 31785 11734 31841
rect 11790 31785 11800 31841
rect 11724 31699 11800 31785
rect 11724 31643 11734 31699
rect 11790 31643 11800 31699
rect 11724 31557 11800 31643
rect 11724 31501 11734 31557
rect 11790 31501 11800 31557
rect 11724 31415 11800 31501
rect 11724 31359 11734 31415
rect 11790 31359 11800 31415
rect 11724 31273 11800 31359
rect 11724 31217 11734 31273
rect 11790 31217 11800 31273
rect 11724 31131 11800 31217
rect 11724 31075 11734 31131
rect 11790 31075 11800 31131
rect 11724 31065 11800 31075
rect 12212 32692 12288 32702
rect 12212 32636 12222 32692
rect 12278 32636 12288 32692
rect 12212 32550 12288 32636
rect 12212 32494 12222 32550
rect 12278 32494 12288 32550
rect 12212 32408 12288 32494
rect 12212 32352 12222 32408
rect 12278 32352 12288 32408
rect 12212 32266 12288 32352
rect 12212 32210 12222 32266
rect 12278 32210 12288 32266
rect 12212 32124 12288 32210
rect 12212 32068 12222 32124
rect 12278 32068 12288 32124
rect 12212 31982 12288 32068
rect 12212 31926 12222 31982
rect 12278 31926 12288 31982
rect 12212 31840 12288 31926
rect 12212 31784 12222 31840
rect 12278 31784 12288 31840
rect 12212 31698 12288 31784
rect 12212 31642 12222 31698
rect 12278 31642 12288 31698
rect 12212 31556 12288 31642
rect 12212 31500 12222 31556
rect 12278 31500 12288 31556
rect 12212 31414 12288 31500
rect 12212 31358 12222 31414
rect 12278 31358 12288 31414
rect 12212 31272 12288 31358
rect 12212 31216 12222 31272
rect 12278 31216 12288 31272
rect 12212 31130 12288 31216
rect 12212 31074 12222 31130
rect 12278 31074 12288 31130
rect 11236 31014 11312 31024
rect 10998 30993 11074 31003
rect 7976 30932 7986 30988
rect 8042 30932 8052 30988
rect 7976 30846 8052 30932
rect 7976 30790 7986 30846
rect 8042 30790 8052 30846
rect 7976 30704 8052 30790
rect 7976 30648 7986 30704
rect 8042 30648 8052 30704
rect 7976 30562 8052 30648
rect 7976 30506 7986 30562
rect 8042 30506 8052 30562
rect 7976 30496 8052 30506
rect 12212 30988 12288 31074
rect 12212 30932 12222 30988
rect 12278 30932 12288 30988
rect 12212 30846 12288 30932
rect 12212 30790 12222 30846
rect 12278 30790 12288 30846
rect 12212 30704 12288 30790
rect 12212 30648 12222 30704
rect 12278 30648 12288 30704
rect 12212 30562 12288 30648
rect 12212 30506 12222 30562
rect 12278 30506 12288 30562
rect 12212 30496 12288 30506
rect 12628 32692 12704 32702
rect 12628 32636 12638 32692
rect 12694 32636 12704 32692
rect 12628 32550 12704 32636
rect 12628 32494 12638 32550
rect 12694 32494 12704 32550
rect 12628 32408 12704 32494
rect 12628 32352 12638 32408
rect 12694 32352 12704 32408
rect 12628 32266 12704 32352
rect 12628 32210 12638 32266
rect 12694 32210 12704 32266
rect 12628 32124 12704 32210
rect 12628 32068 12638 32124
rect 12694 32068 12704 32124
rect 12628 31982 12704 32068
rect 12628 31926 12638 31982
rect 12694 31926 12704 31982
rect 12628 31840 12704 31926
rect 12628 31784 12638 31840
rect 12694 31784 12704 31840
rect 12628 31698 12704 31784
rect 12628 31642 12638 31698
rect 12694 31642 12704 31698
rect 12628 31556 12704 31642
rect 12628 31500 12638 31556
rect 12694 31500 12704 31556
rect 12628 31414 12704 31500
rect 12628 31358 12638 31414
rect 12694 31358 12704 31414
rect 12628 31272 12704 31358
rect 12628 31216 12638 31272
rect 12694 31216 12704 31272
rect 12628 31130 12704 31216
rect 12628 31074 12638 31130
rect 12694 31074 12704 31130
rect 12628 30988 12704 31074
rect 12628 30932 12638 30988
rect 12694 30932 12704 30988
rect 12628 30846 12704 30932
rect 12628 30790 12638 30846
rect 12694 30790 12704 30846
rect 12628 30704 12704 30790
rect 12628 30648 12638 30704
rect 12694 30648 12704 30704
rect 12628 30562 12704 30648
rect 12628 30506 12638 30562
rect 12694 30506 12704 30562
rect 12628 30496 12704 30506
rect 14020 32692 14096 32702
rect 14020 32636 14030 32692
rect 14086 32636 14096 32692
rect 14020 32550 14096 32636
rect 14020 32494 14030 32550
rect 14086 32494 14096 32550
rect 14020 32408 14096 32494
rect 14020 32352 14030 32408
rect 14086 32352 14096 32408
rect 14020 32266 14096 32352
rect 14020 32210 14030 32266
rect 14086 32210 14096 32266
rect 14020 32124 14096 32210
rect 14020 32068 14030 32124
rect 14086 32068 14096 32124
rect 14020 31982 14096 32068
rect 14020 31926 14030 31982
rect 14086 31926 14096 31982
rect 14020 31840 14096 31926
rect 14020 31784 14030 31840
rect 14086 31784 14096 31840
rect 14020 31698 14096 31784
rect 14020 31642 14030 31698
rect 14086 31642 14096 31698
rect 14020 31556 14096 31642
rect 14020 31500 14030 31556
rect 14086 31500 14096 31556
rect 14020 31414 14096 31500
rect 14020 31358 14030 31414
rect 14086 31358 14096 31414
rect 14020 31272 14096 31358
rect 14020 31216 14030 31272
rect 14086 31216 14096 31272
rect 14020 31130 14096 31216
rect 14020 31074 14030 31130
rect 14086 31074 14096 31130
rect 14020 30988 14096 31074
rect 14020 30932 14030 30988
rect 14086 30932 14096 30988
rect 14020 30846 14096 30932
rect 14020 30790 14030 30846
rect 14086 30790 14096 30846
rect 14020 30704 14096 30790
rect 14020 30648 14030 30704
rect 14086 30648 14096 30704
rect 14020 30562 14096 30648
rect 14020 30506 14030 30562
rect 14086 30506 14096 30562
rect 14020 30496 14096 30506
rect 14400 32638 14760 32724
rect 14400 32582 14410 32638
rect 14466 32582 14552 32638
rect 14608 32582 14694 32638
rect 14750 32582 14760 32638
rect 14400 32496 14760 32582
rect 14400 32440 14410 32496
rect 14466 32440 14552 32496
rect 14608 32440 14694 32496
rect 14750 32440 14760 32496
rect 14400 32354 14760 32440
rect 14400 32298 14410 32354
rect 14466 32298 14552 32354
rect 14608 32298 14694 32354
rect 14750 32298 14760 32354
rect 14400 32212 14760 32298
rect 14400 32156 14410 32212
rect 14466 32156 14552 32212
rect 14608 32156 14694 32212
rect 14750 32156 14760 32212
rect 14400 32070 14760 32156
rect 14400 32014 14410 32070
rect 14466 32014 14552 32070
rect 14608 32014 14694 32070
rect 14750 32014 14760 32070
rect 14400 31928 14760 32014
rect 14400 31872 14410 31928
rect 14466 31872 14552 31928
rect 14608 31872 14694 31928
rect 14750 31872 14760 31928
rect 14400 31786 14760 31872
rect 14400 31730 14410 31786
rect 14466 31730 14552 31786
rect 14608 31730 14694 31786
rect 14750 31730 14760 31786
rect 14400 31644 14760 31730
rect 14400 31588 14410 31644
rect 14466 31588 14552 31644
rect 14608 31588 14694 31644
rect 14750 31588 14760 31644
rect 14400 31502 14760 31588
rect 14400 31446 14410 31502
rect 14466 31446 14552 31502
rect 14608 31446 14694 31502
rect 14750 31446 14760 31502
rect 14400 31360 14760 31446
rect 14400 31304 14410 31360
rect 14466 31304 14552 31360
rect 14608 31304 14694 31360
rect 14750 31304 14760 31360
rect 14400 31218 14760 31304
rect 14400 31162 14410 31218
rect 14466 31162 14552 31218
rect 14608 31162 14694 31218
rect 14750 31162 14760 31218
rect 14400 31076 14760 31162
rect 14400 31020 14410 31076
rect 14466 31020 14552 31076
rect 14608 31020 14694 31076
rect 14750 31020 14760 31076
rect 14400 30934 14760 31020
rect 14400 30878 14410 30934
rect 14466 30878 14552 30934
rect 14608 30878 14694 30934
rect 14750 30878 14760 30934
rect 14400 30792 14760 30878
rect 14400 30736 14410 30792
rect 14466 30736 14552 30792
rect 14608 30736 14694 30792
rect 14750 30736 14760 30792
rect 14400 30650 14760 30736
rect 14400 30594 14410 30650
rect 14466 30594 14552 30650
rect 14608 30594 14694 30650
rect 14750 30594 14760 30650
rect 14400 30508 14760 30594
rect 486 30442 562 30452
rect 14400 30452 14410 30508
rect 14466 30452 14552 30508
rect 14608 30452 14694 30508
rect 14750 30452 14760 30508
rect 14400 30442 14760 30452
rect 14400 30167 14760 30177
rect 1985 30109 3339 30119
rect 1985 30053 1995 30109
rect 2051 30053 2137 30109
rect 2193 30053 2279 30109
rect 2335 30053 2421 30109
rect 2477 30053 2563 30109
rect 2619 30053 2705 30109
rect 2761 30053 2847 30109
rect 2903 30053 2989 30109
rect 3045 30053 3131 30109
rect 3187 30053 3273 30109
rect 3329 30053 3339 30109
rect 1985 30043 3339 30053
rect 11922 30109 13276 30119
rect 11922 30053 11932 30109
rect 11988 30053 12074 30109
rect 12130 30053 12216 30109
rect 12272 30053 12358 30109
rect 12414 30053 12500 30109
rect 12556 30053 12642 30109
rect 12698 30053 12784 30109
rect 12840 30053 12926 30109
rect 12982 30053 13068 30109
rect 13124 30053 13210 30109
rect 13266 30053 13276 30109
rect 11922 30043 13276 30053
rect 14400 30111 14410 30167
rect 14466 30111 14552 30167
rect 14608 30111 14694 30167
rect 14750 30111 14760 30167
rect 14400 30025 14760 30111
rect 14400 29969 14410 30025
rect 14466 29969 14552 30025
rect 14608 29969 14694 30025
rect 14750 29969 14760 30025
rect 14400 29883 14760 29969
rect 14400 29827 14410 29883
rect 14466 29827 14552 29883
rect 14608 29827 14694 29883
rect 14750 29827 14760 29883
rect 14400 29741 14760 29827
rect 14400 29685 14410 29741
rect 14466 29685 14552 29741
rect 14608 29685 14694 29741
rect 14750 29685 14760 29741
rect 14400 29599 14760 29685
rect 14400 29543 14410 29599
rect 14466 29543 14552 29599
rect 14608 29543 14694 29599
rect 14750 29543 14760 29599
rect 14400 29457 14760 29543
rect 14400 29401 14410 29457
rect 14466 29401 14552 29457
rect 14608 29401 14694 29457
rect 14750 29401 14760 29457
rect 14400 29315 14760 29401
rect 14400 29259 14410 29315
rect 14466 29259 14552 29315
rect 14608 29259 14694 29315
rect 14750 29259 14760 29315
rect 14400 29173 14760 29259
rect 14400 29117 14410 29173
rect 14466 29117 14552 29173
rect 14608 29117 14694 29173
rect 14750 29117 14760 29173
rect 14400 29031 14760 29117
rect 14400 28975 14410 29031
rect 14466 28975 14552 29031
rect 14608 28975 14694 29031
rect 14750 28975 14760 29031
rect 14400 28889 14760 28975
rect 14400 28833 14410 28889
rect 14466 28833 14552 28889
rect 14608 28833 14694 28889
rect 14750 28833 14760 28889
rect 14400 28823 14760 28833
rect 165 28567 383 28577
rect 165 28511 175 28567
rect 231 28511 317 28567
rect 373 28511 383 28567
rect 165 28425 383 28511
rect 165 28369 175 28425
rect 231 28369 317 28425
rect 373 28369 383 28425
rect 165 28283 383 28369
rect 165 28227 175 28283
rect 231 28227 317 28283
rect 373 28227 383 28283
rect 165 28141 383 28227
rect 165 28085 175 28141
rect 231 28085 317 28141
rect 373 28085 383 28141
rect 165 27999 383 28085
rect 165 27943 175 27999
rect 231 27943 317 27999
rect 373 27943 383 27999
rect 165 27857 383 27943
rect 165 27801 175 27857
rect 231 27801 317 27857
rect 373 27801 383 27857
rect 165 27715 383 27801
rect 165 27659 175 27715
rect 231 27659 317 27715
rect 373 27659 383 27715
rect 165 27573 383 27659
rect 165 27517 175 27573
rect 231 27517 317 27573
rect 373 27517 383 27573
rect 165 27431 383 27517
rect 165 27375 175 27431
rect 231 27375 317 27431
rect 373 27375 383 27431
rect 165 27289 383 27375
rect 165 27233 175 27289
rect 231 27233 317 27289
rect 373 27233 383 27289
rect 165 27223 383 27233
rect 14400 26948 14760 26958
rect 14400 26892 14410 26948
rect 14466 26892 14552 26948
rect 14608 26892 14694 26948
rect 14750 26892 14760 26948
rect 14400 26806 14760 26892
rect 14400 26750 14410 26806
rect 14466 26750 14552 26806
rect 14608 26750 14694 26806
rect 14750 26750 14760 26806
rect 14400 26664 14760 26750
rect 14400 26608 14410 26664
rect 14466 26608 14552 26664
rect 14608 26608 14694 26664
rect 14750 26608 14760 26664
rect 14400 26522 14760 26608
rect 14400 26466 14410 26522
rect 14466 26466 14552 26522
rect 14608 26466 14694 26522
rect 14750 26466 14760 26522
rect 14400 26380 14760 26466
rect 14400 26324 14410 26380
rect 14466 26324 14552 26380
rect 14608 26324 14694 26380
rect 14750 26324 14760 26380
rect 14400 26238 14760 26324
rect 14400 26182 14410 26238
rect 14466 26182 14552 26238
rect 14608 26182 14694 26238
rect 14750 26182 14760 26238
rect 14400 26096 14760 26182
rect 14400 26040 14410 26096
rect 14466 26040 14552 26096
rect 14608 26040 14694 26096
rect 14750 26040 14760 26096
rect 14400 25954 14760 26040
rect 14400 25898 14410 25954
rect 14466 25898 14552 25954
rect 14608 25898 14694 25954
rect 14750 25898 14760 25954
rect 14400 25812 14760 25898
rect 14400 25756 14410 25812
rect 14466 25756 14552 25812
rect 14608 25756 14694 25812
rect 14750 25756 14760 25812
rect 14400 25670 14760 25756
rect 14400 25614 14410 25670
rect 14466 25614 14552 25670
rect 14608 25614 14694 25670
rect 14750 25614 14760 25670
rect 14400 25528 14760 25614
rect 14400 25472 14410 25528
rect 14466 25472 14552 25528
rect 14608 25472 14694 25528
rect 14750 25472 14760 25528
rect 14400 25386 14760 25472
rect 14400 25330 14410 25386
rect 14466 25330 14552 25386
rect 14608 25330 14694 25386
rect 14750 25330 14760 25386
rect 14400 25244 14760 25330
rect 14400 25188 14410 25244
rect 14466 25188 14552 25244
rect 14608 25188 14694 25244
rect 14750 25188 14760 25244
rect 14400 25102 14760 25188
rect 14400 25046 14410 25102
rect 14466 25046 14552 25102
rect 14608 25046 14694 25102
rect 14750 25046 14760 25102
rect 14400 24960 14760 25046
rect 14400 24904 14410 24960
rect 14466 24904 14552 24960
rect 14608 24904 14694 24960
rect 14750 24904 14760 24960
rect 14400 24818 14760 24904
rect 14400 24762 14410 24818
rect 14466 24762 14552 24818
rect 14608 24762 14694 24818
rect 14750 24762 14760 24818
rect 14400 24676 14760 24762
rect 14400 24620 14410 24676
rect 14466 24620 14552 24676
rect 14608 24620 14694 24676
rect 14750 24620 14760 24676
rect 14400 24534 14760 24620
rect 14400 24478 14410 24534
rect 14466 24478 14552 24534
rect 14608 24478 14694 24534
rect 14750 24478 14760 24534
rect 14400 24392 14760 24478
rect 14400 24336 14410 24392
rect 14466 24336 14552 24392
rect 14608 24336 14694 24392
rect 14750 24336 14760 24392
rect 14400 24250 14760 24336
rect 14400 24194 14410 24250
rect 14466 24194 14552 24250
rect 14608 24194 14694 24250
rect 14750 24194 14760 24250
rect 14400 24108 14760 24194
rect 14400 24052 14410 24108
rect 14466 24052 14552 24108
rect 14608 24052 14694 24108
rect 14750 24052 14760 24108
rect 14400 24042 14760 24052
rect 14400 23748 14760 23758
rect 14400 23692 14410 23748
rect 14466 23692 14552 23748
rect 14608 23692 14694 23748
rect 14750 23692 14760 23748
rect 14400 23606 14760 23692
rect 14400 23550 14410 23606
rect 14466 23550 14552 23606
rect 14608 23550 14694 23606
rect 14750 23550 14760 23606
rect 14400 23464 14760 23550
rect 14400 23408 14410 23464
rect 14466 23408 14552 23464
rect 14608 23408 14694 23464
rect 14750 23408 14760 23464
rect 14400 23322 14760 23408
rect 14400 23266 14410 23322
rect 14466 23266 14552 23322
rect 14608 23266 14694 23322
rect 14750 23266 14760 23322
rect 14400 23180 14760 23266
rect 14400 23124 14410 23180
rect 14466 23124 14552 23180
rect 14608 23124 14694 23180
rect 14750 23124 14760 23180
rect 14400 23038 14760 23124
rect 14400 22982 14410 23038
rect 14466 22982 14552 23038
rect 14608 22982 14694 23038
rect 14750 22982 14760 23038
rect 14400 22896 14760 22982
rect 14400 22840 14410 22896
rect 14466 22840 14552 22896
rect 14608 22840 14694 22896
rect 14750 22840 14760 22896
rect 14400 22754 14760 22840
rect 14400 22698 14410 22754
rect 14466 22698 14552 22754
rect 14608 22698 14694 22754
rect 14750 22698 14760 22754
rect 14400 22612 14760 22698
rect 14400 22556 14410 22612
rect 14466 22556 14552 22612
rect 14608 22556 14694 22612
rect 14750 22556 14760 22612
rect 14400 22470 14760 22556
rect 14400 22414 14410 22470
rect 14466 22414 14552 22470
rect 14608 22414 14694 22470
rect 14750 22414 14760 22470
rect 14400 22328 14760 22414
rect 14400 22272 14410 22328
rect 14466 22272 14552 22328
rect 14608 22272 14694 22328
rect 14750 22272 14760 22328
rect 14400 22186 14760 22272
rect 14400 22130 14410 22186
rect 14466 22130 14552 22186
rect 14608 22130 14694 22186
rect 14750 22130 14760 22186
rect 14400 22044 14760 22130
rect 14400 21988 14410 22044
rect 14466 21988 14552 22044
rect 14608 21988 14694 22044
rect 14750 21988 14760 22044
rect 14400 21902 14760 21988
rect 14400 21846 14410 21902
rect 14466 21846 14552 21902
rect 14608 21846 14694 21902
rect 14750 21846 14760 21902
rect 14400 21760 14760 21846
rect 14400 21704 14410 21760
rect 14466 21704 14552 21760
rect 14608 21704 14694 21760
rect 14750 21704 14760 21760
rect 14400 21618 14760 21704
rect 14400 21562 14410 21618
rect 14466 21562 14552 21618
rect 14608 21562 14694 21618
rect 14750 21562 14760 21618
rect 14400 21476 14760 21562
rect 14400 21420 14410 21476
rect 14466 21420 14552 21476
rect 14608 21420 14694 21476
rect 14750 21420 14760 21476
rect 14400 21334 14760 21420
rect 14400 21278 14410 21334
rect 14466 21278 14552 21334
rect 14608 21278 14694 21334
rect 14750 21278 14760 21334
rect 14400 21192 14760 21278
rect 14400 21136 14410 21192
rect 14466 21136 14552 21192
rect 14608 21136 14694 21192
rect 14750 21136 14760 21192
rect 14400 21050 14760 21136
rect 14400 20994 14410 21050
rect 14466 20994 14552 21050
rect 14608 20994 14694 21050
rect 14750 20994 14760 21050
rect 14400 20908 14760 20994
rect 14400 20852 14410 20908
rect 14466 20852 14552 20908
rect 14608 20852 14694 20908
rect 14750 20852 14760 20908
rect 14400 20842 14760 20852
rect 14400 20548 14760 20558
rect 14400 20492 14410 20548
rect 14466 20492 14552 20548
rect 14608 20492 14694 20548
rect 14750 20492 14760 20548
rect 14400 20406 14760 20492
rect 14400 20350 14410 20406
rect 14466 20350 14552 20406
rect 14608 20350 14694 20406
rect 14750 20350 14760 20406
rect 14400 20264 14760 20350
rect 14400 20208 14410 20264
rect 14466 20208 14552 20264
rect 14608 20208 14694 20264
rect 14750 20208 14760 20264
rect 14400 20122 14760 20208
rect 14400 20066 14410 20122
rect 14466 20066 14552 20122
rect 14608 20066 14694 20122
rect 14750 20066 14760 20122
rect 14400 19980 14760 20066
rect 14400 19924 14410 19980
rect 14466 19924 14552 19980
rect 14608 19924 14694 19980
rect 14750 19924 14760 19980
rect 14400 19838 14760 19924
rect 14400 19782 14410 19838
rect 14466 19782 14552 19838
rect 14608 19782 14694 19838
rect 14750 19782 14760 19838
rect 14400 19696 14760 19782
rect 14400 19640 14410 19696
rect 14466 19640 14552 19696
rect 14608 19640 14694 19696
rect 14750 19640 14760 19696
rect 14400 19554 14760 19640
rect 14400 19498 14410 19554
rect 14466 19498 14552 19554
rect 14608 19498 14694 19554
rect 14750 19498 14760 19554
rect 14400 19412 14760 19498
rect 14400 19356 14410 19412
rect 14466 19356 14552 19412
rect 14608 19356 14694 19412
rect 14750 19356 14760 19412
rect 14400 19270 14760 19356
rect 14400 19214 14410 19270
rect 14466 19214 14552 19270
rect 14608 19214 14694 19270
rect 14750 19214 14760 19270
rect 14400 19128 14760 19214
rect 14400 19072 14410 19128
rect 14466 19072 14552 19128
rect 14608 19072 14694 19128
rect 14750 19072 14760 19128
rect 14400 18986 14760 19072
rect 14400 18930 14410 18986
rect 14466 18930 14552 18986
rect 14608 18930 14694 18986
rect 14750 18930 14760 18986
rect 14400 18844 14760 18930
rect 14400 18788 14410 18844
rect 14466 18788 14552 18844
rect 14608 18788 14694 18844
rect 14750 18788 14760 18844
rect 14400 18702 14760 18788
rect 14400 18646 14410 18702
rect 14466 18646 14552 18702
rect 14608 18646 14694 18702
rect 14750 18646 14760 18702
rect 14400 18560 14760 18646
rect 14400 18504 14410 18560
rect 14466 18504 14552 18560
rect 14608 18504 14694 18560
rect 14750 18504 14760 18560
rect 14400 18418 14760 18504
rect 14400 18362 14410 18418
rect 14466 18362 14552 18418
rect 14608 18362 14694 18418
rect 14750 18362 14760 18418
rect 14400 18276 14760 18362
rect 14400 18220 14410 18276
rect 14466 18220 14552 18276
rect 14608 18220 14694 18276
rect 14750 18220 14760 18276
rect 14400 18134 14760 18220
rect 14400 18078 14410 18134
rect 14466 18078 14552 18134
rect 14608 18078 14694 18134
rect 14750 18078 14760 18134
rect 14400 17992 14760 18078
rect 14400 17936 14410 17992
rect 14466 17936 14552 17992
rect 14608 17936 14694 17992
rect 14750 17936 14760 17992
rect 14400 17850 14760 17936
rect 14400 17794 14410 17850
rect 14466 17794 14552 17850
rect 14608 17794 14694 17850
rect 14750 17794 14760 17850
rect 14400 17708 14760 17794
rect 14400 17652 14410 17708
rect 14466 17652 14552 17708
rect 14608 17652 14694 17708
rect 14750 17652 14760 17708
rect 14400 17642 14760 17652
rect 14400 17348 14760 17358
rect 14400 17292 14410 17348
rect 14466 17292 14552 17348
rect 14608 17292 14694 17348
rect 14750 17292 14760 17348
rect 14400 17206 14760 17292
rect 14400 17150 14410 17206
rect 14466 17150 14552 17206
rect 14608 17150 14694 17206
rect 14750 17150 14760 17206
rect 14400 17064 14760 17150
rect 14400 17008 14410 17064
rect 14466 17008 14552 17064
rect 14608 17008 14694 17064
rect 14750 17008 14760 17064
rect 14400 16922 14760 17008
rect 14400 16866 14410 16922
rect 14466 16866 14552 16922
rect 14608 16866 14694 16922
rect 14750 16866 14760 16922
rect 14400 16780 14760 16866
rect 14400 16724 14410 16780
rect 14466 16724 14552 16780
rect 14608 16724 14694 16780
rect 14750 16724 14760 16780
rect 14400 16638 14760 16724
rect 14400 16582 14410 16638
rect 14466 16582 14552 16638
rect 14608 16582 14694 16638
rect 14750 16582 14760 16638
rect 14400 16496 14760 16582
rect 14400 16440 14410 16496
rect 14466 16440 14552 16496
rect 14608 16440 14694 16496
rect 14750 16440 14760 16496
rect 14400 16354 14760 16440
rect 14400 16298 14410 16354
rect 14466 16298 14552 16354
rect 14608 16298 14694 16354
rect 14750 16298 14760 16354
rect 14400 16212 14760 16298
rect 14400 16156 14410 16212
rect 14466 16156 14552 16212
rect 14608 16156 14694 16212
rect 14750 16156 14760 16212
rect 14400 16070 14760 16156
rect 14400 16014 14410 16070
rect 14466 16014 14552 16070
rect 14608 16014 14694 16070
rect 14750 16014 14760 16070
rect 14400 15928 14760 16014
rect 14400 15872 14410 15928
rect 14466 15872 14552 15928
rect 14608 15872 14694 15928
rect 14750 15872 14760 15928
rect 14400 15786 14760 15872
rect 14400 15730 14410 15786
rect 14466 15730 14552 15786
rect 14608 15730 14694 15786
rect 14750 15730 14760 15786
rect 14400 15644 14760 15730
rect 14400 15588 14410 15644
rect 14466 15588 14552 15644
rect 14608 15588 14694 15644
rect 14750 15588 14760 15644
rect 14400 15502 14760 15588
rect 14400 15446 14410 15502
rect 14466 15446 14552 15502
rect 14608 15446 14694 15502
rect 14750 15446 14760 15502
rect 14400 15360 14760 15446
rect 14400 15304 14410 15360
rect 14466 15304 14552 15360
rect 14608 15304 14694 15360
rect 14750 15304 14760 15360
rect 14400 15218 14760 15304
rect 14400 15162 14410 15218
rect 14466 15162 14552 15218
rect 14608 15162 14694 15218
rect 14750 15162 14760 15218
rect 14400 15076 14760 15162
rect 14400 15020 14410 15076
rect 14466 15020 14552 15076
rect 14608 15020 14694 15076
rect 14750 15020 14760 15076
rect 14400 14934 14760 15020
rect 14400 14878 14410 14934
rect 14466 14878 14552 14934
rect 14608 14878 14694 14934
rect 14750 14878 14760 14934
rect 14400 14792 14760 14878
rect 14400 14736 14410 14792
rect 14466 14736 14552 14792
rect 14608 14736 14694 14792
rect 14750 14736 14760 14792
rect 14400 14650 14760 14736
rect 14400 14594 14410 14650
rect 14466 14594 14552 14650
rect 14608 14594 14694 14650
rect 14750 14594 14760 14650
rect 14400 14508 14760 14594
rect 14400 14452 14410 14508
rect 14466 14452 14552 14508
rect 14608 14452 14694 14508
rect 14750 14452 14760 14508
rect 14400 14442 14760 14452
rect 165 10948 383 10958
rect 165 10892 175 10948
rect 231 10892 317 10948
rect 373 10892 383 10948
rect 165 10806 383 10892
rect 165 10750 175 10806
rect 231 10750 317 10806
rect 373 10750 383 10806
rect 165 10664 383 10750
rect 165 10608 175 10664
rect 231 10608 317 10664
rect 373 10608 383 10664
rect 165 10522 383 10608
rect 165 10466 175 10522
rect 231 10466 317 10522
rect 373 10466 383 10522
rect 165 10380 383 10466
rect 165 10324 175 10380
rect 231 10324 317 10380
rect 373 10324 383 10380
rect 165 10238 383 10324
rect 165 10182 175 10238
rect 231 10182 317 10238
rect 373 10182 383 10238
rect 165 10096 383 10182
rect 165 10040 175 10096
rect 231 10040 317 10096
rect 373 10040 383 10096
rect 165 9954 383 10040
rect 165 9898 175 9954
rect 231 9898 317 9954
rect 373 9898 383 9954
rect 165 9812 383 9898
rect 165 9756 175 9812
rect 231 9756 317 9812
rect 373 9756 383 9812
rect 165 9670 383 9756
rect 165 9614 175 9670
rect 231 9614 317 9670
rect 373 9614 383 9670
rect 165 9528 383 9614
rect 165 9472 175 9528
rect 231 9472 317 9528
rect 373 9472 383 9528
rect 165 9386 383 9472
rect 165 9330 175 9386
rect 231 9330 317 9386
rect 373 9330 383 9386
rect 165 9244 383 9330
rect 165 9188 175 9244
rect 231 9188 317 9244
rect 373 9188 383 9244
rect 165 9102 383 9188
rect 165 9046 175 9102
rect 231 9046 317 9102
rect 373 9046 383 9102
rect 165 8960 383 9046
rect 165 8904 175 8960
rect 231 8904 317 8960
rect 373 8904 383 8960
rect 165 8818 383 8904
rect 165 8762 175 8818
rect 231 8762 317 8818
rect 373 8762 383 8818
rect 165 8676 383 8762
rect 165 8620 175 8676
rect 231 8620 317 8676
rect 373 8620 383 8676
rect 165 8534 383 8620
rect 165 8478 175 8534
rect 231 8478 317 8534
rect 373 8478 383 8534
rect 165 8392 383 8478
rect 165 8336 175 8392
rect 231 8336 317 8392
rect 373 8336 383 8392
rect 165 8250 383 8336
rect 165 8194 175 8250
rect 231 8194 317 8250
rect 373 8194 383 8250
rect 165 8108 383 8194
rect 165 8052 175 8108
rect 231 8052 317 8108
rect 373 8052 383 8108
rect 165 8042 383 8052
rect 165 7748 383 7758
rect 165 7692 175 7748
rect 231 7692 317 7748
rect 373 7692 383 7748
rect 165 7606 383 7692
rect 165 7550 175 7606
rect 231 7550 317 7606
rect 373 7550 383 7606
rect 165 7464 383 7550
rect 165 7408 175 7464
rect 231 7408 317 7464
rect 373 7408 383 7464
rect 165 7322 383 7408
rect 165 7266 175 7322
rect 231 7266 317 7322
rect 373 7266 383 7322
rect 165 7180 383 7266
rect 165 7124 175 7180
rect 231 7124 317 7180
rect 373 7124 383 7180
rect 165 7038 383 7124
rect 165 6982 175 7038
rect 231 6982 317 7038
rect 373 6982 383 7038
rect 165 6896 383 6982
rect 165 6840 175 6896
rect 231 6840 317 6896
rect 373 6840 383 6896
rect 165 6754 383 6840
rect 165 6698 175 6754
rect 231 6698 317 6754
rect 373 6698 383 6754
rect 165 6612 383 6698
rect 165 6556 175 6612
rect 231 6556 317 6612
rect 373 6556 383 6612
rect 165 6470 383 6556
rect 165 6414 175 6470
rect 231 6414 317 6470
rect 373 6414 383 6470
rect 165 6328 383 6414
rect 165 6272 175 6328
rect 231 6272 317 6328
rect 373 6272 383 6328
rect 165 6186 383 6272
rect 165 6130 175 6186
rect 231 6130 317 6186
rect 373 6130 383 6186
rect 165 6044 383 6130
rect 165 5988 175 6044
rect 231 5988 317 6044
rect 373 5988 383 6044
rect 165 5902 383 5988
rect 165 5846 175 5902
rect 231 5846 317 5902
rect 373 5846 383 5902
rect 165 5760 383 5846
rect 165 5704 175 5760
rect 231 5704 317 5760
rect 373 5704 383 5760
rect 165 5618 383 5704
rect 165 5562 175 5618
rect 231 5562 317 5618
rect 373 5562 383 5618
rect 165 5476 383 5562
rect 165 5420 175 5476
rect 231 5420 317 5476
rect 373 5420 383 5476
rect 165 5334 383 5420
rect 165 5278 175 5334
rect 231 5278 317 5334
rect 373 5278 383 5334
rect 165 5192 383 5278
rect 165 5136 175 5192
rect 231 5136 317 5192
rect 373 5136 383 5192
rect 165 5050 383 5136
rect 165 4994 175 5050
rect 231 4994 317 5050
rect 373 4994 383 5050
rect 165 4908 383 4994
rect 165 4852 175 4908
rect 231 4852 317 4908
rect 373 4852 383 4908
rect 165 4842 383 4852
rect 165 4548 383 4558
rect 165 4492 175 4548
rect 231 4492 317 4548
rect 373 4492 383 4548
rect 165 4406 383 4492
rect 165 4350 175 4406
rect 231 4350 317 4406
rect 373 4350 383 4406
rect 165 4264 383 4350
rect 165 4208 175 4264
rect 231 4208 317 4264
rect 373 4208 383 4264
rect 165 4122 383 4208
rect 165 4066 175 4122
rect 231 4066 317 4122
rect 373 4066 383 4122
rect 165 3980 383 4066
rect 165 3924 175 3980
rect 231 3924 317 3980
rect 373 3924 383 3980
rect 165 3838 383 3924
rect 165 3782 175 3838
rect 231 3782 317 3838
rect 373 3782 383 3838
rect 165 3696 383 3782
rect 165 3640 175 3696
rect 231 3640 317 3696
rect 373 3640 383 3696
rect 165 3554 383 3640
rect 165 3498 175 3554
rect 231 3498 317 3554
rect 373 3498 383 3554
rect 165 3412 383 3498
rect 165 3356 175 3412
rect 231 3356 317 3412
rect 373 3356 383 3412
rect 165 3270 383 3356
rect 165 3214 175 3270
rect 231 3214 317 3270
rect 373 3214 383 3270
rect 165 3128 383 3214
rect 165 3072 175 3128
rect 231 3072 317 3128
rect 373 3072 383 3128
rect 165 2986 383 3072
rect 165 2930 175 2986
rect 231 2930 317 2986
rect 373 2930 383 2986
rect 165 2844 383 2930
rect 165 2788 175 2844
rect 231 2788 317 2844
rect 373 2788 383 2844
rect 165 2702 383 2788
rect 165 2646 175 2702
rect 231 2646 317 2702
rect 373 2646 383 2702
rect 165 2560 383 2646
rect 165 2504 175 2560
rect 231 2504 317 2560
rect 373 2504 383 2560
rect 165 2418 383 2504
rect 165 2362 175 2418
rect 231 2362 317 2418
rect 373 2362 383 2418
rect 165 2276 383 2362
rect 165 2220 175 2276
rect 231 2220 317 2276
rect 373 2220 383 2276
rect 165 2134 383 2220
rect 165 2078 175 2134
rect 231 2078 317 2134
rect 373 2078 383 2134
rect 165 1992 383 2078
rect 165 1936 175 1992
rect 231 1936 317 1992
rect 373 1936 383 1992
rect 165 1850 383 1936
rect 165 1794 175 1850
rect 231 1794 317 1850
rect 373 1794 383 1850
rect 165 1708 383 1794
rect 165 1652 175 1708
rect 231 1652 317 1708
rect 373 1652 383 1708
rect 165 1642 383 1652
use comp018green_esd_cdm  comp018green_esd_cdm_0
timestamp 1698431365
transform 1 0 4583 0 -1 49459
box -205 -83 5981 8547
use comp018green_inpath_cms_smt  comp018green_inpath_cms_smt_0
timestamp 1698431365
transform 1 0 848 0 -1 55852
box -144 -83 13504 14940
use comp018green_out_paddrv_16T  comp018green_out_paddrv_16T_0
timestamp 1698431365
transform 1 0 794 0 1 1465
box -360 -1465 13796 27678
use comp018green_out_predrv  comp018green_out_predrv_0
timestamp 1698431365
transform 1 0 479 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_1
timestamp 1698431365
transform -1 0 14585 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_2
timestamp 1698431365
transform 1 0 7487 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_predrv  comp018green_out_predrv_3
timestamp 1698431365
transform -1 0 7577 0 -1 35969
box -83 -83 3677 6020
use comp018green_out_sigbuf_a  comp018green_out_sigbuf_a_0
timestamp 1698431365
transform -1 0 11282 0 1 37501
box -83 -83 2701 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_0
timestamp 1698431365
transform 1 0 798 0 1 37501
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_1
timestamp 1698431365
transform -1 0 6132 0 1 37501
box -83 -803 2795 2911
use comp018green_out_sigbuf_oe  comp018green_out_sigbuf_oe_2
timestamp 1698431365
transform 1 0 6042 0 1 37501
box -83 -803 2795 2911
use comp018green_sigbuf_1  comp018green_sigbuf_1_0
timestamp 1698431365
transform 1 0 11192 0 1 37501
box -83 -83 2889 2911
use M1_NWELL_CDNS_40661953145322  M1_NWELL_CDNS_40661953145322_0
timestamp 1698431365
transform 1 0 999 0 1 55135
box 0 0 1 1
use M1_NWELL_CDNS_40661953145377  M1_NWELL_CDNS_40661953145377_0
timestamp 1698431365
transform 1 0 482 0 1 55900
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145165  M1_PACTIVE_CDNS_40661953145165_0
timestamp 1698431365
transform 1 0 12098 0 1 42332
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145165  M1_PACTIVE_CDNS_40661953145165_1
timestamp 1698431365
transform 1 0 14615 0 1 42332
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145166  M1_PACTIVE_CDNS_40661953145166_0
timestamp 1698431365
transform 1 0 13333 0 1 41110
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145166  M1_PACTIVE_CDNS_40661953145166_1
timestamp 1698431365
transform 1 0 13333 0 1 43554
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145167  M1_PACTIVE_CDNS_40661953145167_0
timestamp 1698431365
transform 1 0 2376 0 1 56639
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145167  M1_PACTIVE_CDNS_40661953145167_1
timestamp 1698431365
transform 1 0 14690 0 1 56639
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145168  M1_PACTIVE_CDNS_40661953145168_0
timestamp 1698431365
transform 0 -1 8533 1 0 56099
box 0 0 1 1
use M1_PACTIVE_CDNS_40661953145168  M1_PACTIVE_CDNS_40661953145168_1
timestamp 1698431365
transform 0 -1 8533 1 0 57179
box 0 0 1 1
use M1_PSUB_CDNS_40661953145215  M1_PSUB_CDNS_40661953145215_0
timestamp 1698431365
transform 1 0 11300 0 1 43149
box 0 0 1 1
use M1_PSUB_CDNS_40661953145338  M1_PSUB_CDNS_40661953145338_0
timestamp 1698431365
transform 1 0 7502 0 1 1121
box 0 0 1 1
use M1_PSUB_CDNS_40661953145339  M1_PSUB_CDNS_40661953145339_0
timestamp 1698431365
transform 1 0 14768 0 1 6174
box 0 0 1 1
use M1_PSUB_CDNS_40661953145339  M1_PSUB_CDNS_40661953145339_1
timestamp 1698431365
transform -1 0 234 0 1 6174
box 0 0 1 1
use M2_M1_CDNS_40661953145112  M2_M1_CDNS_40661953145112_0
timestamp 1698431365
transform 1 0 4980 0 1 52653
box 0 0 1 1
use M2_M1_CDNS_40661953145112  M2_M1_CDNS_40661953145112_1
timestamp 1698431365
transform 1 0 6684 0 1 52653
box 0 0 1 1
use M2_M1_CDNS_40661953145114  M2_M1_CDNS_40661953145114_0
timestamp 1698431365
transform 1 0 10941 0 1 37542
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_0
timestamp 1698431365
transform 1 0 2760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_1
timestamp 1698431365
transform 1 0 7260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_2
timestamp 1698431365
transform 1 0 6760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_3
timestamp 1698431365
transform 1 0 5260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_4
timestamp 1698431365
transform 1 0 4260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_5
timestamp 1698431365
transform 1 0 5760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_6
timestamp 1698431365
transform 1 0 3760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_7
timestamp 1698431365
transform 1 0 8260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_8
timestamp 1698431365
transform 1 0 9760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_9
timestamp 1698431365
transform 1 0 10260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_10
timestamp 1698431365
transform 1 0 8760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_11
timestamp 1698431365
transform 1 0 11760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_12
timestamp 1698431365
transform 1 0 12760 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_13
timestamp 1698431365
transform 1 0 13260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_14
timestamp 1698431365
transform 1 0 14470 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_15
timestamp 1698431365
transform 1 0 11260 0 1 56637
box 0 0 1 1
use M2_M1_CDNS_40661953145116  M2_M1_CDNS_40661953145116_0
timestamp 1698431365
transform 1 0 524 0 1 31953
box 0 0 1 1
use M2_M1_CDNS_40661953145116  M2_M1_CDNS_40661953145116_1
timestamp 1698431365
transform 1 0 14540 0 1 31953
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_0
timestamp 1698431365
transform -1 0 4927 0 1 40708
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_1
timestamp 1698431365
transform -1 0 7143 0 1 40708
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_2
timestamp 1698431365
transform 1 0 5656 0 1 40542
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_3
timestamp 1698431365
transform -1 0 5484 0 1 36328
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_4
timestamp 1698431365
transform 1 0 6522 0 1 29791
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_5
timestamp 1698431365
transform -1 0 6144 0 1 36464
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_6
timestamp 1698431365
transform -1 0 5900 0 1 36600
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_7
timestamp 1698431365
transform -1 0 4551 0 1 36600
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_8
timestamp 1698431365
transform -1 0 6656 0 1 36192
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_9
timestamp 1698431365
transform 1 0 6766 0 1 29611
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_10
timestamp 1698431365
transform -1 0 4580 0 1 36056
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_11
timestamp 1698431365
transform 1 0 3476 0 1 36056
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_12
timestamp 1698431365
transform 1 0 1400 0 1 36192
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_13
timestamp 1698431365
transform 1 0 3181 0 1 36464
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_14
timestamp 1698431365
transform 1 0 2003 0 1 40708
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_15
timestamp 1698431365
transform 1 0 2572 0 1 36328
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_16
timestamp 1698431365
transform 1 0 1912 0 1 36464
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_17
timestamp 1698431365
transform 1 0 1686 0 1 40542
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_18
timestamp 1698431365
transform 1 0 1457 0 1 29791
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_19
timestamp 1698431365
transform 1 0 1637 0 1 29611
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_20
timestamp 1698431365
transform 1 0 3586 0 1 29404
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_21
timestamp 1698431365
transform 1 0 3456 0 1 52981
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_22
timestamp 1698431365
transform 1 0 1564 0 1 57301
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_23
timestamp 1698431365
transform 1 0 2683 0 1 55437
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_24
timestamp 1698431365
transform 1 0 7344 0 1 52653
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_25
timestamp 1698431365
transform 1 0 3773 0 1 52981
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_26
timestamp 1698431365
transform -1 0 3749 0 1 36464
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_27
timestamp 1698431365
transform -1 0 11480 0 1 29404
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_28
timestamp 1698431365
transform -1 0 12596 0 1 36328
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_29
timestamp 1698431365
transform 1 0 13012 0 1 36736
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_30
timestamp 1698431365
transform 1 0 13152 0 1 36872
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_31
timestamp 1698431365
transform -1 0 13664 0 1 36192
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_32
timestamp 1698431365
transform 1 0 13752 0 1 40572
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_33
timestamp 1698431365
transform 1 0 13898 0 1 40436
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_34
timestamp 1698431365
transform 1 0 11792 0 1 40857
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_35
timestamp 1698431365
transform 1 0 13425 0 1 36056
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_36
timestamp 1698431365
transform -1 0 11588 0 1 36056
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_37
timestamp 1698431365
transform 0 -1 11558 1 0 38607
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_38
timestamp 1698431365
transform 0 -1 14096 1 0 40760
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_39
timestamp 1698431365
transform 1 0 11506 0 1 40572
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_40
timestamp 1698431365
transform -1 0 13429 0 1 29611
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_41
timestamp 1698431365
transform -1 0 13609 0 1 29791
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_42
timestamp 1698431365
transform 1 0 12074 0 1 40436
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_43
timestamp 1698431365
transform 1 0 8408 0 1 36192
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_44
timestamp 1698431365
transform 1 0 8657 0 1 35920
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_45
timestamp 1698431365
transform 1 0 8383 0 1 36736
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_46
timestamp 1698431365
transform 1 0 10978 0 1 40708
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_47
timestamp 1698431365
transform 1 0 10484 0 1 36056
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_48
timestamp 1698431365
transform 1 0 8542 0 1 29611
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_49
timestamp 1698431365
transform 1 0 8786 0 1 29791
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_50
timestamp 1698431365
transform 1 0 10734 0 1 40436
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_51
timestamp 1698431365
transform 1 0 9580 0 1 36328
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_52
timestamp 1698431365
transform 1 0 8920 0 1 36464
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_53
timestamp 1698431365
transform -1 0 9060 0 1 36600
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_54
timestamp 1698431365
transform 0 -1 8477 1 0 36924
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_55
timestamp 1698431365
transform 1 0 12512 0 1 44027
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_0
timestamp 1698431365
transform 1 0 3646 0 1 42293
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_1
timestamp 1698431365
transform 1 0 84 0 1 37493
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_2
timestamp 1698431365
transform 1 0 3646 0 1 43893
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_3
timestamp 1698431365
transform 1 0 84 0 1 51893
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_4
timestamp 1698431365
transform 1 0 14980 0 1 37493
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_0
timestamp 1698431365
transform 1 0 14980 0 1 51893
box 0 0 1 1
use M2_M1_CDNS_40661953145125  M2_M1_CDNS_40661953145125_0
timestamp 1698431365
transform 1 0 13952 0 1 57301
box 0 0 1 1
use M2_M1_CDNS_40661953145161  M2_M1_CDNS_40661953145161_0
timestamp 1698431365
transform 1 0 13278 0 1 40288
box 0 0 1 1
use M2_M1_CDNS_40661953145163  M2_M1_CDNS_40661953145163_0
timestamp 1698431365
transform 1 0 3275 0 1 46270
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_0
timestamp 1698431365
transform -1 0 5952 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_1
timestamp 1698431365
transform 1 0 6196 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_2
timestamp 1698431365
transform 1 0 5952 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_3
timestamp 1698431365
transform -1 0 5536 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_4
timestamp 1698431365
transform 1 0 4193 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_5
timestamp 1698431365
transform -1 0 4998 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_6
timestamp 1698431365
transform -1 0 4185 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_7
timestamp 1698431365
transform -1 0 3697 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_8
timestamp 1698431365
transform 1 0 2520 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_9
timestamp 1698431365
transform 1 0 1860 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_10
timestamp 1698431365
transform 1 0 2104 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_11
timestamp 1698431365
transform 1 0 3233 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_12
timestamp 1698431365
transform 1 0 2745 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_13
timestamp 1698431365
transform 1 0 742 0 1 57249
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_14
timestamp 1698431365
transform 1 0 2347 0 1 55633
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_15
timestamp 1698431365
transform 1 0 13341 0 1 38597
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_16
timestamp 1698431365
transform 1 0 11609 0 1 41737
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_17
timestamp 1698431365
transform 1 0 11609 0 1 41263
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_18
timestamp 1698431365
transform 1 0 13134 0 1 42790
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_19
timestamp 1698431365
transform 1 0 13134 0 1 41863
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_20
timestamp 1698431365
transform 1 0 13570 0 1 41863
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_21
timestamp 1698431365
transform 1 0 13570 0 1 42790
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_22
timestamp 1698431365
transform 1 0 11324 0 1 41085
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_23
timestamp 1698431365
transform -1 0 13204 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_24
timestamp 1698431365
transform -1 0 12960 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_25
timestamp 1698431365
transform 1 0 13477 0 1 37945
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_26
timestamp 1698431365
transform -1 0 12544 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_27
timestamp 1698431365
transform -1 0 10873 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_28
timestamp 1698431365
transform -1 0 8868 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_29
timestamp 1698431365
transform -1 0 8477 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_30
timestamp 1698431365
transform -1 0 8331 0 1 38610
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_31
timestamp 1698431365
transform 1 0 10926 0 1 38968
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_32
timestamp 1698431365
transform 1 0 9528 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_33
timestamp 1698431365
transform 1 0 9112 0 1 34357
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_34
timestamp 1698431365
transform 1 0 10068 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_35
timestamp 1698431365
transform 1 0 9114 0 1 29391
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_36
timestamp 1698431365
transform 1 0 10682 0 1 38968
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_37
timestamp 1698431365
transform 1 0 8933 0 1 37861
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_38
timestamp 1698431365
transform 1 0 11055 0 1 40894
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_39
timestamp 1698431365
transform 1 0 14242 0 1 45915
box 0 0 1 1
use M2_M1_CDNS_40661953145164  M2_M1_CDNS_40661953145164_40
timestamp 1698431365
transform 1 0 11656 0 1 47864
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_0
timestamp 1698431365
transform 1 0 4200 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_1
timestamp 1698431365
transform 1 0 4788 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_2
timestamp 1698431365
transform 1 0 7480 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_3
timestamp 1698431365
transform 1 0 7292 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_4
timestamp 1698431365
transform 1 0 6804 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_5
timestamp 1698431365
transform 1 0 6316 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_6
timestamp 1698431365
transform 1 0 5952 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_7
timestamp 1698431365
transform 1 0 5464 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_8
timestamp 1698431365
transform 1 0 4976 0 1 55368
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_9
timestamp 1698431365
transform 1 0 8068 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_10
timestamp 1698431365
transform 1 0 10032 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_11
timestamp 1698431365
transform 1 0 11196 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_12
timestamp 1698431365
transform 1 0 10220 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_13
timestamp 1698431365
transform 1 0 10708 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_14
timestamp 1698431365
transform 1 0 12724 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_15
timestamp 1698431365
transform 1 0 13312 0 1 53773
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_16
timestamp 1698431365
transform 1 0 12048 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_17
timestamp 1698431365
transform 1 0 11560 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145169  M2_M1_CDNS_40661953145169_18
timestamp 1698431365
transform 1 0 12536 0 1 55377
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_0
timestamp 1698431365
transform 1 0 7480 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_1
timestamp 1698431365
transform 1 0 6134 0 1 53825
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_2
timestamp 1698431365
transform 1 0 6134 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_3
timestamp 1698431365
transform 1 0 4788 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_4
timestamp 1698431365
transform 1 0 10032 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_5
timestamp 1698431365
transform 1 0 12724 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_6
timestamp 1698431365
transform 1 0 13312 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_7
timestamp 1698431365
transform 1 0 11378 0 1 53825
box 0 0 1 1
use M2_M1_CDNS_40661953145171  M2_M1_CDNS_40661953145171_8
timestamp 1698431365
transform 1 0 11378 0 1 55287
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_0
timestamp 1698431365
transform 1 0 5121 0 1 39472
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_1
timestamp 1698431365
transform 1 0 7053 0 1 39472
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_2
timestamp 1698431365
transform 1 0 1809 0 1 39502
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_3
timestamp 1698431365
transform 1 0 5952 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_4
timestamp 1698431365
transform 1 0 6316 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_5
timestamp 1698431365
transform 1 0 6804 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_6
timestamp 1698431365
transform 1 0 7292 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_7
timestamp 1698431365
transform 1 0 4976 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_8
timestamp 1698431365
transform 1 0 5464 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_9
timestamp 1698431365
transform 1 0 11196 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_10
timestamp 1698431365
transform 1 0 11039 0 1 47432
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_11
timestamp 1698431365
transform 1 0 10220 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_12
timestamp 1698431365
transform 1 0 10708 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_13
timestamp 1698431365
transform 1 0 12536 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_14
timestamp 1698431365
transform 1 0 12048 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145173  M2_M1_CDNS_40661953145173_15
timestamp 1698431365
transform 1 0 11560 0 1 53716
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_0
timestamp 1698431365
transform 1 0 6087 0 1 38018
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_1
timestamp 1698431365
transform 1 0 6087 0 1 39264
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_2
timestamp 1698431365
transform 1 0 3465 0 1 38018
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_3
timestamp 1698431365
transform 1 0 843 0 1 38018
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_4
timestamp 1698431365
transform 1 0 3508 0 1 53877
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_5
timestamp 1698431365
transform 1 0 10365 0 1 39294
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_6
timestamp 1698431365
transform 1 0 8709 0 1 38018
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_7
timestamp 1698431365
transform 1 0 8068 0 1 55335
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_8
timestamp 1698431365
transform 1 0 9444 0 1 55335
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_9
timestamp 1698431365
transform 1 0 8975 0 1 55335
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_10
timestamp 1698431365
transform 1 0 8537 0 1 55335
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_11
timestamp 1698431365
transform 1 0 8752 0 1 55335
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_12
timestamp 1698431365
transform 1 0 8756 0 1 53877
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_13
timestamp 1698431365
transform 1 0 10820 0 1 48866
box 0 0 1 1
use M2_M1_CDNS_40661953145176  M2_M1_CDNS_40661953145176_14
timestamp 1698431365
transform 1 0 11238 0 1 39294
box 0 0 1 1
use M2_M1_CDNS_40661953145177  M2_M1_CDNS_40661953145177_0
timestamp 1698431365
transform 1 0 4794 0 1 48654
box 0 0 1 1
use M2_M1_CDNS_40661953145178  M2_M1_CDNS_40661953145178_0
timestamp 1698431365
transform 1 0 384 0 1 54945
box 0 0 1 1
use M2_M1_CDNS_40661953145178  M2_M1_CDNS_40661953145178_1
timestamp 1698431365
transform 1 0 384 0 1 54036
box 0 0 1 1
use M2_M1_CDNS_40661953145181  M2_M1_CDNS_40661953145181_0
timestamp 1698431365
transform 1 0 384 0 1 40280
box 0 0 1 1
use M2_M1_CDNS_40661953145181  M2_M1_CDNS_40661953145181_1
timestamp 1698431365
transform 1 0 2270 0 1 36600
box 0 0 1 1
use M2_M1_CDNS_40661953145181  M2_M1_CDNS_40661953145181_2
timestamp 1698431365
transform 1 0 904 0 1 52981
box 0 0 1 1
use M2_M1_CDNS_40661953145181  M2_M1_CDNS_40661953145181_3
timestamp 1698431365
transform 1 0 7914 0 1 50243
box 0 0 1 1
use M2_M1_CDNS_40661953145181  M2_M1_CDNS_40661953145181_4
timestamp 1698431365
transform 1 0 8616 0 1 50243
box 0 0 1 1
use M2_M1_CDNS_40661953145182  M2_M1_CDNS_40661953145182_0
timestamp 1698431365
transform 1 0 6616 0 1 49268
box 0 0 1 1
use M2_M1_CDNS_40661953145182  M2_M1_CDNS_40661953145182_1
timestamp 1698431365
transform 1 0 5713 0 1 49268
box 0 0 1 1
use M2_M1_CDNS_40661953145182  M2_M1_CDNS_40661953145182_2
timestamp 1698431365
transform 1 0 7914 0 1 49268
box 0 0 1 1
use M2_M1_CDNS_40661953145182  M2_M1_CDNS_40661953145182_3
timestamp 1698431365
transform 1 0 8616 0 1 49268
box 0 0 1 1
use M2_M1_CDNS_40661953145185  M2_M1_CDNS_40661953145185_0
timestamp 1698431365
transform 1 0 3646 0 1 47242
box 0 0 1 1
use M2_M1_CDNS_40661953145187  M2_M1_CDNS_40661953145187_0
timestamp 1698431365
transform 1 0 2758 0 1 41044
box 0 0 1 1
use M2_M1_CDNS_40661953145187  M2_M1_CDNS_40661953145187_1
timestamp 1698431365
transform 1 0 8810 0 1 40288
box 0 0 1 1
use M2_M1_CDNS_40661953145189  M2_M1_CDNS_40661953145189_0
timestamp 1698431365
transform 1 0 4028 0 1 31915
box 0 0 1 1
use M2_M1_CDNS_40661953145189  M2_M1_CDNS_40661953145189_1
timestamp 1698431365
transform 1 0 524 0 1 35036
box 0 0 1 1
use M2_M1_CDNS_40661953145189  M2_M1_CDNS_40661953145189_2
timestamp 1698431365
transform 1 0 11036 0 1 31915
box 0 0 1 1
use M2_M1_CDNS_40661953145195  M2_M1_CDNS_40661953145195_0
timestamp 1698431365
transform 1 0 4926 0 1 35244
box 0 0 1 1
use M2_M1_CDNS_40661953145195  M2_M1_CDNS_40661953145195_1
timestamp 1698431365
transform 1 0 3130 0 1 35244
box 0 0 1 1
use M2_M1_CDNS_40661953145195  M2_M1_CDNS_40661953145195_2
timestamp 1698431365
transform 1 0 762 0 1 35244
box 0 0 1 1
use M2_M1_CDNS_40661953145195  M2_M1_CDNS_40661953145195_3
timestamp 1698431365
transform 1 0 11934 0 1 35244
box 0 0 1 1
use M2_M1_CDNS_40661953145195  M2_M1_CDNS_40661953145195_4
timestamp 1698431365
transform 1 0 10138 0 1 35244
box 0 0 1 1
use M2_M1_CDNS_40661953145198  M2_M1_CDNS_40661953145198_0
timestamp 1698431365
transform 1 0 4028 0 1 34620
box 0 0 1 1
use M2_M1_CDNS_40661953145198  M2_M1_CDNS_40661953145198_1
timestamp 1698431365
transform 1 0 11036 0 1 34620
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_0
timestamp 1698431365
transform 1 0 7050 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_1
timestamp 1698431365
transform 1 0 1006 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_2
timestamp 1698431365
transform 1 0 2398 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_3
timestamp 1698431365
transform 1 0 2814 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_4
timestamp 1698431365
transform 1 0 12250 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_5
timestamp 1698431365
transform 1 0 12666 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_6
timestamp 1698431365
transform 1 0 14058 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145201  M2_M1_CDNS_40661953145201_7
timestamp 1698431365
transform 1 0 8014 0 1 31572
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_0
timestamp 1698431365
transform 1 0 5658 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_1
timestamp 1698431365
transform 1 0 5242 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_2
timestamp 1698431365
transform 1 0 4754 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_3
timestamp 1698431365
transform 1 0 4266 0 1 31834
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_4
timestamp 1698431365
transform 1 0 3302 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_5
timestamp 1698431365
transform 1 0 3790 0 1 31834
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_6
timestamp 1698431365
transform 1 0 11762 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_7
timestamp 1698431365
transform 1 0 10798 0 1 31834
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_8
timestamp 1698431365
transform 1 0 10310 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_9
timestamp 1698431365
transform 1 0 9822 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_10
timestamp 1698431365
transform 1 0 9406 0 1 31884
box 0 0 1 1
use M2_M1_CDNS_40661953145203  M2_M1_CDNS_40661953145203_11
timestamp 1698431365
transform 1 0 11274 0 1 31834
box 0 0 1 1
use M2_M1_CDNS_40661953145205  M2_M1_CDNS_40661953145205_0
timestamp 1698431365
transform 1 0 2662 0 1 30081
box 0 0 1 1
use M2_M1_CDNS_40661953145205  M2_M1_CDNS_40661953145205_1
timestamp 1698431365
transform 1 0 12599 0 1 30081
box 0 0 1 1
use M2_M1_CDNS_40661953145211  M2_M1_CDNS_40661953145211_0
timestamp 1698431365
transform 1 0 8066 0 1 56268
box 0 0 1 1
use M2_M1_CDNS_40661953145211  M2_M1_CDNS_40661953145211_1
timestamp 1698431365
transform 1 0 8066 0 1 57010
box 0 0 1 1
use M2_M1_CDNS_40661953145214  M2_M1_CDNS_40661953145214_0
timestamp 1698431365
transform 1 0 3459 0 1 40288
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_0
timestamp 1698431365
transform 1 0 6562 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_1
timestamp 1698431365
transform 1 0 4510 0 1 30676
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_2
timestamp 1698431365
transform 1 0 6806 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_3
timestamp 1698431365
transform 1 0 4998 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_4
timestamp 1698431365
transform 1 0 3546 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_5
timestamp 1698431365
transform 1 0 3058 0 1 30676
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_6
timestamp 1698431365
transform 1 0 1738 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_7
timestamp 1698431365
transform 1 0 1494 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_8
timestamp 1698431365
transform -1 0 11518 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_9
timestamp 1698431365
transform -1 0 12006 0 1 30676
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_10
timestamp 1698431365
transform -1 0 13570 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_11
timestamp 1698431365
transform -1 0 13814 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_12
timestamp 1698431365
transform -1 0 10554 0 1 30676
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_13
timestamp 1698431365
transform -1 0 10066 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_14
timestamp 1698431365
transform 1 0 8502 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145216  M2_M1_CDNS_40661953145216_15
timestamp 1698431365
transform 1 0 8746 0 1 30496
box 0 0 1 1
use M2_M1_CDNS_40661953145329  M2_M1_CDNS_40661953145329_0
timestamp 1698431365
transform 1 0 4334 0 1 50243
box 0 0 1 1
use M2_M1_CDNS_40661953145331  M2_M1_CDNS_40661953145331_0
timestamp 1698431365
transform 1 0 12460 0 1 46940
box 0 0 1 1
use M2_M1_CDNS_40661953145333  M2_M1_CDNS_40661953145333_0
timestamp 1698431365
transform 1 0 14472 0 1 49062
box 0 0 1 1
use M2_M1_CDNS_40661953145333  M2_M1_CDNS_40661953145333_1
timestamp 1698431365
transform 1 0 14472 0 1 48094
box 0 0 1 1
use M2_M1_CDNS_40661953145378  M2_M1_CDNS_40661953145378_0
timestamp 1698431365
transform 1 0 3798 0 1 55811
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_0
timestamp 1698431365
transform 1 0 6316 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_1
timestamp 1698431365
transform 1 0 6804 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_2
timestamp 1698431365
transform 1 0 7292 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_3
timestamp 1698431365
transform 1 0 4976 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_4
timestamp 1698431365
transform 1 0 5464 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_5
timestamp 1698431365
transform 1 0 5952 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_6
timestamp 1698431365
transform 1 0 7292 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_7
timestamp 1698431365
transform 1 0 6804 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_8
timestamp 1698431365
transform 1 0 6316 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_9
timestamp 1698431365
transform 1 0 5952 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_10
timestamp 1698431365
transform 1 0 5464 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_11
timestamp 1698431365
transform 1 0 4976 0 1 55368
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_12
timestamp 1698431365
transform 1 0 10708 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_13
timestamp 1698431365
transform 1 0 10220 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_14
timestamp 1698431365
transform 1 0 11196 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_15
timestamp 1698431365
transform 1 0 11196 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_16
timestamp 1698431365
transform 1 0 10220 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_17
timestamp 1698431365
transform 1 0 10708 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_18
timestamp 1698431365
transform 1 0 11560 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_19
timestamp 1698431365
transform 1 0 12048 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_20
timestamp 1698431365
transform 1 0 12536 0 1 53716
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_21
timestamp 1698431365
transform 1 0 12536 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_22
timestamp 1698431365
transform 1 0 12048 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145170  M3_M2_CDNS_40661953145170_23
timestamp 1698431365
transform 1 0 11560 0 1 55377
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_0
timestamp 1698431365
transform 1 0 4788 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_1
timestamp 1698431365
transform 1 0 7480 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_2
timestamp 1698431365
transform 1 0 7480 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_3
timestamp 1698431365
transform 1 0 6134 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_4
timestamp 1698431365
transform 1 0 6134 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_5
timestamp 1698431365
transform 1 0 4788 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_6
timestamp 1698431365
transform 1 0 10032 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_7
timestamp 1698431365
transform 1 0 10032 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_8
timestamp 1698431365
transform 1 0 12724 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_9
timestamp 1698431365
transform 1 0 12724 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_10
timestamp 1698431365
transform 1 0 11378 0 1 53706
box 0 0 1 1
use M3_M2_CDNS_40661953145172  M3_M2_CDNS_40661953145172_11
timestamp 1698431365
transform 1 0 11378 0 1 55287
box 0 0 1 1
use M3_M2_CDNS_40661953145174  M3_M2_CDNS_40661953145174_0
timestamp 1698431365
transform 1 0 11668 0 1 49762
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_0
timestamp 1698431365
transform 1 0 6087 0 1 37493
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_1
timestamp 1698431365
transform 1 0 84 0 1 37500
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_2
timestamp 1698431365
transform 1 0 3646 0 1 42293
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_3
timestamp 1698431365
transform 1 0 84 0 1 51900
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_4
timestamp 1698431365
transform 1 0 1924 0 1 53493
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_5
timestamp 1698431365
transform 1 0 3646 0 1 43893
box 0 0 1 1
use M3_M2_CDNS_40661953145179  M3_M2_CDNS_40661953145179_6
timestamp 1698431365
transform 1 0 14980 0 1 37493
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_0
timestamp 1698431365
transform 1 0 904 0 1 37493
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_1
timestamp 1698431365
transform 1 0 384 0 1 39093
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_2
timestamp 1698431365
transform 1 0 384 0 1 50293
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_3
timestamp 1698431365
transform 1 0 904 0 1 51893
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_4
timestamp 1698431365
transform 1 0 14580 0 1 29500
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_5
timestamp 1698431365
transform 1 0 14580 0 1 40693
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_6
timestamp 1698431365
transform 1 0 9349 0 1 53493
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_7
timestamp 1698431365
transform 1 0 14580 0 1 55100
box 0 0 1 1
use M3_M2_CDNS_40661953145180  M3_M2_CDNS_40661953145180_8
timestamp 1698431365
transform 1 0 14580 0 1 47093
box 0 0 1 1
use M3_M2_CDNS_40661953145186  M3_M2_CDNS_40661953145186_0
timestamp 1698431365
transform 1 0 6087 0 1 39229
box 0 0 1 1
use M3_M2_CDNS_40661953145186  M3_M2_CDNS_40661953145186_1
timestamp 1698431365
transform 1 0 3646 0 1 47235
box 0 0 1 1
use M3_M2_CDNS_40661953145186  M3_M2_CDNS_40661953145186_2
timestamp 1698431365
transform 1 0 10365 0 1 39235
box 0 0 1 1
use M3_M2_CDNS_40661953145186  M3_M2_CDNS_40661953145186_3
timestamp 1698431365
transform 1 0 10820 0 1 48835
box 0 0 1 1
use M3_M2_CDNS_40661953145186  M3_M2_CDNS_40661953145186_4
timestamp 1698431365
transform 1 0 11238 0 1 39235
box 0 0 1 1
use M3_M2_CDNS_40661953145188  M3_M2_CDNS_40661953145188_0
timestamp 1698431365
transform 1 0 2797 0 1 41044
box 0 0 1 1
use M3_M2_CDNS_40661953145190  M3_M2_CDNS_40661953145190_0
timestamp 1698431365
transform 1 0 7053 0 1 39448
box 0 0 1 1
use M3_M2_CDNS_40661953145190  M3_M2_CDNS_40661953145190_1
timestamp 1698431365
transform 1 0 5121 0 1 39448
box 0 0 1 1
use M3_M2_CDNS_40661953145190  M3_M2_CDNS_40661953145190_2
timestamp 1698431365
transform 1 0 1809 0 1 39448
box 0 0 1 1
use M3_M2_CDNS_40661953145190  M3_M2_CDNS_40661953145190_3
timestamp 1698431365
transform 1 0 11039 0 1 47432
box 0 0 1 1
use M3_M2_CDNS_40661953145193  M3_M2_CDNS_40661953145193_0
timestamp 1698431365
transform 1 0 8877 0 1 40288
box 0 0 1 1
use M3_M2_CDNS_40661953145194  M3_M2_CDNS_40661953145194_0
timestamp 1698431365
transform 1 0 13283 0 1 40288
box 0 0 1 1
use M3_M2_CDNS_40661953145194  M3_M2_CDNS_40661953145194_1
timestamp 1698431365
transform 1 0 10960 0 1 37542
box 0 0 1 1
use M3_M2_CDNS_40661953145196  M3_M2_CDNS_40661953145196_0
timestamp 1698431365
transform 1 0 4028 0 1 31954
box 0 0 1 1
use M3_M2_CDNS_40661953145196  M3_M2_CDNS_40661953145196_1
timestamp 1698431365
transform 1 0 524 0 1 35036
box 0 0 1 1
use M3_M2_CDNS_40661953145196  M3_M2_CDNS_40661953145196_2
timestamp 1698431365
transform 1 0 11036 0 1 31954
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_0
timestamp 1698431365
transform 1 0 4926 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_1
timestamp 1698431365
transform 1 0 762 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_2
timestamp 1698431365
transform 1 0 3130 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_3
timestamp 1698431365
transform 1 0 11934 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_4
timestamp 1698431365
transform 1 0 10138 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145197  M3_M2_CDNS_40661953145197_5
timestamp 1698431365
transform 1 0 8709 0 1 35244
box 0 0 1 1
use M3_M2_CDNS_40661953145199  M3_M2_CDNS_40661953145199_0
timestamp 1698431365
transform 1 0 4028 0 1 34851
box 0 0 1 1
use M3_M2_CDNS_40661953145199  M3_M2_CDNS_40661953145199_1
timestamp 1698431365
transform 1 0 11036 0 1 34851
box 0 0 1 1
use M3_M2_CDNS_40661953145200  M3_M2_CDNS_40661953145200_0
timestamp 1698431365
transform 1 0 524 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_0
timestamp 1698431365
transform 1 0 7050 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_1
timestamp 1698431365
transform 1 0 2814 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_2
timestamp 1698431365
transform 1 0 2398 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_3
timestamp 1698431365
transform 1 0 1006 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_4
timestamp 1698431365
transform 1 0 12666 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_5
timestamp 1698431365
transform 1 0 12250 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_6
timestamp 1698431365
transform 1 0 14058 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145202  M3_M2_CDNS_40661953145202_7
timestamp 1698431365
transform 1 0 8014 0 1 31599
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_0
timestamp 1698431365
transform 1 0 5658 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_1
timestamp 1698431365
transform 1 0 5242 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_2
timestamp 1698431365
transform 1 0 4754 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_3
timestamp 1698431365
transform 1 0 4266 0 1 31833
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_4
timestamp 1698431365
transform 1 0 3302 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_5
timestamp 1698431365
transform 1 0 3790 0 1 31833
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_6
timestamp 1698431365
transform 1 0 11762 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_7
timestamp 1698431365
transform 1 0 9406 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_8
timestamp 1698431365
transform 1 0 10798 0 1 31833
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_9
timestamp 1698431365
transform 1 0 10310 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_10
timestamp 1698431365
transform 1 0 9822 0 1 31884
box 0 0 1 1
use M3_M2_CDNS_40661953145204  M3_M2_CDNS_40661953145204_11
timestamp 1698431365
transform 1 0 11274 0 1 31833
box 0 0 1 1
use M3_M2_CDNS_40661953145206  M3_M2_CDNS_40661953145206_0
timestamp 1698431365
transform 1 0 2662 0 1 30081
box 0 0 1 1
use M3_M2_CDNS_40661953145206  M3_M2_CDNS_40661953145206_1
timestamp 1698431365
transform 1 0 12599 0 1 30081
box 0 0 1 1
use M3_M2_CDNS_40661953145207  M3_M2_CDNS_40661953145207_0
timestamp 1698431365
transform 1 0 14580 0 1 15900
box 0 0 1 1
use M3_M2_CDNS_40661953145207  M3_M2_CDNS_40661953145207_1
timestamp 1698431365
transform 1 0 14580 0 1 25500
box 0 0 1 1
use M3_M2_CDNS_40661953145207  M3_M2_CDNS_40661953145207_2
timestamp 1698431365
transform 1 0 14580 0 1 22300
box 0 0 1 1
use M3_M2_CDNS_40661953145207  M3_M2_CDNS_40661953145207_3
timestamp 1698431365
transform 1 0 14580 0 1 19100
box 0 0 1 1
use M3_M2_CDNS_40661953145207  M3_M2_CDNS_40661953145207_4
timestamp 1698431365
transform 1 0 14580 0 1 31900
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_0
timestamp 1698431365
transform 1 0 274 0 1 9500
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_1
timestamp 1698431365
transform 1 0 274 0 1 6300
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_2
timestamp 1698431365
transform 1 0 274 0 1 3100
box 0 0 1 1
use M3_M2_CDNS_40661953145208  M3_M2_CDNS_40661953145208_3
timestamp 1698431365
transform 1 0 274 0 1 35100
box 0 0 1 1
use M3_M2_CDNS_40661953145209  M3_M2_CDNS_40661953145209_0
timestamp 1698431365
transform 1 0 274 0 1 27900
box 0 0 1 1
use M3_M2_CDNS_40661953145209  M3_M2_CDNS_40661953145209_1
timestamp 1698431365
transform 1 0 12515 0 1 37493
box 0 0 1 1
use M3_M2_CDNS_40661953145210  M3_M2_CDNS_40661953145210_0
timestamp 1698431365
transform 1 0 1924 0 1 56639
box 0 0 1 1
use M3_M2_CDNS_40661953145210  M3_M2_CDNS_40661953145210_1
timestamp 1698431365
transform 1 0 14980 0 1 51893
box 0 0 1 1
use M3_M2_CDNS_40661953145212  M3_M2_CDNS_40661953145212_0
timestamp 1698431365
transform 1 0 8066 0 1 57010
box 0 0 1 1
use M3_M2_CDNS_40661953145212  M3_M2_CDNS_40661953145212_1
timestamp 1698431365
transform 1 0 8066 0 1 56268
box 0 0 1 1
use M3_M2_CDNS_40661953145213  M3_M2_CDNS_40661953145213_0
timestamp 1698431365
transform 1 0 13331 0 1 42380
box 0 0 1 1
use M3_M2_CDNS_40661953145314  M3_M2_CDNS_40661953145314_0
timestamp 1698431365
transform 1 0 10514 0 1 48008
box 0 0 1 1
use M3_M2_CDNS_40661953145330  M3_M2_CDNS_40661953145330_0
timestamp 1698431365
transform 1 0 10926 0 1 45474
box 0 0 1 1
use M3_M2_CDNS_40661953145330  M3_M2_CDNS_40661953145330_1
timestamp 1698431365
transform 1 0 11055 0 1 45474
box 0 0 1 1
use M3_M2_CDNS_40661953145332  M3_M2_CDNS_40661953145332_0
timestamp 1698431365
transform 1 0 3460 0 1 40288
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_0
timestamp 1698431365
transform 0 1 12482 1 0 41548
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_1
timestamp 1698431365
transform 0 1 13622 1 0 41548
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_2
timestamp 1698431365
transform 0 1 12482 1 0 42516
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314522  nmoscap_6p0_CDNS_4066195314522_3
timestamp 1698431365
transform 0 1 13622 1 0 42516
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_0
timestamp 1698431365
transform 0 1 4260 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_1
timestamp 1698431365
transform 0 1 5760 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_2
timestamp 1698431365
transform 0 1 2760 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_3
timestamp 1698431365
transform 0 1 8760 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_4
timestamp 1698431365
transform 0 1 13260 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_5
timestamp 1698431365
transform 0 1 11760 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_6
timestamp 1698431365
transform 0 1 10260 1 0 56489
box 0 0 1 1
use nmoscap_6p0_CDNS_4066195314523  nmoscap_6p0_CDNS_4066195314523_7
timestamp 1698431365
transform 0 1 7260 1 0 56489
box 0 0 1 1
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_0
timestamp 1698431365
transform 1 0 11458 0 1 41163
box 0 0 1 1
use pn_6p0_CDNS_4066195314528  pn_6p0_CDNS_4066195314528_1
timestamp 1698431365
transform 1 0 11458 0 1 41627
box 0 0 1 1
use ppolyf_u_CDNS_4066195314551  ppolyf_u_CDNS_4066195314551_0
timestamp 1698431365
transform 0 -1 939 1 0 55401
box 0 0 1 1
use ppolyf_u_CDNS_4066195314551  ppolyf_u_CDNS_4066195314551_1
timestamp 1698431365
transform 0 -1 1219 1 0 55401
box 0 0 1 1
<< labels >>
rlabel metal2 s 11512 29559 11512 29559 4 pdrive_x_<3>
port 1 nsew
rlabel metal2 s 10870 29559 10870 29559 4 pdrive_y_<3>
port 2 nsew
rlabel metal2 s 10062 29559 10062 29559 4 pdrive_y_<2>
port 3 nsew
rlabel metal2 s 9110 29559 9110 29559 4 pdrive_x_<2>
port 4 nsew
rlabel metal2 s 5954 29559 5954 29559 4 pdrive_x_<1>
port 5 nsew
rlabel metal2 s 4995 29559 4995 29559 4 pdrive_y_<1>
port 6 nsew
rlabel metal2 s 4188 29559 4188 29559 4 pdrive_y_<0>
port 7 nsew
rlabel metal2 s 3547 29559 3547 29559 4 pdrive_x_<0>
port 8 nsew
rlabel metal2 s 14010 29559 14010 29559 4 ndrive_Y_<3>
port 9 nsew
rlabel metal2 s 13824 29559 13824 29559 4 ndrive_x_<3>
port 10 nsew
rlabel metal2 s 13647 29559 13647 29559 4 ndrive_y_<2>
port 11 nsew
rlabel metal2 s 13463 29559 13463 29559 4 ndrive_x_<2>
port 12 nsew
rlabel metal2 s 1594 29559 1594 29559 4 ndrive_Y_<1>
port 13 nsew
rlabel metal2 s 1408 29559 1408 29559 4 ndrive_x_<1>
port 14 nsew
rlabel metal2 s 1231 29559 1231 29559 4 ndrive_y_<0>
port 15 nsew
rlabel metal2 s 1047 29559 1047 29559 4 ndrive_x_<0>
port 16 nsew
rlabel metal2 s 14242 57528 14242 57528 4 Y
port 17 nsew
rlabel metal2 s 1263 57483 1263 57483 4 PU
port 18 nsew
rlabel metal2 s 7532 28487 7532 28487 4 PAD
port 19 nsew
rlabel metal2 s 2136 57487 2136 57487 4 PD
port 20 nsew
<< properties >>
string GDS_END 17675458
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 17636180
string path 17.600 1432.525 353.350 1432.525 
<< end >>
