magic
tech gf180mcuD
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 453 2774 1094
<< pwell >>
rect -86 -86 2774 453
<< mvnmos >>
rect 124 138 244 296
rect 392 156 512 296
rect 560 156 680 296
rect 728 156 848 296
rect 952 156 1072 296
rect 1120 156 1240 296
rect 1288 156 1408 296
rect 1548 156 1668 314
rect 1716 156 1836 314
rect 2084 175 2204 333
rect 2352 69 2472 333
<< mvpmos >>
rect 124 573 224 849
rect 484 648 584 848
rect 688 648 788 848
rect 836 648 936 848
rect 1040 648 1140 848
rect 1200 648 1300 848
rect 1404 648 1504 848
rect 1656 574 1756 850
rect 2116 574 2216 850
rect 2356 574 2456 940
<< mvndiff >>
rect 1996 320 2084 333
rect 1468 296 1548 314
rect 36 215 124 296
rect 36 169 49 215
rect 95 169 124 215
rect 36 138 124 169
rect 244 205 392 296
rect 244 159 273 205
rect 319 159 392 205
rect 244 156 392 159
rect 512 156 560 296
rect 680 156 728 296
rect 848 215 952 296
rect 848 169 877 215
rect 923 169 952 215
rect 848 156 952 169
rect 1072 156 1120 296
rect 1240 156 1288 296
rect 1408 215 1548 296
rect 1408 169 1437 215
rect 1483 169 1548 215
rect 1408 156 1548 169
rect 1668 156 1716 314
rect 1836 215 1924 314
rect 1836 169 1865 215
rect 1911 169 1924 215
rect 1996 274 2009 320
rect 2055 274 2084 320
rect 1996 175 2084 274
rect 2204 222 2352 333
rect 2204 175 2277 222
rect 1836 156 1924 169
rect 244 138 332 156
rect 2264 82 2277 175
rect 2323 82 2352 222
rect 2264 69 2352 82
rect 2472 320 2560 333
rect 2472 180 2501 320
rect 2547 180 2560 320
rect 2472 69 2560 180
<< mvpdiff >>
rect 36 831 124 849
rect 36 691 49 831
rect 95 691 124 831
rect 36 573 124 691
rect 224 831 312 849
rect 2276 850 2356 940
rect 1576 848 1656 850
rect 224 691 253 831
rect 299 691 312 831
rect 224 573 312 691
rect 396 831 484 848
rect 396 691 409 831
rect 455 691 484 831
rect 396 648 484 691
rect 584 835 688 848
rect 584 789 613 835
rect 659 789 688 835
rect 584 648 688 789
rect 788 648 836 848
rect 936 831 1040 848
rect 936 691 965 831
rect 1011 691 1040 831
rect 936 648 1040 691
rect 1140 648 1200 848
rect 1300 835 1404 848
rect 1300 789 1329 835
rect 1375 789 1404 835
rect 1300 648 1404 789
rect 1504 831 1656 848
rect 1504 691 1581 831
rect 1627 691 1656 831
rect 1504 648 1656 691
rect 1576 574 1656 648
rect 1756 831 1844 850
rect 1756 691 1785 831
rect 1831 691 1844 831
rect 1756 574 1844 691
rect 2028 831 2116 850
rect 2028 691 2041 831
rect 2087 691 2116 831
rect 2028 574 2116 691
rect 2216 837 2356 850
rect 2216 697 2245 837
rect 2291 697 2356 837
rect 2216 574 2356 697
rect 2456 831 2544 940
rect 2456 691 2485 831
rect 2531 691 2544 831
rect 2456 574 2544 691
<< mvndiffc >>
rect 49 169 95 215
rect 273 159 319 205
rect 877 169 923 215
rect 1437 169 1483 215
rect 1865 169 1911 215
rect 2009 274 2055 320
rect 2277 82 2323 222
rect 2501 180 2547 320
<< mvpdiffc >>
rect 49 691 95 831
rect 253 691 299 831
rect 409 691 455 831
rect 613 789 659 835
rect 965 691 1011 831
rect 1329 789 1375 835
rect 1581 691 1627 831
rect 1785 691 1831 831
rect 2041 691 2087 831
rect 2245 697 2291 837
rect 2485 691 2531 831
<< polysilicon >>
rect 2356 940 2456 984
rect 124 849 224 893
rect 484 848 584 892
rect 688 848 788 892
rect 836 848 936 892
rect 1040 848 1140 892
rect 1200 848 1300 892
rect 1404 848 1504 892
rect 1656 850 1756 894
rect 2116 850 2216 894
rect 484 604 584 648
rect 688 604 788 648
rect 836 604 936 648
rect 124 501 224 573
rect 484 514 524 604
rect 688 514 728 604
rect 896 546 936 604
rect 896 533 992 546
rect 124 455 152 501
rect 198 455 224 501
rect 124 340 224 455
rect 392 501 524 514
rect 392 455 453 501
rect 499 485 524 501
rect 608 501 728 514
rect 499 455 512 485
rect 124 296 244 340
rect 392 296 512 455
rect 608 455 621 501
rect 667 474 728 501
rect 776 501 848 514
rect 667 455 680 474
rect 608 340 680 455
rect 776 455 789 501
rect 835 455 848 501
rect 896 487 909 533
rect 955 487 992 533
rect 896 474 992 487
rect 776 340 848 455
rect 560 296 680 340
rect 728 296 848 340
rect 952 340 992 474
rect 1040 501 1140 648
rect 1040 455 1053 501
rect 1099 455 1140 501
rect 1040 442 1140 455
rect 1200 604 1300 648
rect 1404 615 1504 648
rect 1200 514 1240 604
rect 1404 569 1417 615
rect 1463 569 1504 615
rect 1404 514 1504 569
rect 1656 530 1756 574
rect 1716 514 1756 530
rect 2116 530 2216 574
rect 2116 514 2204 530
rect 2356 514 2456 574
rect 1200 501 1296 514
rect 1200 455 1237 501
rect 1283 455 1296 501
rect 1404 474 1588 514
rect 1200 442 1296 455
rect 1200 340 1240 442
rect 1548 358 1588 474
rect 1716 501 1788 514
rect 1716 455 1729 501
rect 1775 455 1788 501
rect 1716 358 1788 455
rect 2084 501 2204 514
rect 2084 455 2097 501
rect 2143 455 2204 501
rect 952 296 1072 340
rect 1120 296 1240 340
rect 1288 296 1408 340
rect 1548 314 1668 358
rect 1716 314 1836 358
rect 2084 333 2204 455
rect 2324 501 2456 514
rect 2324 455 2337 501
rect 2383 455 2456 501
rect 2324 442 2456 455
rect 2352 377 2456 442
rect 2352 333 2472 377
rect 124 94 244 138
rect 392 64 512 156
rect 560 112 680 156
rect 728 112 848 156
rect 952 112 1072 156
rect 1120 112 1240 156
rect 1288 64 1408 156
rect 1548 112 1668 156
rect 1716 112 1836 156
rect 2084 131 2204 175
rect 392 24 1408 64
rect 2352 25 2472 69
<< polycontact >>
rect 152 455 198 501
rect 453 455 499 501
rect 621 455 667 501
rect 789 455 835 501
rect 909 487 955 533
rect 1053 455 1099 501
rect 1417 569 1463 615
rect 1237 455 1283 501
rect 1729 455 1775 501
rect 2097 455 2143 501
rect 2337 455 2383 501
<< metal1 >>
rect 0 918 2688 1098
rect 49 831 95 842
rect 49 634 95 691
rect 253 831 299 918
rect 253 680 299 691
rect 409 831 455 842
rect 613 835 659 918
rect 613 778 659 789
rect 965 831 1011 842
rect 455 691 965 726
rect 1329 835 1375 918
rect 1329 778 1375 789
rect 1581 831 1627 842
rect 1011 691 1463 726
rect 409 680 1463 691
rect 49 588 955 634
rect 1417 615 1463 680
rect 49 215 95 588
rect 366 501 499 542
rect 141 455 152 501
rect 198 455 320 501
rect 274 308 320 455
rect 366 455 453 501
rect 366 354 499 455
rect 590 501 667 542
rect 909 533 955 588
rect 590 455 621 501
rect 590 354 667 455
rect 789 501 835 512
rect 1145 569 1417 604
rect 1581 634 1627 691
rect 1785 831 1831 918
rect 1785 680 1831 691
rect 2041 831 2087 842
rect 2041 640 2087 691
rect 2245 837 2291 918
rect 2245 686 2291 697
rect 2485 831 2547 842
rect 2531 691 2547 831
rect 1581 588 1911 634
rect 2041 594 2383 640
rect 1145 558 1463 569
rect 909 476 955 487
rect 1053 501 1099 512
rect 789 430 835 455
rect 1053 430 1099 455
rect 789 354 1099 430
rect 789 308 835 354
rect 274 262 835 308
rect 1145 226 1191 558
rect 1237 501 1283 512
rect 1237 308 1283 455
rect 1710 501 1775 542
rect 1710 455 1729 501
rect 1710 354 1775 455
rect 1865 512 1911 588
rect 1865 501 2143 512
rect 1865 455 2097 501
rect 1865 444 2143 455
rect 2337 501 2383 594
rect 1865 308 1911 444
rect 2337 331 2383 455
rect 1237 262 1911 308
rect 2009 320 2383 331
rect 2055 285 2383 320
rect 2485 320 2547 691
rect 2009 263 2055 274
rect 49 158 95 169
rect 273 205 319 216
rect 273 90 319 159
rect 877 215 1191 226
rect 1865 215 1911 262
rect 923 169 1191 215
rect 877 158 1191 169
rect 1426 169 1437 215
rect 1483 169 1494 215
rect 1426 90 1494 169
rect 1865 158 1911 169
rect 2277 222 2323 233
rect 0 82 2277 90
rect 2485 180 2501 320
rect 2485 169 2547 180
rect 2323 82 2688 90
rect 0 -90 2688 82
<< labels >>
flabel metal1 s 590 354 667 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 1053 501 1099 512 0 FreeSans 200 0 0 0 E
port 2 nsew clock input
flabel metal1 s 2485 169 2547 842 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 366 354 499 542 0 FreeSans 200 0 0 0 RN
port 3 nsew default input
flabel metal1 s 1710 354 1775 542 0 FreeSans 200 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 0 918 2688 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2277 216 2323 233 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 7 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 8 nsew ground bidirectional
rlabel metal1 s 789 501 835 512 1 E
port 2 nsew clock input
rlabel metal1 s 1053 455 1099 501 1 E
port 2 nsew clock input
rlabel metal1 s 789 455 835 501 1 E
port 2 nsew clock input
rlabel metal1 s 141 455 320 501 1 E
port 2 nsew clock input
rlabel metal1 s 1053 430 1099 455 1 E
port 2 nsew clock input
rlabel metal1 s 789 430 835 455 1 E
port 2 nsew clock input
rlabel metal1 s 274 430 320 455 1 E
port 2 nsew clock input
rlabel metal1 s 789 354 1099 430 1 E
port 2 nsew clock input
rlabel metal1 s 274 354 320 430 1 E
port 2 nsew clock input
rlabel metal1 s 789 308 835 354 1 E
port 2 nsew clock input
rlabel metal1 s 274 308 320 354 1 E
port 2 nsew clock input
rlabel metal1 s 274 262 835 308 1 E
port 2 nsew clock input
rlabel metal1 s 2245 778 2291 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1785 778 1831 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1329 778 1375 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 613 778 659 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 778 299 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2245 686 2291 778 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1785 686 1831 778 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 686 299 778 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1785 680 1831 686 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 680 299 686 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2277 215 2323 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 215 319 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2277 90 2323 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1426 90 1494 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2688 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2688 1008
string GDS_END 1031682
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1024720
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
