magic
tech gf180mcuC
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 407 3894 870
rect -86 352 575 407
rect 943 352 3894 407
<< pwell >>
rect 575 352 943 407
rect -86 -86 3894 352
<< metal1 >>
rect 0 724 3808 844
rect 290 652 358 724
rect 1058 657 1126 724
rect 109 355 335 437
rect 1466 657 1534 724
rect 1874 657 1942 724
rect 2078 553 2146 676
rect 2282 657 2350 724
rect 2486 553 2554 676
rect 2690 657 2758 724
rect 2894 553 2962 676
rect 3098 657 3166 724
rect 3302 553 3370 676
rect 3506 657 3574 724
rect 2078 485 3370 553
rect 1015 360 1886 424
rect 2684 227 2814 485
rect 2080 173 3510 227
rect 262 60 330 131
rect 934 60 1002 95
rect 1426 60 1494 127
rect 1874 60 1942 127
rect 2322 60 2390 127
rect 2770 60 2838 127
rect 3218 60 3286 127
rect 3666 60 3734 127
rect 0 -60 3808 60
<< obsm1 >>
rect 536 632 965 678
rect 84 556 431 602
rect 385 504 431 556
rect 385 447 730 504
rect 385 265 431 447
rect 778 401 846 586
rect 38 219 431 265
rect 641 355 846 401
rect 919 552 965 632
rect 1273 552 1319 676
rect 1681 552 1727 676
rect 919 506 1997 552
rect 38 170 106 219
rect 641 152 687 355
rect 919 309 965 506
rect 1951 439 1997 506
rect 1951 393 2452 439
rect 754 263 965 309
rect 1951 273 2504 319
rect 754 228 822 263
rect 1951 219 1997 273
rect 3010 393 3486 439
rect 3083 273 3598 319
rect 1139 187 1997 219
rect 843 173 1997 187
rect 843 152 1189 173
rect 478 141 1189 152
rect 478 106 888 141
<< labels >>
rlabel metal1 s 109 355 335 437 6 EN
port 1 nsew default input
rlabel metal1 s 1015 360 1886 424 6 I
port 2 nsew default input
rlabel metal1 s 2080 173 3510 227 6 Z
port 3 nsew default output
rlabel metal1 s 2684 227 2814 485 6 Z
port 3 nsew default output
rlabel metal1 s 2078 485 3370 553 6 Z
port 3 nsew default output
rlabel metal1 s 3302 553 3370 676 6 Z
port 3 nsew default output
rlabel metal1 s 2894 553 2962 676 6 Z
port 3 nsew default output
rlabel metal1 s 2486 553 2554 676 6 Z
port 3 nsew default output
rlabel metal1 s 2078 553 2146 676 6 Z
port 3 nsew default output
rlabel metal1 s 3506 657 3574 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3098 657 3166 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2690 657 2758 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2282 657 2350 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1874 657 1942 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1466 657 1534 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1058 657 1126 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 290 652 358 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 724 3808 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel nwell s 943 352 3894 407 6 VNW
port 5 nsew power bidirectional
rlabel nwell s -86 352 575 407 6 VNW
port 5 nsew power bidirectional
rlabel nwell s -86 407 3894 870 6 VNW
port 5 nsew power bidirectional
rlabel pwell s -86 -86 3894 352 6 VPW
port 6 nsew ground bidirectional
rlabel pwell s 575 352 943 407 6 VPW
port 6 nsew ground bidirectional
rlabel metal1 s 0 -60 3808 60 8 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3666 60 3734 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3218 60 3286 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2770 60 2838 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2322 60 2390 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1874 60 1942 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1426 60 1494 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 95 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 131 6 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1417210
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1408920
<< end >>
