magic
tech gf180mcuC
magscale 1 5
timestamp 1698431365
<< nwell >>
rect -43 176 3627 435
<< pwell >>
rect -43 -43 3627 176
<< metal1 >>
rect 0 362 3584 422
rect 0 -30 3584 30
<< labels >>
flabel metal1 s 0 362 3584 422 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 0 -30 3584 30 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell s 5 367 55 417 0 FreeSans 200 0 0 0 VNW
port 2 nsew power bidirectional
flabel pwell s 5 -25 55 25 0 FreeSans 200 0 0 0 VPW
port 3 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 3584 392
string GDS_END 1154596
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1153436
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
