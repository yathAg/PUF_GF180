magic
tech gf180mcuA
magscale 1 10
timestamp 1698431365
<< nwell >>
rect -86 377 3110 870
rect -86 352 988 377
rect 2799 352 3110 377
<< pwell >>
rect -86 -86 3110 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1164 93 1284 257
rect 1388 93 1508 257
rect 1612 93 1732 257
rect 1836 93 1956 257
rect 2060 93 2180 257
rect 2284 93 2404 257
rect 2508 93 2628 257
rect 2776 68 2896 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 572 497 672 716
rect 816 497 916 716
rect 1184 497 1284 716
rect 1408 497 1508 716
rect 1612 497 1712 716
rect 1836 497 1936 716
rect 2080 497 2180 716
rect 2304 497 2404 716
rect 2508 497 2608 716
rect 2776 497 2876 716
<< mvndiff >>
rect 36 158 124 232
rect 36 112 49 158
rect 95 112 124 158
rect 36 68 124 112
rect 244 219 348 232
rect 244 173 273 219
rect 319 173 348 219
rect 244 68 348 173
rect 468 127 572 232
rect 468 81 497 127
rect 543 81 572 127
rect 468 68 572 81
rect 692 219 796 232
rect 692 173 721 219
rect 767 173 796 219
rect 692 68 796 173
rect 916 127 1004 232
rect 916 81 945 127
rect 991 81 1004 127
rect 1076 152 1164 257
rect 1076 106 1089 152
rect 1135 106 1164 152
rect 1076 93 1164 106
rect 1284 244 1388 257
rect 1284 198 1313 244
rect 1359 198 1388 244
rect 1284 93 1388 198
rect 1508 152 1612 257
rect 1508 106 1537 152
rect 1583 106 1612 152
rect 1508 93 1612 106
rect 1732 244 1836 257
rect 1732 198 1761 244
rect 1807 198 1836 244
rect 1732 93 1836 198
rect 1956 152 2060 257
rect 1956 106 1985 152
rect 2031 106 2060 152
rect 1956 93 2060 106
rect 2180 244 2284 257
rect 2180 198 2209 244
rect 2255 198 2284 244
rect 2180 93 2284 198
rect 2404 152 2508 257
rect 2404 106 2433 152
rect 2479 106 2508 152
rect 2404 93 2508 106
rect 2628 244 2716 257
rect 2628 198 2657 244
rect 2703 232 2716 244
rect 2703 198 2776 232
rect 2628 93 2776 198
rect 916 68 1004 81
rect 2696 68 2776 93
rect 2896 152 2984 232
rect 2896 106 2925 152
rect 2971 106 2984 152
rect 2896 68 2984 106
<< mvpdiff >>
rect 56 611 144 716
rect 56 565 69 611
rect 115 565 144 611
rect 56 497 144 565
rect 244 497 368 716
rect 468 703 572 716
rect 468 657 497 703
rect 543 657 572 703
rect 468 497 572 657
rect 672 497 816 716
rect 916 639 1184 716
rect 916 593 945 639
rect 991 593 1109 639
rect 1155 593 1184 639
rect 916 497 1184 593
rect 1284 497 1408 716
rect 1508 703 1612 716
rect 1508 657 1537 703
rect 1583 657 1612 703
rect 1508 497 1612 657
rect 1712 497 1836 716
rect 1936 639 2080 716
rect 1936 593 1985 639
rect 2031 593 2080 639
rect 1936 497 2080 593
rect 2180 497 2304 716
rect 2404 703 2508 716
rect 2404 657 2433 703
rect 2479 657 2508 703
rect 2404 497 2508 657
rect 2608 497 2776 716
rect 2876 639 2964 716
rect 2876 593 2905 639
rect 2951 593 2964 639
rect 2876 497 2964 593
<< mvndiffc >>
rect 49 112 95 158
rect 273 173 319 219
rect 497 81 543 127
rect 721 173 767 219
rect 945 81 991 127
rect 1089 106 1135 152
rect 1313 198 1359 244
rect 1537 106 1583 152
rect 1761 198 1807 244
rect 1985 106 2031 152
rect 2209 198 2255 244
rect 2433 106 2479 152
rect 2657 198 2703 244
rect 2925 106 2971 152
<< mvpdiffc >>
rect 69 565 115 611
rect 497 657 543 703
rect 945 593 991 639
rect 1109 593 1155 639
rect 1537 657 1583 703
rect 1985 593 2031 639
rect 2433 657 2479 703
rect 2905 593 2951 639
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 1184 716 1284 760
rect 1408 716 1508 760
rect 1612 716 1712 760
rect 1836 716 1936 760
rect 2080 716 2180 760
rect 2304 716 2404 760
rect 2508 716 2608 760
rect 2776 716 2876 760
rect 144 402 244 497
rect 368 415 468 497
rect 368 402 395 415
rect 124 365 244 402
rect 124 319 144 365
rect 190 319 244 365
rect 124 232 244 319
rect 348 369 395 402
rect 441 394 468 415
rect 572 415 672 497
rect 572 394 599 415
rect 441 369 599 394
rect 645 402 672 415
rect 816 402 916 497
rect 1184 415 1284 497
rect 1184 402 1211 415
rect 645 369 692 402
rect 348 348 692 369
rect 348 232 468 348
rect 572 232 692 348
rect 796 365 916 402
rect 796 319 819 365
rect 865 319 916 365
rect 796 232 916 319
rect 1164 369 1211 402
rect 1257 369 1284 415
rect 1408 415 1508 497
rect 1408 402 1435 415
rect 1164 257 1284 369
rect 1388 369 1435 402
rect 1481 394 1508 415
rect 1612 415 1712 497
rect 1612 394 1639 415
rect 1481 369 1639 394
rect 1685 402 1712 415
rect 1836 415 1936 497
rect 1685 369 1732 402
rect 1388 348 1732 369
rect 1388 257 1508 348
rect 1612 257 1732 348
rect 1836 369 1865 415
rect 1911 402 1936 415
rect 2080 402 2180 497
rect 2304 415 2404 497
rect 2304 402 2331 415
rect 1911 369 1956 402
rect 1836 257 1956 369
rect 2060 394 2180 402
rect 2060 348 2115 394
rect 2161 348 2180 394
rect 2060 257 2180 348
rect 2284 369 2331 402
rect 2377 394 2404 415
rect 2508 415 2608 497
rect 2508 394 2535 415
rect 2377 369 2535 394
rect 2581 402 2608 415
rect 2776 415 2876 497
rect 2581 369 2628 402
rect 2284 348 2628 369
rect 2284 257 2404 348
rect 2508 257 2628 348
rect 2776 369 2806 415
rect 2852 402 2876 415
rect 2852 369 2896 402
rect 2776 232 2896 369
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1164 24 1284 93
rect 1388 24 1508 93
rect 1612 24 1732 93
rect 1836 24 1956 93
rect 2060 24 2180 93
rect 2284 24 2404 93
rect 2508 24 2628 93
rect 2776 24 2896 68
<< polycontact >>
rect 144 319 190 365
rect 395 369 441 415
rect 599 369 645 415
rect 819 319 865 365
rect 1211 369 1257 415
rect 1435 369 1481 415
rect 1639 369 1685 415
rect 1865 369 1911 415
rect 2115 348 2161 394
rect 2331 369 2377 415
rect 2535 369 2581 415
rect 2806 369 2852 415
<< metal1 >>
rect 0 724 3024 844
rect 486 703 554 724
rect 486 657 497 703
rect 543 657 554 703
rect 1526 703 1594 724
rect 1526 657 1537 703
rect 1583 657 1594 703
rect 2422 703 2490 724
rect 2422 657 2433 703
rect 2479 657 2490 703
rect 625 639 1468 648
rect 625 611 945 639
rect 56 565 69 611
rect 115 593 945 611
rect 991 593 1109 639
rect 1155 611 1468 639
rect 1689 639 2355 648
rect 1689 611 1985 639
rect 1155 593 1985 611
rect 2031 611 2355 639
rect 2544 639 2964 648
rect 2544 611 2905 639
rect 2031 593 2905 611
rect 2951 593 2964 639
rect 115 584 2964 593
rect 115 565 684 584
rect 1418 565 2590 584
rect 1014 519 1348 538
rect 1014 473 1876 519
rect 132 365 204 438
rect 132 319 144 365
rect 190 319 204 365
rect 306 415 692 424
rect 306 369 395 415
rect 441 369 599 415
rect 645 369 692 415
rect 306 360 692 369
rect 802 365 1003 424
rect 132 314 204 319
rect 802 319 819 365
rect 865 360 1003 365
rect 1208 415 1260 473
rect 1820 430 1876 473
rect 1208 369 1211 415
rect 1257 369 1260 415
rect 865 319 876 360
rect 1208 358 1260 369
rect 1354 415 1774 424
rect 1354 369 1435 415
rect 1481 369 1639 415
rect 1685 369 1774 415
rect 1354 360 1774 369
rect 1820 415 1936 430
rect 1820 369 1865 415
rect 1911 369 1936 415
rect 1820 354 1936 369
rect 802 314 876 319
rect 132 267 876 314
rect 1986 244 2032 565
rect 2657 519 2892 538
rect 2105 473 2892 519
rect 2105 394 2212 473
rect 2105 348 2115 394
rect 2161 348 2212 394
rect 2258 415 2678 424
rect 2258 369 2331 415
rect 2377 369 2535 415
rect 2581 369 2678 415
rect 2258 360 2678 369
rect 2801 415 2892 473
rect 2801 369 2806 415
rect 2852 369 2892 415
rect 2105 329 2212 348
rect 976 219 1313 244
rect 262 173 273 219
rect 319 173 721 219
rect 767 198 1313 219
rect 1359 198 1761 244
rect 1807 198 1818 244
rect 1986 198 2209 244
rect 2255 198 2657 244
rect 2703 198 2714 244
rect 2801 232 2892 369
rect 767 173 1026 198
rect 49 158 95 169
rect 49 60 95 112
rect 486 81 497 127
rect 543 81 554 127
rect 486 60 554 81
rect 934 81 945 127
rect 991 81 1002 127
rect 1078 106 1089 152
rect 1135 106 1537 152
rect 1583 106 1985 152
rect 2031 106 2433 152
rect 2479 106 2925 152
rect 2971 106 2984 152
rect 934 60 1002 81
rect 0 -60 3024 60
<< labels >>
flabel metal1 s 1014 519 1348 538 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 1354 360 1774 424 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel metal1 s 132 424 204 438 0 FreeSans 400 0 0 0 C1
port 5 nsew default input
flabel metal1 s 306 360 692 424 0 FreeSans 400 0 0 0 C2
port 6 nsew default input
flabel metal1 s 0 724 3024 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 49 127 95 169 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 2544 611 2964 648 0 FreeSans 400 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 2657 519 2892 538 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 2258 360 2678 424 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell s 10 734 110 834 0 FreeSans 400 0 0 0 VNW
port 9 nsew power bidirectional
flabel pwell s 10 -50 110 50 0 FreeSans 400 0 0 0 VPW
port 10 nsew ground bidirectional
rlabel metal1 s 2105 473 2892 519 1 A1
port 1 nsew default input
rlabel metal1 s 2801 329 2892 473 1 A1
port 1 nsew default input
rlabel metal1 s 2105 329 2212 473 1 A1
port 1 nsew default input
rlabel metal1 s 2801 232 2892 329 1 A1
port 1 nsew default input
rlabel metal1 s 1014 473 1876 519 1 B1
port 3 nsew default input
rlabel metal1 s 1820 430 1876 473 1 B1
port 3 nsew default input
rlabel metal1 s 1208 430 1260 473 1 B1
port 3 nsew default input
rlabel metal1 s 1820 358 1936 430 1 B1
port 3 nsew default input
rlabel metal1 s 1208 358 1260 430 1 B1
port 3 nsew default input
rlabel metal1 s 1820 354 1936 358 1 B1
port 3 nsew default input
rlabel metal1 s 802 360 1003 424 1 C1
port 5 nsew default input
rlabel metal1 s 132 360 204 424 1 C1
port 5 nsew default input
rlabel metal1 s 802 314 876 360 1 C1
port 5 nsew default input
rlabel metal1 s 132 314 204 360 1 C1
port 5 nsew default input
rlabel metal1 s 132 267 876 314 1 C1
port 5 nsew default input
rlabel metal1 s 1689 611 2355 648 1 ZN
port 7 nsew default output
rlabel metal1 s 625 611 1468 648 1 ZN
port 7 nsew default output
rlabel metal1 s 56 584 2964 611 1 ZN
port 7 nsew default output
rlabel metal1 s 1418 565 2590 584 1 ZN
port 7 nsew default output
rlabel metal1 s 56 565 684 584 1 ZN
port 7 nsew default output
rlabel metal1 s 1986 244 2032 565 1 ZN
port 7 nsew default output
rlabel metal1 s 1986 198 2714 244 1 ZN
port 7 nsew default output
rlabel metal1 s 2422 657 2490 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1526 657 1594 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 486 657 554 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 934 60 1002 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 1 VSS
port 11 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3024 60 1 VSS
port 11 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3024 784
string GDS_END 133736
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 127598
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
